magic
tech scmos
timestamp 1607319584
<< metal1 >>
rect 1048 4903 1050 4907
rect 1054 4903 1057 4907
rect 1061 4903 1064 4907
rect 2072 4903 2074 4907
rect 2078 4903 2081 4907
rect 2085 4903 2088 4907
rect 3096 4903 3098 4907
rect 3102 4903 3105 4907
rect 3109 4903 3112 4907
rect 4112 4903 4114 4907
rect 4118 4903 4121 4907
rect 4125 4903 4128 4907
rect 726 4878 738 4881
rect 834 4878 841 4881
rect 734 4877 738 4878
rect 70 4868 78 4871
rect 250 4858 257 4861
rect 310 4858 318 4861
rect 686 4862 689 4871
rect 1262 4871 1265 4881
rect 3398 4878 3417 4881
rect 3422 4878 3434 4881
rect 3838 4878 3857 4881
rect 1830 4876 1834 4878
rect 3430 4877 3434 4878
rect 1262 4868 1281 4871
rect 1562 4868 1570 4871
rect 642 4858 649 4861
rect 702 4858 710 4861
rect 878 4858 881 4868
rect 1174 4858 1190 4861
rect 1378 4858 1385 4861
rect 1534 4858 1542 4861
rect 1790 4862 1793 4871
rect 1890 4868 1897 4871
rect 2566 4868 2598 4871
rect 2898 4868 2905 4871
rect 3518 4868 3530 4871
rect 4230 4871 4233 4881
rect 4214 4868 4233 4871
rect 4494 4868 4502 4871
rect 4574 4868 4585 4871
rect 1806 4858 1814 4861
rect 2102 4858 2121 4861
rect 2286 4858 2294 4861
rect 2426 4858 2433 4861
rect 2438 4858 2446 4861
rect 2686 4858 2694 4861
rect 2706 4858 2713 4861
rect 2718 4858 2726 4861
rect 3074 4858 3081 4861
rect 3086 4858 3094 4861
rect 3358 4858 3366 4861
rect 3398 4858 3401 4868
rect 3786 4858 3793 4861
rect 4574 4862 4577 4868
rect 570 4848 574 4852
rect 2102 4848 2105 4858
rect 2682 4848 2686 4852
rect 955 4838 958 4842
rect 1211 4838 1214 4842
rect 1714 4838 1717 4842
rect 2230 4838 2242 4841
rect 2253 4838 2254 4842
rect 3043 4838 3046 4842
rect 3187 4838 3190 4842
rect 3226 4838 3227 4842
rect 3315 4838 3318 4842
rect 4086 4818 4094 4821
rect 5021 4818 5022 4822
rect 536 4803 538 4807
rect 542 4803 545 4807
rect 549 4803 552 4807
rect 1560 4803 1562 4807
rect 1566 4803 1569 4807
rect 1573 4803 1576 4807
rect 2584 4803 2586 4807
rect 2590 4803 2593 4807
rect 2597 4803 2600 4807
rect 3608 4803 3610 4807
rect 3614 4803 3617 4807
rect 3621 4803 3624 4807
rect 4632 4803 4634 4807
rect 4638 4803 4641 4807
rect 4645 4803 4648 4807
rect 194 4788 195 4792
rect 322 4788 323 4792
rect 482 4788 483 4792
rect 562 4788 563 4792
rect 1685 4788 1686 4792
rect 1738 4788 1739 4792
rect 2506 4788 2507 4792
rect 3397 4788 3398 4792
rect 3461 4788 3462 4792
rect 4677 4788 4678 4792
rect 4101 4778 4102 4782
rect 730 4768 738 4771
rect 2147 4768 2150 4772
rect 3429 4768 3430 4772
rect 3914 4768 3917 4772
rect 4619 4768 4622 4772
rect 3806 4766 3810 4768
rect 4694 4766 4698 4768
rect 126 4751 129 4761
rect 126 4748 145 4751
rect 334 4751 337 4761
rect 334 4748 353 4751
rect 426 4748 433 4751
rect 494 4751 497 4761
rect 690 4758 694 4762
rect 810 4758 814 4762
rect 1618 4758 1622 4762
rect 2186 4758 2190 4762
rect 2218 4758 2222 4762
rect 494 4748 513 4751
rect 518 4748 558 4751
rect 726 4751 729 4758
rect 726 4748 745 4751
rect 782 4748 790 4751
rect 882 4748 889 4751
rect 958 4748 966 4751
rect 1570 4748 1585 4751
rect 1642 4748 1649 4751
rect 1654 4748 1670 4751
rect 1686 4748 1702 4751
rect 1810 4748 1817 4751
rect 1962 4748 1969 4751
rect 2270 4748 2278 4751
rect 2366 4751 2369 4761
rect 2350 4748 2369 4751
rect 2574 4748 2582 4751
rect 2726 4751 2729 4761
rect 2738 4758 2742 4762
rect 3586 4758 3590 4762
rect 2710 4748 2729 4751
rect 3254 4742 3257 4751
rect 3598 4751 3601 4761
rect 3598 4748 3633 4751
rect 3862 4751 3865 4761
rect 3846 4748 3865 4751
rect 4042 4748 4049 4751
rect 4166 4751 4169 4761
rect 4150 4748 4169 4751
rect 4250 4748 4257 4751
rect 4454 4748 4470 4751
rect 4770 4748 4777 4751
rect 4982 4748 4990 4751
rect 5050 4748 5057 4751
rect 5146 4748 5153 4751
rect 1174 4738 1182 4741
rect 1270 4732 1273 4742
rect 1318 4738 1337 4741
rect 3778 4738 3785 4741
rect 1142 4728 1161 4731
rect 1334 4728 1337 4738
rect 1878 4728 1897 4731
rect 2022 4728 2025 4738
rect 2526 4728 2529 4738
rect 2534 4728 2553 4731
rect 3190 4728 3193 4738
rect 3286 4731 3290 4733
rect 3254 4728 3273 4731
rect 3278 4728 3290 4731
rect 3302 4732 3306 4736
rect 3758 4728 3777 4731
rect 4822 4728 4841 4731
rect 1197 4718 1198 4722
rect 1550 4718 1566 4721
rect 1709 4718 1710 4722
rect 3813 4718 3814 4722
rect 1048 4703 1050 4707
rect 1054 4703 1057 4707
rect 1061 4703 1064 4707
rect 2072 4703 2074 4707
rect 2078 4703 2081 4707
rect 2085 4703 2088 4707
rect 3096 4703 3098 4707
rect 3102 4703 3105 4707
rect 3109 4703 3112 4707
rect 4112 4703 4114 4707
rect 4118 4703 4121 4707
rect 4125 4703 4128 4707
rect 126 4671 129 4681
rect 406 4678 425 4681
rect 126 4668 145 4671
rect 442 4668 449 4671
rect 510 4668 518 4671
rect 746 4668 753 4671
rect 1166 4671 1169 4681
rect 1166 4668 1185 4671
rect 1222 4668 1241 4671
rect 1270 4671 1273 4681
rect 2030 4678 2049 4681
rect 2214 4678 2225 4681
rect 2742 4678 2761 4681
rect 2958 4678 2969 4681
rect 3158 4678 3177 4681
rect 3398 4678 3417 4681
rect 2214 4677 2218 4678
rect 2958 4677 2962 4678
rect 3422 4672 3425 4681
rect 1270 4668 1289 4671
rect 1562 4668 1577 4671
rect 1630 4668 1649 4671
rect 278 4658 297 4661
rect 342 4658 361 4661
rect 510 4658 529 4661
rect 658 4658 665 4661
rect 670 4658 678 4661
rect 1202 4658 1209 4661
rect 1294 4658 1302 4661
rect 1366 4658 1374 4661
rect 1590 4658 1598 4661
rect 1782 4658 1790 4661
rect 1958 4662 1961 4671
rect 2262 4668 2270 4671
rect 2318 4668 2326 4671
rect 2974 4668 2985 4671
rect 3618 4668 3641 4671
rect 2382 4658 2401 4661
rect 2542 4658 2561 4661
rect 2658 4658 2665 4661
rect 3018 4658 3025 4661
rect 3038 4658 3057 4661
rect 3398 4658 3401 4668
rect 3610 4658 3646 4661
rect 3654 4658 3673 4661
rect 3754 4658 3761 4661
rect 3958 4658 3974 4661
rect 4022 4658 4041 4661
rect 4326 4662 4329 4671
rect 4718 4668 4745 4671
rect 4454 4658 4473 4661
rect 4542 4658 4561 4661
rect 4630 4658 4638 4661
rect 4854 4658 4873 4661
rect 4946 4658 4953 4661
rect 4994 4658 5001 4661
rect 5038 4658 5054 4661
rect 5070 4658 5078 4661
rect 5138 4658 5145 4661
rect 278 4648 281 4658
rect 342 4648 345 4658
rect 510 4648 513 4658
rect 858 4648 862 4652
rect 1810 4648 1814 4652
rect 1938 4648 1942 4652
rect 2398 4648 2401 4658
rect 2558 4648 2561 4658
rect 3038 4648 3041 4658
rect 3278 4652 3282 4657
rect 3062 4648 3073 4651
rect 3082 4648 3086 4652
rect 3670 4648 3673 4658
rect 4038 4648 4041 4658
rect 4470 4648 4473 4658
rect 4542 4648 4545 4658
rect 4658 4648 4665 4651
rect 4766 4648 4785 4651
rect 4854 4648 4857 4658
rect 3062 4642 3065 4648
rect 266 4638 267 4642
rect 2843 4638 2846 4642
rect 2994 4638 2995 4642
rect 3515 4638 3518 4642
rect 3925 4638 3926 4642
rect 4149 4638 4150 4642
rect 4309 4638 4310 4642
rect 4373 4638 4374 4642
rect 4426 4638 4433 4641
rect 1314 4618 1315 4622
rect 3026 4618 3027 4622
rect 3605 4618 3606 4622
rect 4709 4618 4710 4622
rect 4813 4618 4814 4622
rect 536 4603 538 4607
rect 542 4603 545 4607
rect 549 4603 552 4607
rect 1560 4603 1562 4607
rect 1566 4603 1569 4607
rect 1573 4603 1576 4607
rect 2584 4603 2586 4607
rect 2590 4603 2593 4607
rect 2597 4603 2600 4607
rect 3608 4603 3610 4607
rect 3614 4603 3617 4607
rect 3621 4603 3624 4607
rect 4632 4603 4634 4607
rect 4638 4603 4641 4607
rect 4645 4603 4648 4607
rect 669 4588 670 4592
rect 1445 4588 1446 4592
rect 1605 4588 1606 4592
rect 3034 4588 3035 4592
rect 5077 4588 5078 4592
rect 282 4568 283 4572
rect 939 4568 942 4572
rect 1206 4568 1217 4571
rect 1214 4562 1217 4568
rect 1958 4568 1966 4571
rect 2230 4568 2238 4571
rect 2734 4568 2745 4571
rect 3747 4568 3750 4572
rect 1422 4566 1426 4568
rect 4078 4566 4082 4568
rect 4246 4566 4250 4568
rect 4382 4568 4390 4571
rect 4402 4568 4409 4571
rect 4286 4566 4290 4568
rect 4414 4566 4418 4568
rect 4470 4566 4474 4568
rect 4558 4566 4562 4568
rect 4582 4566 4586 4568
rect 4734 4566 4738 4568
rect 294 4551 297 4561
rect 294 4548 313 4551
rect 358 4551 361 4561
rect 342 4548 361 4551
rect 774 4551 777 4561
rect 758 4548 777 4551
rect 838 4551 841 4561
rect 1422 4558 1433 4561
rect 1930 4558 1934 4562
rect 2466 4558 2470 4562
rect 822 4548 841 4551
rect 1034 4548 1049 4551
rect 1286 4548 1294 4551
rect 2478 4551 2481 4561
rect 2558 4558 2566 4561
rect 2722 4558 2726 4562
rect 2478 4548 2497 4551
rect 2530 4548 2545 4551
rect 14 4538 33 4541
rect 262 4538 273 4541
rect 1366 4538 1374 4541
rect 1646 4538 1665 4541
rect 1778 4538 1785 4541
rect 1802 4538 1809 4541
rect 2106 4538 2121 4541
rect 2214 4538 2222 4541
rect 2454 4538 2457 4548
rect 2694 4548 2702 4551
rect 2714 4548 2721 4551
rect 3046 4551 3049 4561
rect 3550 4553 3554 4558
rect 3046 4548 3065 4551
rect 3070 4548 3078 4551
rect 3322 4548 3329 4551
rect 3642 4548 3657 4551
rect 3890 4548 3897 4551
rect 3950 4551 3953 4561
rect 4006 4558 4014 4561
rect 4054 4558 4073 4561
rect 3934 4548 3953 4551
rect 3986 4548 3993 4551
rect 3998 4548 4006 4551
rect 4090 4548 4097 4551
rect 4254 4551 4257 4561
rect 4522 4558 4526 4562
rect 4566 4558 4577 4561
rect 4566 4552 4569 4558
rect 4238 4548 4257 4551
rect 4306 4548 4313 4551
rect 4498 4548 4521 4551
rect 4538 4548 4553 4551
rect 4654 4548 4662 4551
rect 4842 4548 4849 4551
rect 4854 4548 4862 4551
rect 4902 4551 4905 4561
rect 4886 4548 4905 4551
rect 5062 4551 5065 4561
rect 5046 4548 5065 4551
rect 2558 4538 2574 4541
rect 3878 4538 3889 4541
rect 4022 4538 4033 4541
rect 30 4528 33 4538
rect 246 4531 250 4533
rect 246 4528 257 4531
rect 510 4528 529 4531
rect 534 4528 550 4531
rect 1374 4528 1393 4531
rect 1646 4528 1649 4538
rect 2150 4528 2158 4531
rect 2342 4528 2345 4538
rect 2926 4531 2930 4533
rect 2926 4528 2937 4531
rect 3134 4528 3153 4531
rect 3350 4528 3369 4531
rect 3862 4531 3866 4533
rect 4966 4532 4969 4542
rect 3862 4528 3873 4531
rect 4598 4528 4614 4531
rect 4730 4528 4734 4532
rect 725 4518 726 4522
rect 973 4518 974 4522
rect 1418 4518 1419 4522
rect 1562 4518 1577 4521
rect 2173 4518 2174 4522
rect 2522 4518 2523 4522
rect 2957 4518 2958 4522
rect 3010 4518 3011 4522
rect 3285 4518 3286 4522
rect 4610 4518 4625 4521
rect 5173 4518 5174 4522
rect 1048 4503 1050 4507
rect 1054 4503 1057 4507
rect 1061 4503 1064 4507
rect 2072 4503 2074 4507
rect 2078 4503 2081 4507
rect 2085 4503 2088 4507
rect 3096 4503 3098 4507
rect 3102 4503 3105 4507
rect 3109 4503 3112 4507
rect 4112 4503 4114 4507
rect 4118 4503 4121 4507
rect 4125 4503 4128 4507
rect 1610 4488 1611 4492
rect 4066 4488 4067 4492
rect 126 4478 145 4481
rect 390 4478 409 4481
rect 1334 4478 1345 4481
rect 1758 4478 1766 4481
rect 2838 4478 2850 4481
rect 3294 4478 3306 4481
rect 3610 4478 3625 4481
rect 3946 4478 3954 4481
rect 214 4468 217 4478
rect 1334 4477 1338 4478
rect 2846 4477 2850 4478
rect 3302 4477 3306 4478
rect 3950 4477 3954 4478
rect 5078 4472 5081 4481
rect 410 4468 417 4471
rect 1018 4468 1025 4471
rect 494 4458 502 4461
rect 894 4458 913 4461
rect 986 4458 993 4461
rect 998 4458 1014 4461
rect 1118 4458 1137 4461
rect 1150 4458 1166 4461
rect 1198 4458 1217 4461
rect 1298 4458 1305 4461
rect 1462 4458 1489 4461
rect 1626 4458 1633 4461
rect 1790 4458 1798 4461
rect 1878 4458 1905 4461
rect 1982 4458 1990 4461
rect 2486 4462 2489 4471
rect 2510 4468 2518 4471
rect 3142 4468 3153 4471
rect 3246 4468 3254 4471
rect 3810 4468 3817 4471
rect 4110 4468 4118 4471
rect 4130 4468 4142 4471
rect 4766 4468 4777 4471
rect 4874 4468 4881 4471
rect 5066 4468 5073 4471
rect 2318 4458 2337 4461
rect 2710 4458 2729 4461
rect 2750 4458 2769 4461
rect 2782 4458 2790 4461
rect 3206 4458 3225 4461
rect 3282 4458 3289 4461
rect 3526 4458 3534 4461
rect 3558 4458 3577 4461
rect 3590 4458 3598 4461
rect 3786 4458 3793 4461
rect 3802 4458 3825 4461
rect 3830 4458 3849 4461
rect 3894 4458 3902 4461
rect 4002 4458 4009 4461
rect 4274 4458 4281 4461
rect 4286 4458 4294 4461
rect 4422 4458 4441 4461
rect 4486 4458 4505 4461
rect 4558 4458 4566 4461
rect 4894 4458 4913 4461
rect 4926 4458 4934 4461
rect 4994 4458 5001 4461
rect 266 4448 270 4452
rect 750 4448 761 4451
rect 894 4448 897 4458
rect 1134 4448 1137 4458
rect 1214 4448 1217 4458
rect 1830 4448 1838 4451
rect 1982 4448 1985 4458
rect 2318 4448 2321 4458
rect 2410 4448 2414 4452
rect 2710 4448 2713 4458
rect 2766 4448 2769 4458
rect 3222 4448 3225 4458
rect 3234 4448 3238 4452
rect 3502 4448 3505 4458
rect 3574 4448 3577 4458
rect 3846 4448 3849 4458
rect 4262 4451 4266 4454
rect 4262 4448 4273 4451
rect 4422 4448 4425 4458
rect 4486 4448 4489 4458
rect 4690 4448 4694 4452
rect 4910 4448 4913 4458
rect 4922 4448 4926 4452
rect 5050 4448 5054 4452
rect 750 4442 754 4444
rect 675 4438 678 4442
rect 1723 4438 1726 4442
rect 2390 4441 2393 4448
rect 2390 4438 2402 4441
rect 2477 4438 2478 4442
rect 2566 4438 2574 4441
rect 3589 4438 3590 4442
rect 3934 4438 3942 4441
rect 3970 4438 3973 4442
rect 4371 4438 4374 4442
rect 4410 4438 4411 4442
rect 4826 4438 4833 4441
rect 882 4428 883 4432
rect 2306 4428 2307 4432
rect 2954 4428 2955 4432
rect 550 4418 566 4421
rect 714 4418 715 4422
rect 1789 4418 1790 4422
rect 1866 4418 1867 4422
rect 2365 4418 2366 4422
rect 2698 4418 2699 4422
rect 2986 4418 2987 4422
rect 3133 4418 3134 4422
rect 3266 4418 3267 4422
rect 3525 4418 3526 4422
rect 4757 4418 4758 4422
rect 536 4403 538 4407
rect 542 4403 545 4407
rect 549 4403 552 4407
rect 1560 4403 1562 4407
rect 1566 4403 1569 4407
rect 1573 4403 1576 4407
rect 2584 4403 2586 4407
rect 2590 4403 2593 4407
rect 2597 4403 2600 4407
rect 3608 4403 3610 4407
rect 3614 4403 3617 4407
rect 3621 4403 3624 4407
rect 4632 4403 4634 4407
rect 4638 4403 4641 4407
rect 4645 4403 4648 4407
rect 1029 4388 1030 4392
rect 1698 4388 1699 4392
rect 2066 4388 2067 4392
rect 4101 4388 4102 4392
rect 1446 4368 1458 4371
rect 1469 4368 1470 4372
rect 2003 4368 2006 4372
rect 2114 4368 2115 4372
rect 2126 4368 2137 4371
rect 3086 4368 3114 4371
rect 198 4358 217 4361
rect 286 4351 289 4361
rect 578 4358 582 4362
rect 286 4348 305 4351
rect 374 4348 382 4351
rect 590 4351 593 4361
rect 766 4361 769 4368
rect 758 4358 769 4361
rect 590 4348 609 4351
rect 618 4348 633 4351
rect 806 4351 809 4361
rect 990 4361 993 4368
rect 2134 4362 2137 4368
rect 3110 4366 3114 4368
rect 3326 4368 3337 4371
rect 3445 4368 3446 4372
rect 3606 4368 3622 4371
rect 3326 4366 3330 4368
rect 3606 4366 3610 4368
rect 3646 4366 3650 4368
rect 3670 4368 3681 4371
rect 3670 4366 3674 4368
rect 3790 4366 3794 4368
rect 4022 4368 4033 4371
rect 4022 4366 4026 4368
rect 4030 4362 4033 4368
rect 4046 4366 4050 4368
rect 4342 4366 4346 4368
rect 982 4358 993 4361
rect 778 4348 785 4351
rect 790 4348 809 4351
rect 974 4348 982 4351
rect 14 4338 33 4341
rect 238 4338 257 4341
rect 546 4338 569 4341
rect 1486 4338 1489 4348
rect 1678 4348 1686 4351
rect 1838 4351 1841 4361
rect 2022 4358 2033 4361
rect 2022 4356 2026 4358
rect 2150 4352 2153 4361
rect 2870 4358 2878 4361
rect 3146 4358 3150 4362
rect 3350 4353 3354 4358
rect 1838 4348 1857 4351
rect 1862 4348 1870 4351
rect 2090 4348 2110 4351
rect 2154 4348 2169 4351
rect 2482 4348 2489 4351
rect 2766 4348 2774 4351
rect 3030 4348 3046 4351
rect 3546 4348 3553 4351
rect 1510 4338 1518 4341
rect 1658 4338 1665 4341
rect 1682 4338 1689 4341
rect 1770 4338 1771 4342
rect 2098 4338 2105 4341
rect 2302 4338 2314 4341
rect 2594 4338 2610 4341
rect 2722 4338 2737 4341
rect 2806 4338 2825 4341
rect 2990 4338 3002 4341
rect 3158 4338 3166 4341
rect 30 4328 33 4338
rect 534 4328 553 4331
rect 1630 4328 1633 4338
rect 1638 4328 1657 4331
rect 2214 4331 2218 4333
rect 2206 4328 2218 4331
rect 2534 4328 2553 4331
rect 2822 4328 2825 4338
rect 3078 4336 3082 4338
rect 3214 4331 3218 4333
rect 3206 4328 3218 4331
rect 3366 4332 3369 4342
rect 3462 4338 3465 4348
rect 3918 4351 3921 4361
rect 4382 4358 4390 4361
rect 3898 4348 3905 4351
rect 3918 4348 3937 4351
rect 4138 4348 4145 4351
rect 4150 4348 4158 4351
rect 4582 4351 4585 4361
rect 4738 4358 4742 4362
rect 4566 4348 4585 4351
rect 4842 4348 4854 4351
rect 4886 4351 4889 4361
rect 4898 4358 4902 4362
rect 4870 4348 4889 4351
rect 5062 4351 5065 4361
rect 5046 4348 5065 4351
rect 3717 4338 3718 4342
rect 3990 4338 3998 4341
rect 4070 4338 4078 4341
rect 4110 4338 4118 4341
rect 4290 4338 4297 4341
rect 4374 4338 4385 4341
rect 4606 4338 4622 4341
rect 4758 4338 4761 4348
rect 4398 4331 4402 4333
rect 4390 4328 4402 4331
rect 325 4318 326 4322
rect 534 4321 537 4328
rect 526 4318 537 4321
rect 845 4318 846 4322
rect 1917 4318 1918 4322
rect 2037 4318 2038 4322
rect 2578 4318 2579 4322
rect 2714 4318 2715 4322
rect 3117 4318 3118 4322
rect 3602 4318 3603 4322
rect 3642 4318 3643 4322
rect 3666 4318 3667 4322
rect 4018 4318 4019 4322
rect 4042 4318 4043 4322
rect 4338 4318 4339 4322
rect 1048 4303 1050 4307
rect 1054 4303 1057 4307
rect 1061 4303 1064 4307
rect 2072 4303 2074 4307
rect 2078 4303 2081 4307
rect 2085 4303 2088 4307
rect 3096 4303 3098 4307
rect 3102 4303 3105 4307
rect 3109 4303 3112 4307
rect 4112 4303 4114 4307
rect 4118 4303 4121 4307
rect 4125 4303 4128 4307
rect 3098 4288 3099 4292
rect 3978 4288 3979 4292
rect 4213 4288 4214 4292
rect 30 4271 33 4281
rect 222 4278 233 4281
rect 342 4278 353 4281
rect 390 4278 409 4281
rect 702 4278 721 4281
rect 894 4278 913 4281
rect 1318 4278 1337 4281
rect 1926 4278 1937 4281
rect 222 4277 226 4278
rect 342 4277 346 4278
rect 1926 4277 1930 4278
rect 14 4268 33 4271
rect 422 4262 425 4271
rect 1258 4268 1262 4271
rect 1630 4268 1638 4271
rect 1942 4268 1953 4271
rect 2006 4271 2009 4281
rect 2726 4278 2745 4281
rect 3054 4278 3073 4281
rect 3294 4278 3305 4281
rect 4274 4278 4286 4281
rect 3294 4277 3298 4278
rect 2006 4268 2025 4271
rect 2230 4268 2241 4271
rect 2542 4268 2570 4271
rect 2926 4268 2953 4271
rect 3306 4268 3313 4271
rect 3502 4268 3513 4271
rect 166 4258 174 4261
rect 566 4258 585 4261
rect 1006 4258 1025 4261
rect 1038 4258 1054 4261
rect 2238 4262 2241 4268
rect 1250 4258 1273 4261
rect 1598 4258 1617 4261
rect 1622 4258 1646 4261
rect 1654 4258 1673 4261
rect 1870 4258 1878 4261
rect 1966 4258 1974 4261
rect 2030 4258 2038 4261
rect 2262 4258 2270 4261
rect 2898 4258 2905 4261
rect 3354 4258 3361 4261
rect 3510 4262 3513 4268
rect 3574 4262 3577 4271
rect 3598 4268 3606 4271
rect 3814 4262 3817 4271
rect 3862 4268 3870 4271
rect 3962 4268 3969 4271
rect 4174 4268 4182 4271
rect 4230 4262 4233 4271
rect 4310 4271 4313 4281
rect 4294 4268 4313 4271
rect 4446 4268 4454 4271
rect 4458 4268 4465 4271
rect 4638 4268 4665 4271
rect 4054 4258 4062 4261
rect 4502 4258 4510 4261
rect 4570 4258 4577 4261
rect 4814 4258 4833 4261
rect 4974 4258 4993 4261
rect 5074 4258 5081 4261
rect 566 4248 569 4258
rect 774 4248 793 4251
rect 1022 4248 1025 4258
rect 1034 4248 1038 4252
rect 1166 4251 1169 4258
rect 1166 4248 1177 4251
rect 1206 4251 1209 4258
rect 1206 4248 1217 4251
rect 1222 4248 1233 4251
rect 1598 4248 1601 4258
rect 1670 4248 1673 4258
rect 1682 4248 1686 4252
rect 2902 4248 2905 4258
rect 2914 4248 2918 4252
rect 3122 4248 3129 4251
rect 3138 4248 3142 4252
rect 3878 4248 3889 4251
rect 3894 4248 3902 4251
rect 4682 4248 4689 4251
rect 4694 4248 4697 4258
rect 4830 4248 4833 4258
rect 4990 4248 4993 4258
rect 1222 4242 1225 4248
rect 3878 4242 3881 4248
rect 1419 4238 1422 4242
rect 4882 4238 4885 4242
rect 5005 4238 5006 4242
rect 554 4218 555 4222
rect 2189 4218 2190 4222
rect 2261 4218 2262 4222
rect 2362 4218 2363 4222
rect 2874 4218 2875 4222
rect 3178 4218 3179 4222
rect 3549 4218 3550 4222
rect 3794 4218 3795 4222
rect 4021 4218 4022 4222
rect 4053 4218 4054 4222
rect 4154 4218 4155 4222
rect 4629 4218 4630 4222
rect 536 4203 538 4207
rect 542 4203 545 4207
rect 549 4203 552 4207
rect 1560 4203 1562 4207
rect 1566 4203 1569 4207
rect 1573 4203 1576 4207
rect 2584 4203 2586 4207
rect 2590 4203 2593 4207
rect 2597 4203 2600 4207
rect 3608 4203 3610 4207
rect 3614 4203 3617 4207
rect 3621 4203 3624 4207
rect 4632 4203 4634 4207
rect 4638 4203 4641 4207
rect 4645 4203 4648 4207
rect 786 4188 787 4192
rect 1378 4188 1379 4192
rect 2346 4188 2347 4192
rect 2730 4188 2731 4192
rect 4498 4188 4499 4192
rect 1330 4178 1331 4182
rect 2314 4178 2315 4182
rect 1226 4168 1234 4171
rect 2026 4168 2029 4172
rect 3434 4168 3435 4172
rect 3965 4168 3966 4172
rect 4090 4168 4097 4171
rect 4205 4168 4206 4172
rect 5058 4168 5059 4172
rect 3286 4166 3290 4168
rect 3558 4166 3562 4168
rect 3782 4166 3786 4168
rect 3998 4166 4002 4168
rect 4462 4166 4466 4168
rect 206 4148 214 4151
rect 238 4151 241 4161
rect 238 4148 257 4151
rect 318 4151 321 4161
rect 390 4158 409 4161
rect 418 4158 422 4162
rect 510 4158 518 4161
rect 318 4148 337 4151
rect 442 4148 449 4151
rect 502 4148 529 4151
rect 662 4148 670 4151
rect 798 4151 801 4161
rect 1186 4158 1190 4162
rect 798 4148 817 4151
rect 862 4148 878 4151
rect 1226 4148 1241 4151
rect 1286 4151 1289 4161
rect 1270 4148 1289 4151
rect 1334 4148 1342 4151
rect 1526 4148 1545 4151
rect 1550 4148 1558 4151
rect 1562 4148 1582 4151
rect 1622 4151 1625 4161
rect 1714 4158 1718 4162
rect 1622 4148 1641 4151
rect 526 4142 529 4148
rect 1526 4142 1529 4148
rect 1902 4148 1910 4151
rect 1974 4151 1977 4161
rect 1986 4158 1990 4162
rect 2114 4158 2121 4161
rect 2282 4158 2286 4162
rect 1958 4148 1977 4151
rect 2158 4148 2166 4151
rect 2538 4148 2553 4151
rect 2622 4148 2649 4151
rect 2742 4151 2745 4161
rect 3262 4158 3281 4161
rect 3746 4158 3750 4162
rect 3782 4158 3793 4161
rect 3846 4158 3858 4161
rect 3854 4156 3858 4158
rect 2742 4148 2761 4151
rect 206 4138 217 4141
rect 622 4138 634 4141
rect 770 4138 777 4141
rect 1558 4138 1601 4141
rect 1622 4138 1630 4141
rect 2094 4138 2102 4141
rect 2122 4138 2129 4141
rect 2714 4138 2721 4141
rect 2862 4138 2865 4148
rect 3806 4148 3830 4151
rect 3838 4148 3846 4151
rect 3886 4148 3894 4151
rect 2886 4138 2913 4141
rect 2981 4138 2982 4142
rect 3066 4138 3078 4141
rect 3094 4138 3129 4141
rect 3462 4138 3481 4141
rect 3782 4141 3785 4148
rect 3966 4148 3974 4151
rect 4226 4148 4233 4151
rect 4306 4148 4313 4151
rect 4374 4142 4377 4151
rect 4430 4151 4433 4161
rect 4414 4148 4433 4151
rect 4482 4148 4497 4151
rect 4690 4148 4697 4151
rect 4918 4151 4921 4161
rect 4930 4158 4934 4162
rect 4902 4148 4921 4151
rect 3782 4138 3793 4141
rect 4070 4138 4078 4141
rect 4293 4138 4294 4142
rect 190 4131 194 4133
rect 718 4131 722 4133
rect 190 4128 201 4131
rect 718 4128 729 4131
rect 1570 4128 1585 4131
rect 1862 4128 1881 4131
rect 2174 4131 2178 4133
rect 2166 4128 2178 4131
rect 2366 4132 2369 4138
rect 2366 4128 2374 4132
rect 2446 4128 2465 4131
rect 3094 4128 3097 4138
rect 3478 4128 3481 4138
rect 4374 4128 4393 4131
rect 277 4118 278 4122
rect 461 4118 462 4122
rect 850 4118 851 4122
rect 1213 4118 1214 4122
rect 1741 4118 1742 4122
rect 2413 4118 2414 4122
rect 3573 4118 3574 4122
rect 3778 4118 3779 4122
rect 3994 4118 3995 4122
rect 1048 4103 1050 4107
rect 1054 4103 1057 4107
rect 1061 4103 1064 4107
rect 2072 4103 2074 4107
rect 2078 4103 2081 4107
rect 2085 4103 2088 4107
rect 3096 4103 3098 4107
rect 3102 4103 3105 4107
rect 3109 4103 3112 4107
rect 4112 4103 4114 4107
rect 4118 4103 4121 4107
rect 4125 4103 4128 4107
rect 1973 4088 1974 4092
rect 3322 4088 3323 4092
rect 4074 4088 4075 4092
rect 5077 4088 5078 4092
rect 126 4078 145 4081
rect 246 4078 257 4081
rect 1358 4078 1369 4081
rect 246 4077 250 4078
rect 1358 4077 1362 4078
rect 118 4068 126 4071
rect 262 4068 273 4071
rect 582 4068 590 4071
rect 670 4068 678 4071
rect 898 4068 905 4071
rect 1126 4062 1129 4071
rect 1262 4062 1265 4071
rect 1498 4068 1505 4071
rect 1858 4068 1865 4071
rect 2110 4068 2118 4071
rect 2274 4068 2281 4071
rect 2582 4071 2585 4078
rect 2582 4068 2593 4071
rect 3054 4071 3057 4081
rect 4606 4078 4641 4081
rect 4798 4078 4810 4081
rect 3038 4068 3057 4071
rect 3246 4068 3249 4078
rect 4806 4077 4810 4078
rect 3726 4068 3734 4071
rect 3838 4068 3854 4071
rect 3966 4068 3974 4071
rect 4174 4068 4182 4071
rect 4446 4068 4457 4071
rect 4790 4068 4798 4071
rect 274 4058 281 4061
rect 294 4058 313 4061
rect 406 4058 433 4061
rect 574 4058 582 4061
rect 594 4058 601 4061
rect 878 4058 886 4061
rect 890 4058 897 4061
rect 970 4058 977 4061
rect 1154 4058 1161 4061
rect 1194 4058 1201 4061
rect 1506 4058 1513 4061
rect 1570 4058 1585 4061
rect 1790 4058 1809 4061
rect 1838 4058 1865 4061
rect 1950 4058 1958 4061
rect 2006 4058 2014 4061
rect 2182 4058 2201 4061
rect 2650 4058 2657 4061
rect 4446 4062 4449 4068
rect 2778 4058 2785 4061
rect 2790 4058 2809 4061
rect 3358 4058 3377 4061
rect 3522 4058 3545 4061
rect 3582 4058 3617 4061
rect 3674 4058 3681 4061
rect 3878 4058 3886 4061
rect 4130 4058 4161 4061
rect 4206 4058 4225 4061
rect 4270 4058 4289 4061
rect 4774 4058 4782 4061
rect 282 4048 286 4052
rect 294 4048 297 4058
rect 486 4048 497 4051
rect 538 4048 561 4051
rect 570 4048 574 4052
rect 894 4048 897 4058
rect 1790 4048 1793 4058
rect 2182 4048 2185 4058
rect 2238 4048 2257 4051
rect 2806 4048 2809 4058
rect 2818 4048 2822 4052
rect 3358 4048 3361 4058
rect 3486 4048 3505 4051
rect 3614 4048 3617 4058
rect 4206 4048 4209 4058
rect 4286 4048 4289 4058
rect 4298 4048 4302 4052
rect 494 4042 497 4048
rect 227 4038 230 4042
rect 1253 4038 1254 4042
rect 2586 4038 2594 4041
rect 3098 4038 3105 4041
rect 3789 4038 3790 4042
rect 3517 4028 3518 4032
rect 3757 4028 3758 4032
rect 602 4018 603 4022
rect 989 4018 990 4022
rect 1202 4018 1203 4022
rect 1418 4018 1419 4022
rect 1597 4018 1598 4022
rect 1741 4018 1742 4022
rect 2226 4018 2227 4022
rect 2378 4018 2379 4022
rect 2658 4018 2659 4022
rect 3546 4018 3547 4022
rect 3629 4018 3630 4022
rect 3925 4018 3926 4022
rect 3997 4018 3998 4022
rect 4106 4018 4107 4022
rect 536 4003 538 4007
rect 542 4003 545 4007
rect 549 4003 552 4007
rect 1560 4003 1562 4007
rect 1566 4003 1569 4007
rect 1573 4003 1576 4007
rect 2584 4003 2586 4007
rect 2590 4003 2593 4007
rect 2597 4003 2600 4007
rect 3608 4003 3610 4007
rect 3614 4003 3617 4007
rect 3621 4003 3624 4007
rect 4632 4003 4634 4007
rect 4638 4003 4641 4007
rect 4645 4003 4648 4007
rect 1141 3988 1142 3992
rect 1658 3988 1659 3992
rect 2538 3988 2539 3992
rect 2757 3988 2758 3992
rect 4274 3988 4275 3992
rect 4397 3988 4398 3992
rect 4930 3988 4931 3992
rect 979 3968 982 3972
rect 1166 3968 1174 3971
rect 1690 3968 1691 3972
rect 2090 3968 2093 3972
rect 2357 3968 2358 3972
rect 2725 3968 2726 3972
rect 2786 3968 2787 3972
rect 2874 3968 2875 3972
rect 1710 3966 1714 3968
rect 3062 3966 3066 3968
rect 3374 3966 3378 3968
rect 4574 3966 4578 3968
rect 4662 3968 4670 3971
rect 4733 3968 4734 3972
rect 4970 3968 4973 3972
rect 4662 3966 4666 3968
rect 362 3958 366 3962
rect 454 3951 457 3961
rect 454 3948 473 3951
rect 870 3951 873 3961
rect 870 3948 889 3951
rect 942 3948 950 3951
rect 1046 3948 1062 3951
rect 1294 3948 1305 3951
rect 1478 3948 1486 3951
rect 1614 3951 1617 3961
rect 1702 3958 1713 3961
rect 1598 3948 1617 3951
rect 1630 3948 1654 3951
rect 1790 3951 1793 3961
rect 1730 3948 1737 3951
rect 1774 3948 1793 3951
rect 1866 3948 1873 3951
rect 1302 3942 1305 3948
rect 2026 3948 2033 3951
rect 2286 3951 2289 3961
rect 2706 3958 2713 3961
rect 3410 3958 3414 3962
rect 2270 3948 2289 3951
rect 2858 3948 2870 3951
rect 3066 3948 3081 3951
rect 3270 3951 3273 3958
rect 3262 3948 3273 3951
rect 3422 3951 3425 3961
rect 3578 3958 3582 3962
rect 3394 3948 3409 3951
rect 3422 3948 3441 3951
rect 3590 3951 3593 3961
rect 4106 3958 4113 3961
rect 4202 3958 4209 3961
rect 3590 3948 3609 3951
rect 4058 3948 4065 3951
rect 4286 3948 4313 3951
rect 4566 3951 4569 3961
rect 4594 3958 4601 3961
rect 4566 3948 4585 3951
rect 4718 3951 4721 3961
rect 4702 3948 4721 3951
rect 4902 3948 4918 3951
rect 5070 3951 5073 3961
rect 5070 3948 5089 3951
rect 5158 3951 5161 3961
rect 5142 3948 5161 3951
rect 118 3938 126 3941
rect 342 3938 353 3941
rect 410 3938 417 3941
rect 1150 3938 1158 3941
rect 1434 3938 1441 3941
rect 1750 3938 1758 3941
rect 1842 3938 1849 3941
rect 2158 3938 2170 3941
rect 2282 3938 2289 3941
rect 2310 3938 2329 3941
rect 2686 3938 2697 3941
rect 3006 3938 3014 3941
rect 3098 3938 3121 3941
rect 3246 3938 3254 3941
rect 3558 3938 3569 3941
rect 4138 3938 4145 3941
rect 4218 3938 4225 3941
rect 4378 3938 4401 3941
rect 4538 3938 4545 3941
rect 4742 3938 4753 3941
rect 5182 3938 5190 3941
rect 126 3928 145 3931
rect 182 3928 201 3931
rect 1102 3928 1105 3938
rect 1422 3931 1426 3933
rect 1422 3928 1433 3931
rect 1874 3928 1881 3931
rect 3134 3931 3138 3933
rect 3126 3928 3138 3931
rect 3278 3931 3282 3933
rect 3270 3928 3282 3931
rect 3542 3931 3546 3933
rect 3542 3928 3553 3931
rect 3958 3928 3977 3931
rect 4342 3928 4361 3931
rect 317 3918 318 3922
rect 389 3918 390 3922
rect 1834 3918 1835 3922
rect 1858 3918 1859 3922
rect 2402 3918 2403 3922
rect 2997 3918 2998 3922
rect 3058 3918 3059 3922
rect 4658 3918 4659 3922
rect 4682 3918 4683 3922
rect 1048 3903 1050 3907
rect 1054 3903 1057 3907
rect 1061 3903 1064 3907
rect 2072 3903 2074 3907
rect 2078 3903 2081 3907
rect 2085 3903 2088 3907
rect 3096 3903 3098 3907
rect 3102 3903 3105 3907
rect 3109 3903 3112 3907
rect 4112 3903 4114 3907
rect 4118 3903 4121 3907
rect 4125 3903 4128 3907
rect 3082 3888 3083 3892
rect 4118 3888 4134 3891
rect 4181 3888 4182 3892
rect 646 3878 657 3881
rect 758 3878 769 3881
rect 990 3878 1009 3881
rect 2118 3878 2137 3881
rect 2478 3878 2497 3881
rect 2846 3878 2858 3881
rect 646 3877 650 3878
rect 758 3877 762 3878
rect 2854 3877 2858 3878
rect 3198 3878 3209 3881
rect 3214 3878 3222 3881
rect 3198 3877 3202 3878
rect 206 3868 217 3871
rect 422 3868 433 3871
rect 1422 3868 1430 3871
rect 1718 3868 1729 3871
rect 2030 3868 2041 3871
rect 2170 3868 2177 3871
rect 2382 3868 2393 3871
rect 2522 3868 2537 3871
rect 2798 3868 2809 3871
rect 3286 3868 3305 3871
rect 3510 3871 3513 3881
rect 3982 3878 4001 3881
rect 4558 3878 4570 3881
rect 4566 3877 4570 3878
rect 3494 3868 3513 3871
rect 3678 3868 3697 3871
rect 3994 3868 4009 3871
rect 4605 3868 4606 3872
rect 4674 3868 4681 3871
rect 4742 3868 4753 3871
rect 5026 3868 5033 3871
rect 238 3858 257 3861
rect 590 3858 598 3861
rect 1006 3858 1009 3868
rect 1146 3858 1153 3861
rect 1158 3858 1166 3861
rect 1414 3858 1422 3861
rect 1426 3858 1433 3861
rect 1562 3858 1577 3861
rect 1678 3858 1705 3861
rect 1838 3858 1846 3861
rect 1870 3861 1873 3868
rect 1862 3858 1873 3861
rect 2062 3858 2097 3861
rect 2346 3858 2353 3861
rect 2454 3858 2462 3861
rect 3018 3858 3025 3861
rect 3162 3858 3169 3861
rect 3302 3861 3305 3868
rect 3302 3858 3313 3861
rect 3390 3858 3409 3861
rect 3642 3858 3665 3861
rect 3670 3858 3686 3861
rect 3750 3858 3758 3861
rect 3782 3858 3801 3861
rect 4214 3858 4233 3861
rect 4458 3858 4465 3861
rect 4502 3858 4521 3861
rect 4750 3861 4753 3868
rect 4750 3858 4766 3861
rect 4774 3858 4793 3861
rect 4838 3858 4857 3861
rect 4918 3858 4926 3861
rect 4938 3858 4945 3861
rect 5018 3858 5041 3861
rect 5046 3858 5065 3861
rect 226 3848 230 3852
rect 238 3848 241 3858
rect 1346 3848 1350 3852
rect 1430 3848 1433 3858
rect 1438 3848 1446 3851
rect 2062 3848 2065 3858
rect 2354 3848 2358 3852
rect 2366 3848 2374 3851
rect 2766 3848 2777 3851
rect 3038 3848 3057 3851
rect 3062 3848 3073 3851
rect 3406 3848 3409 3858
rect 3798 3848 3801 3858
rect 4166 3848 4177 3851
rect 4230 3848 4233 3858
rect 4242 3848 4246 3852
rect 4518 3848 4521 3858
rect 4790 3848 4793 3858
rect 4854 3848 4857 3858
rect 5062 3848 5065 3858
rect 5074 3848 5078 3852
rect 2766 3842 2769 3848
rect 3070 3842 3073 3848
rect 3230 3842 3234 3844
rect 3246 3841 3249 3848
rect 3238 3838 3249 3841
rect 3630 3838 3658 3841
rect 2442 3828 2443 3832
rect 378 3818 379 3822
rect 413 3818 414 3822
rect 534 3818 550 3821
rect 805 3818 806 3822
rect 1666 3818 1667 3822
rect 1802 3818 1803 3822
rect 2709 3818 2710 3822
rect 2818 3818 2819 3822
rect 3026 3818 3027 3822
rect 3325 3818 3326 3822
rect 3365 3818 3366 3822
rect 3853 3818 3854 3822
rect 4154 3818 4155 3822
rect 4805 3818 4806 3822
rect 5013 3818 5014 3822
rect 536 3803 538 3807
rect 542 3803 545 3807
rect 549 3803 552 3807
rect 1560 3803 1562 3807
rect 1566 3803 1569 3807
rect 1573 3803 1576 3807
rect 2584 3803 2586 3807
rect 2590 3803 2593 3807
rect 2597 3803 2600 3807
rect 3608 3803 3610 3807
rect 3614 3803 3617 3807
rect 3621 3803 3624 3807
rect 4632 3803 4634 3807
rect 4638 3803 4641 3807
rect 4645 3803 4648 3807
rect 690 3788 691 3792
rect 1002 3788 1003 3792
rect 1749 3788 1750 3792
rect 2658 3788 2659 3792
rect 3413 3788 3414 3792
rect 410 3778 411 3782
rect 2394 3768 2395 3772
rect 2938 3768 2941 3772
rect 3342 3768 3354 3771
rect 3350 3766 3354 3768
rect 4178 3768 4181 3772
rect 3646 3766 3650 3768
rect 3950 3766 3954 3768
rect 4366 3766 4370 3768
rect 4454 3768 4465 3771
rect 4454 3766 4458 3768
rect 4622 3766 4626 3768
rect 4750 3766 4754 3768
rect 350 3758 369 3761
rect 50 3748 65 3751
rect 422 3751 425 3761
rect 422 3748 441 3751
rect 486 3748 502 3751
rect 702 3751 705 3761
rect 702 3748 721 3751
rect 926 3751 929 3761
rect 926 3748 945 3751
rect 1046 3751 1049 3761
rect 1066 3758 1073 3761
rect 1046 3748 1081 3751
rect 1086 3748 1102 3751
rect 1118 3751 1121 3761
rect 1118 3748 1126 3751
rect 1334 3751 1337 3761
rect 1318 3748 1337 3751
rect 1638 3751 1641 3761
rect 1774 3758 1793 3761
rect 1638 3748 1657 3751
rect 1902 3751 1905 3761
rect 2166 3753 2170 3758
rect 1886 3748 1905 3751
rect 94 3738 106 3741
rect 646 3738 654 3741
rect 1086 3738 1089 3748
rect 2214 3742 2217 3751
rect 2406 3751 2409 3761
rect 2582 3758 2590 3761
rect 2386 3748 2393 3751
rect 2406 3748 2425 3751
rect 2522 3748 2529 3751
rect 2670 3751 2673 3761
rect 3638 3758 3649 3761
rect 3674 3758 3681 3761
rect 3326 3753 3330 3758
rect 2670 3748 2689 3751
rect 2714 3748 2721 3751
rect 3606 3748 3614 3751
rect 3870 3748 3889 3751
rect 4130 3748 4137 3751
rect 4210 3748 4217 3751
rect 4358 3751 4361 3761
rect 4734 3758 4745 3761
rect 4734 3752 4737 3758
rect 4358 3748 4377 3751
rect 4446 3748 4454 3751
rect 1606 3738 1617 3741
rect 1662 3738 1670 3741
rect 1758 3738 1766 3741
rect 1814 3738 1822 3741
rect 2594 3738 2606 3741
rect 2870 3738 2889 3741
rect 3078 3738 3086 3741
rect 3690 3738 3697 3741
rect 4078 3741 4081 3748
rect 4070 3738 4081 3741
rect 4150 3738 4153 3748
rect 4706 3748 4713 3751
rect 4818 3748 4833 3751
rect 4970 3748 4977 3751
rect 4982 3748 4990 3751
rect 5042 3748 5057 3751
rect 4298 3738 4305 3741
rect 4394 3738 4401 3741
rect 4558 3741 4561 3748
rect 4558 3738 4569 3741
rect 4654 3738 4673 3741
rect 4750 3741 4753 3748
rect 4750 3738 4761 3741
rect 4862 3738 4874 3741
rect 190 3731 194 3733
rect 1198 3732 1202 3736
rect 190 3728 201 3731
rect 562 3728 569 3731
rect 1582 3728 1601 3731
rect 2182 3731 2186 3733
rect 2286 3731 2290 3733
rect 2182 3728 2193 3731
rect 2198 3728 2217 3731
rect 2278 3728 2290 3731
rect 2886 3728 2889 3738
rect 3222 3728 3241 3731
rect 4670 3728 4673 3738
rect 4782 3736 4786 3738
rect 661 3718 662 3722
rect 757 3718 758 3722
rect 1133 3718 1134 3722
rect 1290 3718 1291 3722
rect 1469 3718 1470 3722
rect 1582 3721 1585 3728
rect 1574 3718 1585 3721
rect 1845 3718 1846 3722
rect 2042 3718 2043 3722
rect 2066 3718 2067 3722
rect 3653 3718 3654 3722
rect 4274 3718 4275 3722
rect 4622 3718 4630 3721
rect 1048 3703 1050 3707
rect 1054 3703 1057 3707
rect 1061 3703 1064 3707
rect 2072 3703 2074 3707
rect 2078 3703 2081 3707
rect 2085 3703 2088 3707
rect 3096 3703 3098 3707
rect 3102 3703 3105 3707
rect 3109 3703 3112 3707
rect 4112 3703 4114 3707
rect 4118 3703 4121 3707
rect 4125 3703 4128 3707
rect 2046 3688 2057 3691
rect 14 3678 33 3681
rect 246 3678 265 3681
rect 614 3678 625 3681
rect 614 3677 618 3678
rect 854 3672 857 3681
rect 965 3678 966 3682
rect 446 3668 457 3671
rect 1046 3671 1049 3681
rect 1821 3678 1822 3682
rect 2046 3681 2049 3688
rect 2574 3681 2577 3688
rect 2030 3678 2049 3681
rect 2494 3678 2505 3681
rect 2574 3678 2593 3681
rect 2662 3678 2674 3681
rect 2494 3677 2498 3678
rect 2670 3677 2674 3678
rect 3054 3678 3065 3681
rect 3102 3678 3137 3681
rect 3054 3677 3058 3678
rect 862 3668 873 3671
rect 1046 3668 1081 3671
rect 1158 3668 1166 3671
rect 1926 3668 1934 3671
rect 1982 3668 1993 3671
rect 2014 3668 2025 3671
rect 2330 3668 2337 3671
rect 446 3662 449 3668
rect 182 3658 201 3661
rect 470 3658 478 3661
rect 630 3658 638 3661
rect 886 3658 894 3661
rect 954 3658 961 3661
rect 1126 3658 1134 3661
rect 1154 3658 1177 3661
rect 1182 3658 1201 3661
rect 1982 3662 1985 3668
rect 1482 3658 1489 3661
rect 1502 3658 1510 3661
rect 1534 3658 1569 3661
rect 1586 3658 1598 3661
rect 1794 3658 1809 3661
rect 1878 3658 1886 3661
rect 2542 3662 2545 3671
rect 2654 3668 2662 3671
rect 3422 3671 3425 3681
rect 3806 3678 3825 3681
rect 4230 3678 4249 3681
rect 4518 3678 4530 3681
rect 4526 3677 4530 3678
rect 3422 3668 3441 3671
rect 3850 3668 3865 3671
rect 3922 3668 3929 3671
rect 4502 3668 4513 3671
rect 4658 3668 4665 3671
rect 4750 3668 4753 3678
rect 4862 3668 4870 3671
rect 4894 3671 4897 3681
rect 4878 3668 4897 3671
rect 5046 3671 5049 3681
rect 5142 3678 5161 3681
rect 5046 3668 5065 3671
rect 2174 3658 2193 3661
rect 2522 3658 2529 3661
rect 2554 3658 2561 3661
rect 2722 3658 2729 3661
rect 2802 3658 2809 3661
rect 2906 3658 2913 3661
rect 2918 3658 2937 3661
rect 3066 3658 3073 3661
rect 3526 3658 3545 3661
rect 3634 3658 3646 3661
rect 3654 3658 3673 3661
rect 3734 3658 3742 3661
rect 3846 3658 3854 3661
rect 3946 3658 3953 3661
rect 3966 3658 3985 3661
rect 4058 3658 4065 3661
rect 4070 3658 4094 3661
rect 4322 3658 4337 3661
rect 4462 3658 4481 3661
rect 4654 3658 4662 3661
rect 5182 3658 5190 3661
rect 182 3648 185 3658
rect 678 3648 697 3651
rect 1126 3648 1129 3658
rect 1198 3648 1201 3658
rect 1486 3648 1489 3658
rect 1542 3648 1558 3651
rect 1566 3648 1569 3658
rect 2174 3648 2177 3658
rect 2686 3652 2690 3657
rect 2586 3648 2593 3651
rect 2778 3648 2782 3652
rect 2934 3648 2937 3658
rect 3038 3652 3042 3657
rect 2946 3648 2950 3652
rect 3270 3648 3289 3651
rect 3526 3648 3529 3658
rect 3670 3648 3673 3658
rect 3966 3648 3969 3658
rect 4478 3648 4481 3658
rect 4490 3648 4494 3652
rect 4654 3651 4657 3658
rect 4638 3648 4657 3651
rect 4694 3648 4697 3658
rect 4818 3648 4825 3651
rect 5102 3648 5121 3651
rect 1614 3641 1618 3644
rect 5126 3642 5130 3644
rect 1614 3638 1625 3641
rect 3685 3638 3686 3642
rect 4122 3638 4125 3642
rect 4546 3638 4549 3642
rect 4702 3638 4710 3641
rect 4946 3638 4949 3642
rect 1213 3628 1214 3632
rect 421 3618 422 3622
rect 650 3618 651 3622
rect 709 3618 710 3622
rect 1149 3618 1150 3622
rect 1501 3618 1502 3622
rect 1581 3618 1582 3622
rect 4026 3618 4027 3622
rect 4426 3618 4427 3622
rect 4853 3618 4854 3622
rect 536 3603 538 3607
rect 542 3603 545 3607
rect 549 3603 552 3607
rect 1560 3603 1562 3607
rect 1566 3603 1569 3607
rect 1573 3603 1576 3607
rect 2584 3603 2586 3607
rect 2590 3603 2593 3607
rect 2597 3603 2600 3607
rect 3608 3603 3610 3607
rect 3614 3603 3617 3607
rect 3621 3603 3624 3607
rect 4632 3603 4634 3607
rect 4638 3603 4641 3607
rect 4645 3603 4648 3607
rect 605 3588 606 3592
rect 2458 3588 2459 3592
rect 3434 3588 3435 3592
rect 4725 3588 4726 3592
rect 2714 3578 2715 3582
rect 147 3568 150 3572
rect 243 3568 246 3572
rect 317 3568 318 3572
rect 1138 3568 1139 3572
rect 2494 3568 2505 3571
rect 3285 3568 3286 3572
rect 2494 3566 2498 3568
rect 3398 3566 3402 3568
rect 3774 3566 3778 3568
rect 4978 3568 4981 3572
rect 3974 3566 3978 3568
rect 5054 3566 5058 3568
rect 302 3552 305 3561
rect 342 3558 350 3561
rect 286 3548 294 3551
rect 590 3551 593 3561
rect 882 3558 886 3562
rect 574 3548 593 3551
rect 894 3551 897 3561
rect 894 3548 913 3551
rect 1006 3548 1022 3551
rect 1062 3548 1078 3551
rect 1366 3548 1374 3551
rect 1462 3551 1465 3561
rect 1818 3558 1822 3562
rect 1446 3548 1465 3551
rect 1614 3548 1622 3551
rect 1830 3551 1833 3561
rect 1830 3548 1849 3551
rect 1990 3551 1993 3561
rect 2070 3558 2105 3561
rect 2110 3558 2121 3561
rect 2130 3558 2134 3562
rect 1990 3548 2009 3551
rect 2154 3548 2161 3551
rect 2398 3551 2401 3561
rect 2470 3558 2489 3561
rect 2874 3558 2878 3562
rect 3150 3558 3162 3561
rect 3158 3556 3162 3558
rect 2382 3548 2401 3551
rect 2846 3548 2854 3551
rect 3014 3548 3022 3551
rect 3142 3548 3150 3551
rect 382 3538 393 3541
rect 662 3538 673 3541
rect 862 3538 873 3541
rect 1582 3538 1590 3541
rect 2022 3538 2030 3541
rect 2038 3538 2049 3541
rect 2221 3538 2222 3542
rect 2422 3538 2449 3541
rect 3006 3541 3009 3548
rect 3446 3551 3449 3561
rect 3502 3551 3505 3561
rect 3418 3548 3433 3551
rect 3446 3548 3465 3551
rect 3486 3548 3505 3551
rect 3518 3548 3526 3551
rect 3686 3551 3689 3561
rect 3906 3558 3910 3562
rect 3658 3548 3673 3551
rect 3686 3548 3705 3551
rect 3710 3548 3729 3551
rect 2998 3538 3009 3541
rect 3106 3538 3126 3541
rect 3294 3538 3302 3541
rect 3362 3538 3377 3541
rect 3526 3538 3537 3541
rect 3726 3541 3729 3548
rect 3726 3538 3737 3541
rect 3790 3541 3793 3548
rect 4166 3551 4169 3561
rect 4178 3558 4182 3562
rect 4150 3548 4169 3551
rect 4194 3548 4209 3551
rect 4366 3551 4369 3561
rect 4378 3558 4382 3562
rect 4350 3548 4369 3551
rect 4518 3548 4526 3551
rect 4566 3551 4569 3561
rect 4666 3558 4673 3561
rect 4754 3558 4758 3562
rect 4550 3548 4569 3551
rect 4582 3548 4590 3551
rect 4618 3548 4625 3551
rect 4690 3548 4697 3551
rect 4726 3548 4734 3551
rect 4910 3551 4913 3561
rect 4922 3558 4926 3562
rect 4894 3548 4913 3551
rect 3782 3538 3793 3541
rect 3950 3538 3961 3541
rect 4037 3538 4038 3542
rect 4190 3538 4198 3541
rect 4230 3538 4238 3541
rect 4390 3538 4401 3541
rect 4590 3538 4598 3541
rect 4606 3538 4617 3541
rect 4682 3538 4689 3541
rect 4766 3538 4777 3541
rect 4938 3538 4945 3541
rect 2518 3533 2522 3538
rect 822 3528 841 3531
rect 2646 3528 2649 3538
rect 3550 3531 3554 3533
rect 3798 3531 3802 3533
rect 3542 3528 3554 3531
rect 3790 3528 3802 3531
rect 4246 3531 4250 3533
rect 4414 3531 4418 3533
rect 4238 3528 4250 3531
rect 4406 3528 4418 3531
rect 4686 3528 4689 3538
rect 4790 3531 4794 3533
rect 4782 3528 4794 3531
rect 4958 3531 4962 3533
rect 4950 3528 4962 3531
rect 5102 3528 5121 3531
rect 1293 3518 1294 3522
rect 1413 3518 1414 3522
rect 3770 3518 3771 3522
rect 4638 3518 4654 3521
rect 5061 3518 5062 3522
rect 5157 3518 5158 3522
rect 1048 3503 1050 3507
rect 1054 3503 1057 3507
rect 1061 3503 1064 3507
rect 2072 3503 2074 3507
rect 2078 3503 2081 3507
rect 2085 3503 2088 3507
rect 3096 3503 3098 3507
rect 3102 3503 3105 3507
rect 3109 3503 3112 3507
rect 4112 3503 4114 3507
rect 4118 3503 4121 3507
rect 4125 3503 4128 3507
rect 1397 3488 1398 3492
rect 2557 3488 2558 3492
rect 4466 3488 4467 3492
rect 4662 3488 4678 3491
rect 446 3468 457 3471
rect 614 3468 622 3471
rect 1050 3468 1062 3471
rect 1278 3471 1281 3481
rect 1370 3478 1377 3481
rect 1278 3468 1297 3471
rect 1306 3468 1313 3471
rect 1446 3471 1449 3481
rect 1430 3468 1449 3471
rect 1518 3468 1526 3471
rect 1686 3468 1697 3471
rect 2002 3468 2009 3471
rect 2062 3468 2078 3471
rect 2110 3468 2121 3471
rect 2518 3468 2526 3471
rect 2902 3471 2905 3481
rect 3422 3478 3430 3481
rect 4766 3478 4785 3481
rect 4918 3478 4937 3481
rect 4942 3478 4954 3481
rect 4950 3477 4954 3478
rect 2902 3468 2921 3471
rect 3406 3468 3417 3471
rect 3646 3468 3662 3471
rect 106 3458 113 3461
rect 150 3458 158 3461
rect 190 3458 209 3461
rect 390 3458 409 3461
rect 438 3458 446 3461
rect 474 3458 481 3461
rect 510 3458 526 3461
rect 782 3458 798 3461
rect 846 3461 849 3468
rect 846 3458 857 3461
rect 982 3458 990 3461
rect 1086 3458 1105 3461
rect 1450 3458 1457 3461
rect 1494 3458 1502 3461
rect 1646 3458 1673 3461
rect 1794 3458 1801 3461
rect 1870 3458 1878 3461
rect 1918 3458 1926 3461
rect 2054 3458 2062 3461
rect 2302 3458 2321 3461
rect 2462 3458 2481 3461
rect 2486 3458 2494 3461
rect 3806 3462 3809 3471
rect 4126 3468 4134 3471
rect 4374 3468 4385 3471
rect 2814 3458 2822 3461
rect 3062 3458 3081 3461
rect 3166 3458 3185 3461
rect 3210 3458 3225 3461
rect 3398 3458 3406 3461
rect 3458 3458 3465 3461
rect 3590 3458 3625 3461
rect 4106 3458 4113 3461
rect 4146 3458 4161 3461
rect 4166 3458 4185 3461
rect 4258 3458 4273 3461
rect 4342 3458 4350 3461
rect 4382 3461 4385 3468
rect 4382 3458 4398 3461
rect 4510 3458 4518 3461
rect 4766 3458 4769 3468
rect 134 3448 137 3458
rect 190 3448 193 3458
rect 390 3448 393 3458
rect 434 3448 438 3452
rect 598 3451 601 3458
rect 590 3448 601 3451
rect 950 3448 969 3451
rect 1086 3448 1089 3458
rect 2038 3448 2041 3458
rect 2098 3448 2102 3452
rect 2302 3448 2305 3458
rect 2462 3448 2465 3458
rect 2646 3448 2649 3458
rect 3078 3448 3081 3458
rect 3182 3448 3185 3458
rect 3194 3448 3198 3452
rect 3622 3448 3625 3458
rect 3922 3448 3926 3452
rect 4082 3448 4086 3452
rect 4182 3448 4185 3458
rect 149 3438 150 3442
rect 262 3441 265 3448
rect 3174 3442 3178 3444
rect 254 3438 265 3441
rect 1227 3438 1230 3442
rect 2053 3438 2054 3442
rect 2251 3438 2254 3442
rect 2634 3438 2635 3442
rect 2669 3438 2670 3442
rect 4197 3438 4198 3442
rect 658 3428 659 3432
rect 3466 3428 3467 3432
rect 493 3418 494 3422
rect 557 3418 558 3422
rect 725 3418 726 3422
rect 981 3418 982 3422
rect 1021 3418 1022 3422
rect 1322 3418 1323 3422
rect 1597 3418 1598 3422
rect 1725 3418 1726 3422
rect 2157 3418 2158 3422
rect 3282 3418 3283 3422
rect 3333 3418 3334 3422
rect 3397 3418 3398 3422
rect 3834 3418 3835 3422
rect 4330 3418 4331 3422
rect 4402 3418 4403 3422
rect 4437 3418 4438 3422
rect 5170 3418 5171 3422
rect 536 3403 538 3407
rect 542 3403 545 3407
rect 549 3403 552 3407
rect 1560 3403 1562 3407
rect 1566 3403 1569 3407
rect 1573 3403 1576 3407
rect 2584 3403 2586 3407
rect 2590 3403 2593 3407
rect 2597 3403 2600 3407
rect 3608 3403 3610 3407
rect 3614 3403 3617 3407
rect 3621 3403 3624 3407
rect 4632 3403 4634 3407
rect 4638 3403 4641 3407
rect 4645 3403 4648 3407
rect 1978 3388 1979 3392
rect 4989 3388 4990 3392
rect 1546 3378 1547 3382
rect 554 3368 562 3371
rect 659 3368 662 3372
rect 1558 3368 1574 3371
rect 1842 3368 1845 3372
rect 2042 3368 2043 3372
rect 2202 3368 2203 3372
rect 2622 3368 2633 3371
rect 3090 3368 3091 3372
rect 3309 3368 3310 3372
rect 2622 3366 2626 3368
rect 2942 3366 2946 3368
rect 3518 3366 3522 3368
rect 4006 3366 4010 3368
rect 4062 3366 4066 3368
rect 4934 3366 4938 3368
rect 242 3358 246 3362
rect 166 3348 174 3351
rect 254 3351 257 3361
rect 522 3358 526 3362
rect 254 3348 273 3351
rect 534 3351 537 3361
rect 534 3348 569 3351
rect 718 3351 721 3361
rect 1114 3358 1118 3362
rect 1126 3352 1129 3361
rect 1146 3358 1150 3362
rect 1222 3358 1241 3361
rect 1434 3358 1441 3361
rect 702 3348 721 3351
rect 1138 3348 1145 3351
rect 1198 3348 1214 3351
rect 1234 3348 1249 3351
rect 1362 3348 1377 3351
rect 1538 3348 1545 3351
rect 1262 3338 1289 3341
rect 1474 3338 1481 3341
rect 1526 3338 1529 3348
rect 1790 3351 1793 3361
rect 1774 3348 1793 3351
rect 1806 3348 1814 3351
rect 1922 3348 1929 3351
rect 1990 3351 1993 3361
rect 1990 3348 2009 3351
rect 2014 3348 2022 3351
rect 2030 3338 2033 3348
rect 2214 3351 2217 3361
rect 2194 3348 2201 3351
rect 2214 3348 2233 3351
rect 2310 3351 2313 3361
rect 2322 3358 2326 3362
rect 2430 3358 2441 3361
rect 2538 3358 2542 3362
rect 2430 3356 2434 3358
rect 2550 3352 2553 3361
rect 2582 3358 2617 3361
rect 2834 3358 2838 3362
rect 2294 3348 2313 3351
rect 2530 3348 2537 3351
rect 2662 3348 2670 3351
rect 2846 3351 2849 3361
rect 2886 3352 2889 3361
rect 2894 3358 2913 3361
rect 2846 3348 2865 3351
rect 3102 3351 3105 3361
rect 3102 3348 3137 3351
rect 3198 3348 3206 3351
rect 3294 3351 3297 3361
rect 3586 3358 3590 3362
rect 3278 3348 3297 3351
rect 3310 3348 3318 3351
rect 3378 3348 3385 3351
rect 3814 3351 3817 3361
rect 3774 3348 3793 3351
rect 3798 3348 3817 3351
rect 4182 3351 4185 3361
rect 4426 3358 4430 3362
rect 4554 3358 4558 3362
rect 4954 3358 4958 3362
rect 4166 3348 4185 3351
rect 4610 3348 4617 3351
rect 4902 3348 4918 3351
rect 5114 3348 5129 3351
rect 2478 3338 2486 3341
rect 2718 3338 2730 3341
rect 2934 3338 2942 3341
rect 2966 3338 2974 3341
rect 3774 3341 3777 3348
rect 3766 3338 3777 3341
rect 4366 3338 4377 3341
rect 5102 3338 5110 3341
rect 86 3328 105 3331
rect 2070 3328 2089 3331
rect 2982 3331 2986 3333
rect 2974 3328 2986 3331
rect 3166 3331 3170 3333
rect 4062 3332 4065 3338
rect 4366 3332 4369 3338
rect 3158 3328 3170 3331
rect 4062 3328 4070 3332
rect 4122 3328 4137 3331
rect 853 3318 854 3322
rect 1421 3318 1422 3322
rect 2086 3321 2089 3328
rect 2086 3318 2097 3321
rect 2949 3318 2950 3322
rect 3525 3318 3526 3322
rect 4770 3318 4771 3322
rect 1048 3303 1050 3307
rect 1054 3303 1057 3307
rect 1061 3303 1064 3307
rect 2072 3303 2074 3307
rect 2078 3303 2081 3307
rect 2085 3303 2088 3307
rect 3096 3303 3098 3307
rect 3102 3303 3105 3307
rect 3109 3303 3112 3307
rect 4112 3303 4114 3307
rect 4118 3303 4121 3307
rect 4125 3303 4128 3307
rect 1309 3288 1310 3292
rect 3610 3288 3611 3292
rect 3626 3288 3641 3291
rect 686 3278 705 3281
rect 1902 3278 1913 3281
rect 3126 3278 3145 3281
rect 3218 3278 3234 3281
rect 3910 3278 3921 3281
rect 4222 3278 4230 3281
rect 4462 3278 4474 3281
rect 4926 3278 4945 3281
rect 4950 3278 4962 3281
rect 1902 3277 1906 3278
rect 3230 3274 3234 3278
rect 3910 3277 3914 3278
rect 4470 3277 4474 3278
rect 4958 3277 4962 3278
rect 5142 3278 5153 3281
rect 5142 3277 5146 3278
rect 830 3272 834 3274
rect 278 3268 286 3271
rect 294 3268 302 3271
rect 902 3268 910 3271
rect 1154 3268 1161 3271
rect 1526 3268 1542 3271
rect 1718 3268 1729 3271
rect 2366 3268 2377 3271
rect 2622 3268 2630 3271
rect 2662 3268 2673 3271
rect 2790 3268 2798 3271
rect 2902 3268 2913 3271
rect 178 3258 185 3261
rect 238 3258 246 3261
rect 270 3258 278 3261
rect 358 3258 377 3261
rect 422 3258 430 3261
rect 622 3258 641 3261
rect 850 3258 857 3261
rect 906 3258 913 3261
rect 1262 3258 1270 3261
rect 1494 3258 1513 3261
rect 1650 3258 1657 3261
rect 1766 3258 1785 3261
rect 1798 3258 1806 3261
rect 2902 3262 2905 3268
rect 2982 3262 2985 3271
rect 3022 3268 3033 3271
rect 3106 3268 3113 3271
rect 3402 3268 3417 3271
rect 3506 3268 3513 3271
rect 3702 3268 3713 3271
rect 3742 3268 3753 3271
rect 4422 3268 4430 3271
rect 5046 3268 5058 3271
rect 5158 3268 5169 3271
rect 3030 3262 3033 3268
rect 2078 3258 2113 3261
rect 2230 3258 2238 3261
rect 2318 3258 2337 3261
rect 2390 3258 2417 3261
rect 2506 3258 2513 3261
rect 2574 3258 2609 3261
rect 2638 3258 2646 3261
rect 2686 3258 2713 3261
rect 2770 3258 2777 3261
rect 2822 3258 2841 3261
rect 3078 3258 3094 3261
rect 3126 3258 3129 3268
rect 3750 3262 3753 3268
rect 3310 3258 3318 3261
rect 3426 3258 3433 3261
rect 3682 3258 3689 3261
rect 4122 3258 4137 3261
rect 4166 3258 4185 3261
rect 4198 3258 4214 3261
rect 4270 3258 4286 3261
rect 4422 3258 4441 3261
rect 4522 3258 4529 3261
rect 4598 3258 4617 3261
rect 4826 3258 4833 3261
rect 4898 3258 4905 3261
rect 4926 3258 4929 3268
rect 4990 3258 4998 3261
rect 5170 3258 5177 3261
rect 5182 3258 5190 3261
rect 358 3248 361 3258
rect 622 3248 625 3258
rect 1494 3248 1497 3258
rect 1782 3248 1785 3258
rect 2078 3248 2081 3258
rect 2318 3248 2321 3258
rect 2574 3248 2577 3258
rect 2594 3248 2601 3251
rect 2822 3248 2825 3258
rect 2962 3248 2966 3252
rect 3270 3251 3273 3258
rect 3894 3252 3898 3257
rect 3262 3248 3273 3251
rect 3802 3248 3806 3252
rect 4114 3248 4129 3251
rect 4182 3248 4185 3258
rect 4194 3248 4198 3252
rect 4422 3248 4425 3258
rect 4614 3248 4617 3258
rect 4626 3248 4630 3252
rect 269 3238 270 3242
rect 838 3238 850 3241
rect 1210 3238 1217 3241
rect 1443 3238 1446 3242
rect 2094 3241 2097 3248
rect 2094 3238 2106 3241
rect 3254 3241 3258 3244
rect 2754 3238 2761 3241
rect 3246 3238 3258 3241
rect 3614 3241 3618 3244
rect 3638 3242 3642 3244
rect 3614 3238 3630 3241
rect 4174 3242 4178 3244
rect 3434 3228 3435 3232
rect 3770 3228 3771 3232
rect 346 3218 347 3222
rect 893 3218 894 3222
rect 1189 3218 1190 3222
rect 1245 3218 1246 3222
rect 1738 3218 1739 3222
rect 2429 3218 2430 3222
rect 2877 3218 2878 3222
rect 3477 3218 3478 3222
rect 3570 3218 3571 3222
rect 3994 3218 3995 3222
rect 536 3203 538 3207
rect 542 3203 545 3207
rect 549 3203 552 3207
rect 1560 3203 1562 3207
rect 1566 3203 1569 3207
rect 1573 3203 1576 3207
rect 2584 3203 2586 3207
rect 2590 3203 2593 3207
rect 2597 3203 2600 3207
rect 3608 3203 3610 3207
rect 3614 3203 3617 3207
rect 3621 3203 3624 3207
rect 4632 3203 4634 3207
rect 4638 3203 4641 3207
rect 4645 3203 4648 3207
rect 434 3188 435 3192
rect 2749 3188 2750 3192
rect 2778 3188 2779 3192
rect 2949 3188 2950 3192
rect 1114 3178 1115 3182
rect 1146 3178 1147 3182
rect 1213 3178 1214 3182
rect 1277 3178 1278 3182
rect 3237 3178 3238 3182
rect 346 3168 347 3172
rect 2062 3168 2078 3171
rect 2610 3168 2618 3171
rect 2810 3168 2811 3172
rect 74 3158 78 3162
rect 54 3148 62 3151
rect 78 3148 86 3151
rect 270 3148 278 3151
rect 446 3151 449 3161
rect 738 3158 745 3161
rect 1166 3152 1169 3161
rect 426 3148 433 3151
rect 446 3148 465 3151
rect 534 3148 550 3151
rect 622 3148 630 3151
rect 1214 3148 1238 3151
rect 1262 3151 1265 3161
rect 1246 3148 1265 3151
rect 46 3138 54 3141
rect 86 3138 94 3141
rect 118 3138 121 3148
rect 1494 3148 1505 3151
rect 1550 3151 1553 3161
rect 1590 3161 1593 3168
rect 2982 3166 2986 3168
rect 3470 3168 3481 3171
rect 3746 3168 3753 3171
rect 4010 3168 4013 3172
rect 4834 3168 4837 3172
rect 4922 3168 4923 3172
rect 3470 3166 3474 3168
rect 3758 3166 3762 3168
rect 4486 3166 4490 3168
rect 4958 3166 4962 3168
rect 1590 3158 1601 3161
rect 1698 3158 1705 3161
rect 1550 3148 1585 3151
rect 1706 3148 1713 3151
rect 1878 3151 1881 3161
rect 1502 3142 1505 3148
rect 1878 3148 1886 3151
rect 1934 3148 1942 3151
rect 2102 3151 2105 3161
rect 2326 3158 2345 3161
rect 2354 3158 2358 3162
rect 2102 3148 2110 3151
rect 2134 3142 2137 3151
rect 2358 3148 2366 3151
rect 2490 3148 2497 3151
rect 2590 3151 2593 3161
rect 2590 3148 2625 3151
rect 3054 3151 3057 3161
rect 3026 3148 3033 3151
rect 3038 3148 3057 3151
rect 3222 3151 3225 3161
rect 3206 3148 3225 3151
rect 3350 3151 3353 3158
rect 3350 3148 3361 3151
rect 3598 3148 3606 3151
rect 3798 3151 3801 3161
rect 3762 3148 3777 3151
rect 3782 3148 3801 3151
rect 3958 3151 3961 3161
rect 3942 3148 3961 3151
rect 4494 3151 4497 3161
rect 4750 3158 4769 3161
rect 4978 3158 4982 3162
rect 4478 3148 4497 3151
rect 4690 3148 4697 3151
rect 5126 3148 5134 3151
rect 230 3138 242 3141
rect 494 3138 513 3141
rect 710 3138 718 3141
rect 854 3138 862 3141
rect 1222 3138 1230 3141
rect 1914 3138 1921 3141
rect 2174 3138 2193 3141
rect 2366 3138 2377 3141
rect 2590 3138 2606 3141
rect 3406 3138 3425 3141
rect 4078 3138 4106 3141
rect 4222 3138 4241 3141
rect 4790 3138 4801 3141
rect 14 3128 33 3131
rect 142 3131 146 3133
rect 134 3128 146 3131
rect 510 3128 513 3138
rect 1894 3128 1913 3131
rect 2118 3128 2137 3131
rect 2190 3128 2193 3138
rect 2390 3131 2394 3133
rect 2382 3128 2394 3131
rect 2918 3131 2922 3133
rect 2918 3128 2929 3131
rect 3342 3131 3346 3133
rect 3342 3128 3353 3131
rect 3422 3128 3425 3138
rect 3646 3131 3650 3133
rect 3598 3128 3633 3131
rect 3638 3128 3650 3131
rect 4222 3128 4225 3138
rect 4714 3128 4715 3132
rect 4814 3131 4818 3133
rect 4806 3128 4818 3131
rect 405 3118 406 3122
rect 725 3118 726 3122
rect 789 3118 790 3122
rect 826 3118 827 3122
rect 909 3118 910 3122
rect 1509 3118 1510 3122
rect 1685 3118 1686 3122
rect 2098 3118 2099 3122
rect 1048 3103 1050 3107
rect 1054 3103 1057 3107
rect 1061 3103 1064 3107
rect 2072 3103 2074 3107
rect 2078 3103 2081 3107
rect 2085 3103 2088 3107
rect 3096 3103 3098 3107
rect 3102 3103 3105 3107
rect 3109 3103 3112 3107
rect 4112 3103 4114 3107
rect 4118 3103 4121 3107
rect 4125 3103 4128 3107
rect 109 3088 110 3092
rect 693 3088 694 3092
rect 1242 3088 1243 3092
rect 3058 3088 3059 3092
rect 3338 3088 3339 3092
rect 270 3072 273 3081
rect 278 3078 297 3081
rect 734 3078 746 3081
rect 1394 3078 1401 3081
rect 1654 3078 1662 3081
rect 2158 3078 2170 3081
rect 742 3077 746 3078
rect 2166 3077 2170 3078
rect 50 3058 65 3061
rect 130 3058 137 3061
rect 294 3058 297 3068
rect 326 3062 329 3071
rect 1186 3068 1193 3071
rect 1430 3068 1438 3071
rect 318 3058 326 3061
rect 350 3058 369 3061
rect 454 3058 462 3061
rect 1694 3062 1697 3071
rect 1850 3068 1857 3071
rect 2082 3068 2097 3071
rect 2118 3068 2126 3071
rect 2438 3071 2441 3081
rect 2446 3078 2465 3081
rect 2566 3072 2569 3081
rect 2806 3072 2809 3081
rect 2814 3078 2833 3081
rect 3270 3078 3281 3081
rect 3454 3078 3465 3081
rect 3630 3078 3642 3081
rect 3838 3078 3857 3081
rect 4398 3078 4417 3081
rect 3270 3077 3274 3078
rect 3462 3072 3465 3078
rect 3638 3077 3642 3078
rect 2434 3068 2441 3071
rect 2478 3068 2486 3071
rect 2834 3068 2841 3071
rect 3286 3068 3297 3071
rect 914 3058 921 3061
rect 934 3058 942 3061
rect 1034 3058 1049 3061
rect 1362 3058 1369 3061
rect 1410 3058 1417 3061
rect 1602 3058 1617 3061
rect 2110 3058 2118 3061
rect 2266 3058 2273 3061
rect 2658 3058 2673 3061
rect 3074 3058 3081 3061
rect 3470 3062 3473 3071
rect 3582 3068 3593 3071
rect 3773 3068 3777 3072
rect 4458 3068 4465 3071
rect 4686 3071 4689 3081
rect 4670 3068 4689 3071
rect 5098 3068 5105 3071
rect 5126 3068 5137 3071
rect 3590 3062 3593 3068
rect 3774 3062 3777 3068
rect 3542 3058 3561 3061
rect 3854 3058 3857 3068
rect 5126 3062 5129 3068
rect 3966 3058 3982 3061
rect 4158 3058 4166 3061
rect 4310 3058 4318 3061
rect 4542 3058 4561 3061
rect 4598 3058 4606 3061
rect 4658 3058 4665 3061
rect 4818 3058 4825 3061
rect 4830 3058 4849 3061
rect 4930 3058 4937 3061
rect 5030 3058 5049 3061
rect 5086 3058 5105 3061
rect 5146 3058 5161 3061
rect 350 3048 353 3058
rect 638 3048 657 3051
rect 918 3048 921 3058
rect 1054 3048 1081 3051
rect 1414 3048 1417 3058
rect 2274 3048 2278 3052
rect 2310 3051 2313 3058
rect 2302 3048 2313 3051
rect 2574 3051 2577 3058
rect 2574 3048 2585 3051
rect 2906 3048 2910 3052
rect 3558 3048 3561 3058
rect 4054 3048 4073 3051
rect 4494 3048 4505 3051
rect 4542 3048 4545 3058
rect 4846 3048 4849 3058
rect 5046 3048 5049 3058
rect 5102 3048 5105 3058
rect 1078 3042 1082 3044
rect 1474 3038 1481 3041
rect 1942 3041 1945 3048
rect 1934 3038 1945 3041
rect 2502 3038 2510 3041
rect 4078 3041 4082 3044
rect 4494 3042 4497 3048
rect 4078 3038 4086 3041
rect 4346 3038 4347 3042
rect 4738 3038 4741 3042
rect 4861 3038 4862 3042
rect 4898 3038 4901 3042
rect 4597 3028 4598 3032
rect 149 3018 150 3022
rect 338 3018 339 3022
rect 669 3018 670 3022
rect 933 3018 934 3022
rect 1157 3018 1158 3022
rect 1370 3018 1371 3022
rect 1714 3018 1715 3022
rect 1821 3018 1822 3022
rect 4005 3018 4006 3022
rect 4530 3018 4531 3022
rect 536 3003 538 3007
rect 542 3003 545 3007
rect 549 3003 552 3007
rect 1560 3003 1562 3007
rect 1566 3003 1569 3007
rect 1573 3003 1576 3007
rect 2584 3003 2586 3007
rect 2590 3003 2593 3007
rect 2597 3003 2600 3007
rect 3608 3003 3610 3007
rect 3614 3003 3617 3007
rect 3621 3003 3624 3007
rect 4632 3003 4634 3007
rect 4638 3003 4641 3007
rect 4645 3003 4648 3007
rect 901 2988 902 2992
rect 3722 2988 3723 2992
rect 3986 2988 3987 2992
rect 1802 2978 1803 2982
rect 565 2968 566 2972
rect 1470 2968 1478 2971
rect 4126 2968 4134 2971
rect 4198 2968 4206 2971
rect 4482 2968 4485 2972
rect 4994 2968 4997 2972
rect 1654 2966 1658 2968
rect 3686 2966 3690 2968
rect 4126 2966 4130 2968
rect 4198 2966 4202 2968
rect 4222 2966 4226 2968
rect 370 2958 374 2962
rect 126 2942 129 2951
rect 382 2951 385 2961
rect 514 2958 518 2962
rect 538 2958 553 2961
rect 738 2958 742 2962
rect 770 2958 774 2962
rect 362 2948 369 2951
rect 382 2948 401 2951
rect 474 2948 481 2951
rect 710 2948 726 2951
rect 838 2948 849 2951
rect 974 2948 982 2951
rect 1074 2948 1081 2951
rect 1166 2951 1169 2961
rect 1362 2958 1366 2962
rect 1630 2958 1649 2961
rect 1654 2958 1665 2961
rect 1674 2958 1678 2962
rect 1834 2958 1838 2962
rect 1846 2952 1849 2961
rect 1942 2958 1953 2961
rect 2302 2958 2321 2961
rect 2474 2958 2478 2962
rect 2562 2958 2569 2961
rect 1942 2956 1946 2958
rect 1162 2948 1169 2951
rect 838 2942 841 2948
rect 218 2938 225 2941
rect 610 2938 625 2941
rect 722 2938 729 2941
rect 978 2938 993 2941
rect 1126 2938 1142 2941
rect 1342 2938 1345 2948
rect 1526 2948 1534 2951
rect 1694 2938 1697 2948
rect 2254 2948 2262 2951
rect 2466 2948 2473 2951
rect 2622 2948 2649 2951
rect 2790 2951 2793 2961
rect 2942 2958 2961 2961
rect 3130 2958 3134 2962
rect 2774 2948 2793 2951
rect 2806 2948 2814 2951
rect 2962 2948 2969 2951
rect 2446 2941 2449 2948
rect 2446 2938 2465 2941
rect 2830 2941 2833 2948
rect 3142 2951 3145 2961
rect 3190 2951 3193 2961
rect 3142 2948 3161 2951
rect 3190 2948 3198 2951
rect 3494 2942 3497 2951
rect 3678 2948 3689 2951
rect 3798 2951 3801 2961
rect 3810 2958 3814 2962
rect 3782 2948 3801 2951
rect 3686 2942 3689 2948
rect 4258 2948 4265 2951
rect 4582 2951 4585 2961
rect 4566 2948 4585 2951
rect 4926 2951 4929 2961
rect 4918 2948 4929 2951
rect 5090 2948 5097 2951
rect 2814 2938 2833 2941
rect 2982 2938 2990 2941
rect 3114 2938 3121 2941
rect 3182 2938 3190 2941
rect 3822 2938 3833 2941
rect 4694 2938 4702 2941
rect 110 2928 129 2931
rect 166 2928 185 2931
rect 934 2928 953 2931
rect 1134 2928 1153 2931
rect 2030 2928 2049 2931
rect 2054 2928 2070 2931
rect 2242 2928 2243 2932
rect 2438 2931 2442 2933
rect 2542 2932 2545 2938
rect 2438 2928 2449 2931
rect 2542 2928 2550 2932
rect 2838 2931 2842 2933
rect 3006 2931 3010 2933
rect 2830 2928 2842 2931
rect 2998 2928 3010 2931
rect 3206 2928 3225 2931
rect 3654 2928 3673 2931
rect 4302 2928 4321 2931
rect 4462 2931 4466 2933
rect 4454 2928 4466 2931
rect 4902 2931 4905 2938
rect 4918 2932 4921 2948
rect 4902 2928 4913 2931
rect 445 2918 446 2922
rect 1173 2918 1174 2922
rect 1957 2918 1958 2922
rect 2194 2918 2195 2922
rect 2573 2918 2574 2922
rect 3654 2921 3657 2928
rect 3646 2918 3657 2921
rect 4122 2918 4123 2922
rect 4218 2918 4219 2922
rect 4933 2918 4934 2922
rect 4962 2918 4963 2922
rect 5077 2918 5078 2922
rect 1048 2903 1050 2907
rect 1054 2903 1057 2907
rect 1061 2903 1064 2907
rect 2072 2903 2074 2907
rect 2078 2903 2081 2907
rect 2085 2903 2088 2907
rect 3096 2903 3098 2907
rect 3102 2903 3105 2907
rect 3109 2903 3112 2907
rect 4112 2903 4114 2907
rect 4118 2903 4121 2907
rect 4125 2903 4128 2907
rect 2082 2888 2089 2891
rect 2277 2888 2278 2892
rect 3354 2888 3355 2892
rect 406 2878 414 2881
rect 510 2878 521 2881
rect 1106 2878 1107 2882
rect 2678 2878 2690 2881
rect 3650 2878 3651 2882
rect 4934 2878 4946 2881
rect 510 2877 514 2878
rect 2686 2877 2690 2878
rect 4942 2877 4946 2878
rect 5118 2872 5121 2878
rect 678 2868 689 2871
rect 946 2868 961 2871
rect 974 2868 990 2871
rect 1566 2868 1574 2871
rect 2086 2868 2105 2871
rect 2126 2868 2134 2871
rect 366 2858 385 2861
rect 526 2858 534 2861
rect 710 2858 729 2861
rect 1074 2858 1089 2861
rect 1318 2858 1337 2861
rect 1478 2858 1497 2861
rect 1682 2858 1697 2861
rect 1702 2858 1721 2861
rect 1802 2858 1809 2861
rect 1922 2858 1937 2861
rect 1962 2858 1969 2861
rect 2126 2858 2145 2861
rect 2258 2858 2265 2861
rect 2294 2858 2302 2861
rect 2414 2862 2417 2871
rect 2662 2868 2678 2871
rect 2438 2858 2457 2861
rect 2490 2858 2505 2861
rect 2782 2862 2785 2871
rect 2986 2868 2993 2871
rect 3030 2868 3049 2871
rect 3254 2868 3262 2871
rect 3314 2868 3329 2871
rect 4026 2868 4041 2871
rect 4278 2868 4294 2871
rect 4678 2868 4697 2871
rect 5038 2868 5057 2871
rect 5118 2868 5122 2872
rect 5174 2868 5182 2871
rect 2806 2858 2825 2861
rect 2862 2858 2881 2861
rect 3050 2858 3057 2861
rect 3234 2858 3241 2861
rect 3302 2858 3310 2861
rect 3662 2858 3689 2861
rect 3734 2858 3742 2861
rect 3830 2858 3838 2861
rect 3930 2858 3937 2861
rect 4114 2858 4137 2861
rect 4614 2858 4649 2861
rect 4718 2858 4737 2861
rect 4986 2858 5001 2861
rect 5138 2858 5145 2861
rect 366 2848 369 2858
rect 710 2848 713 2858
rect 1318 2848 1321 2858
rect 1466 2848 1470 2852
rect 1478 2848 1481 2858
rect 1534 2851 1537 2858
rect 1526 2848 1537 2851
rect 1718 2848 1721 2858
rect 2126 2848 2129 2858
rect 2426 2848 2430 2852
rect 2438 2848 2441 2858
rect 2478 2848 2497 2851
rect 2650 2848 2654 2852
rect 2806 2848 2809 2858
rect 2862 2848 2865 2858
rect 3218 2848 3222 2852
rect 4162 2848 4169 2851
rect 4622 2848 4638 2851
rect 4646 2848 4649 2858
rect 4718 2848 4721 2858
rect 491 2838 494 2842
rect 1267 2838 1270 2842
rect 2706 2838 2709 2842
rect 2794 2838 2795 2842
rect 4213 2838 4214 2842
rect 3386 2828 3387 2832
rect 3938 2828 3939 2832
rect 757 2818 758 2822
rect 1045 2818 1046 2822
rect 1733 2818 1734 2822
rect 1866 2818 1867 2822
rect 2050 2818 2051 2822
rect 2546 2818 2547 2822
rect 2850 2818 2851 2822
rect 2957 2818 2958 2822
rect 3290 2818 3291 2822
rect 4090 2818 4091 2822
rect 4482 2818 4483 2822
rect 4530 2818 4531 2822
rect 4661 2818 4662 2822
rect 536 2803 538 2807
rect 542 2803 545 2807
rect 549 2803 552 2807
rect 1560 2803 1562 2807
rect 1566 2803 1569 2807
rect 1573 2803 1576 2807
rect 2584 2803 2586 2807
rect 2590 2803 2593 2807
rect 2597 2803 2600 2807
rect 3608 2803 3610 2807
rect 3614 2803 3617 2807
rect 3621 2803 3624 2807
rect 4632 2803 4634 2807
rect 4638 2803 4641 2807
rect 4645 2803 4648 2807
rect 3165 2788 3166 2792
rect 3906 2788 3907 2792
rect 4234 2788 4235 2792
rect 4850 2788 4851 2792
rect 4914 2788 4915 2792
rect 4978 2788 4979 2792
rect 219 2768 222 2772
rect 790 2768 802 2771
rect 2022 2768 2033 2771
rect 2910 2768 2921 2771
rect 3626 2768 3627 2772
rect 4270 2768 4281 2771
rect 798 2766 802 2768
rect 2030 2762 2033 2768
rect 3662 2766 3666 2768
rect 4270 2766 4274 2768
rect 490 2758 497 2761
rect 526 2758 542 2761
rect 574 2758 593 2761
rect 598 2758 610 2761
rect 606 2756 610 2758
rect 506 2748 513 2751
rect 734 2748 742 2751
rect 1246 2751 1249 2761
rect 1258 2758 1262 2762
rect 1230 2748 1249 2751
rect 1470 2751 1473 2761
rect 1482 2758 1486 2762
rect 1454 2748 1473 2751
rect 1858 2748 1865 2751
rect 494 2738 505 2741
rect 826 2738 833 2741
rect 1046 2738 1054 2741
rect 1190 2738 1209 2741
rect 1270 2738 1281 2741
rect 1418 2738 1425 2741
rect 1494 2738 1505 2741
rect 1790 2741 1793 2748
rect 2014 2751 2017 2761
rect 2010 2748 2017 2751
rect 2118 2748 2145 2751
rect 2222 2751 2225 2761
rect 2778 2758 2782 2762
rect 2222 2748 2241 2751
rect 2450 2748 2457 2751
rect 2702 2748 2710 2751
rect 2790 2751 2793 2761
rect 2898 2758 2902 2762
rect 2790 2748 2809 2751
rect 2850 2748 2865 2751
rect 2882 2748 2897 2751
rect 3150 2751 3153 2761
rect 3638 2758 3657 2761
rect 3918 2758 3937 2761
rect 2970 2748 2977 2751
rect 3134 2748 3153 2751
rect 3226 2748 3233 2751
rect 3462 2748 3473 2751
rect 3666 2748 3673 2751
rect 3698 2748 3705 2751
rect 1774 2738 1793 2741
rect 1846 2738 1862 2741
rect 1990 2738 2001 2741
rect 2182 2738 2201 2741
rect 2222 2738 2230 2741
rect 2394 2738 2402 2741
rect 2550 2738 2561 2741
rect 2654 2738 2662 2741
rect 3102 2738 3118 2741
rect 3230 2741 3233 2748
rect 3470 2742 3473 2748
rect 3890 2748 3897 2751
rect 3982 2751 3985 2761
rect 4246 2758 4265 2761
rect 3946 2748 3961 2751
rect 3966 2748 3985 2751
rect 4066 2748 4073 2751
rect 4158 2748 4169 2751
rect 3174 2738 3193 2741
rect 3230 2738 3241 2741
rect 3602 2738 3617 2741
rect 3718 2738 3726 2741
rect 3894 2738 3897 2748
rect 4166 2741 4169 2748
rect 4402 2748 4409 2751
rect 4550 2748 4569 2751
rect 4842 2748 4849 2751
rect 4166 2738 4185 2741
rect 4366 2738 4374 2741
rect 4606 2738 4614 2741
rect 4694 2738 4713 2741
rect 478 2731 482 2733
rect 478 2728 489 2731
rect 862 2728 870 2731
rect 1190 2728 1193 2738
rect 1294 2731 1298 2733
rect 1990 2732 1993 2738
rect 1286 2728 1298 2731
rect 1510 2728 1529 2731
rect 1654 2728 1673 2731
rect 2486 2731 2490 2733
rect 2934 2732 2938 2736
rect 4294 2732 4298 2736
rect 2486 2728 2497 2731
rect 4710 2728 4713 2738
rect 373 2718 374 2722
rect 1397 2718 1398 2722
rect 1526 2721 1529 2728
rect 1526 2718 1537 2721
rect 1693 2718 1694 2722
rect 1797 2718 1798 2722
rect 2370 2718 2371 2722
rect 2582 2718 2590 2721
rect 2837 2718 2838 2722
rect 4146 2718 4147 2722
rect 1048 2703 1050 2707
rect 1054 2703 1057 2707
rect 1061 2703 1064 2707
rect 2072 2703 2074 2707
rect 2078 2703 2081 2707
rect 2085 2703 2088 2707
rect 3096 2703 3098 2707
rect 3102 2703 3105 2707
rect 3109 2703 3112 2707
rect 4112 2703 4114 2707
rect 4118 2703 4121 2707
rect 4125 2703 4128 2707
rect 546 2688 561 2691
rect 701 2688 702 2692
rect 4610 2688 4611 2692
rect 4930 2688 4931 2692
rect 94 2678 102 2681
rect 110 2678 129 2681
rect 197 2678 198 2682
rect 286 2678 305 2681
rect 326 2678 345 2681
rect 462 2678 473 2681
rect 734 2678 746 2681
rect 878 2678 890 2681
rect 1078 2678 1097 2681
rect 1350 2678 1361 2681
rect 1525 2678 1526 2682
rect 1550 2678 1558 2682
rect 1902 2678 1913 2681
rect 1918 2678 1937 2681
rect 2038 2678 2057 2681
rect 2062 2678 2078 2681
rect 2242 2678 2246 2682
rect 3262 2678 3273 2681
rect 3494 2678 3505 2681
rect 3750 2678 3769 2681
rect 94 2677 98 2678
rect 462 2677 466 2678
rect 742 2677 746 2678
rect 886 2677 890 2678
rect 1350 2677 1354 2678
rect 1550 2672 1553 2678
rect 1902 2677 1906 2678
rect 3262 2677 3266 2678
rect 3494 2677 3498 2678
rect 1894 2672 1898 2674
rect 130 2668 137 2671
rect 478 2668 489 2671
rect 510 2668 518 2671
rect 1070 2668 1086 2671
rect 1370 2668 1377 2671
rect 1454 2668 1465 2671
rect 1774 2668 1785 2671
rect 2066 2668 2097 2671
rect 2226 2668 2233 2671
rect 2274 2668 2281 2671
rect 2298 2668 2305 2671
rect 2718 2668 2726 2671
rect 174 2658 182 2661
rect 510 2658 529 2661
rect 1006 2658 1025 2661
rect 1050 2658 1057 2661
rect 1414 2658 1433 2661
rect 1622 2658 1638 2661
rect 1690 2658 1697 2661
rect 1786 2658 1793 2661
rect 1846 2658 1854 2661
rect 2038 2658 2041 2668
rect 2162 2658 2169 2661
rect 2390 2658 2409 2661
rect 2830 2662 2833 2671
rect 3090 2668 3121 2671
rect 3278 2668 3289 2671
rect 3510 2668 3521 2671
rect 3610 2668 3617 2671
rect 3650 2668 3657 2671
rect 3918 2671 3921 2681
rect 4054 2678 4073 2681
rect 4326 2678 4345 2681
rect 4702 2672 4706 2674
rect 3902 2668 3921 2671
rect 2582 2658 2598 2661
rect 2602 2658 2609 2661
rect 2666 2658 2673 2661
rect 2866 2658 2873 2661
rect 2926 2658 2934 2661
rect 3006 2658 3022 2661
rect 3206 2658 3214 2661
rect 3310 2658 3329 2661
rect 3358 2658 3374 2661
rect 3518 2662 3521 2668
rect 4486 2662 4489 2671
rect 4498 2668 4505 2671
rect 4594 2668 4601 2671
rect 5014 2668 5022 2671
rect 5054 2668 5062 2671
rect 5094 2671 5097 2681
rect 5102 2678 5121 2681
rect 5090 2668 5097 2671
rect 3602 2658 3625 2661
rect 3630 2658 3657 2661
rect 4002 2658 4009 2661
rect 4126 2658 4134 2661
rect 4142 2658 4153 2661
rect 4210 2658 4217 2661
rect 4446 2658 4465 2661
rect 4626 2658 4649 2661
rect 4654 2658 4662 2661
rect 4726 2658 4734 2661
rect 4866 2658 4881 2661
rect 4950 2658 4966 2661
rect 510 2648 513 2658
rect 850 2648 854 2652
rect 994 2648 998 2652
rect 1006 2648 1009 2658
rect 1214 2648 1233 2651
rect 1386 2648 1390 2652
rect 2082 2648 2089 2651
rect 2406 2648 2409 2658
rect 3310 2648 3313 2658
rect 4142 2652 4145 2658
rect 3338 2648 3345 2651
rect 3386 2648 3390 2652
rect 4462 2648 4465 2658
rect 4670 2651 4673 2658
rect 4670 2648 4681 2651
rect 5034 2648 5038 2652
rect 5074 2648 5081 2651
rect 2206 2642 2210 2644
rect 762 2638 765 2642
rect 906 2638 909 2642
rect 1179 2638 1182 2642
rect 1474 2638 1481 2641
rect 1659 2638 1662 2642
rect 2246 2642 2250 2644
rect 2534 2642 2538 2644
rect 3698 2638 3705 2641
rect 4686 2641 4690 2644
rect 4686 2638 4697 2641
rect 1445 2618 1446 2622
rect 1794 2618 1795 2622
rect 1986 2618 1987 2622
rect 2874 2618 2875 2622
rect 3357 2618 3358 2622
rect 536 2603 538 2607
rect 542 2603 545 2607
rect 549 2603 552 2607
rect 1560 2603 1562 2607
rect 1566 2603 1569 2607
rect 1573 2603 1576 2607
rect 2584 2603 2586 2607
rect 2590 2603 2593 2607
rect 2597 2603 2600 2607
rect 3608 2603 3610 2607
rect 3614 2603 3617 2607
rect 3621 2603 3624 2607
rect 4632 2603 4634 2607
rect 4638 2603 4641 2607
rect 4645 2603 4648 2607
rect 778 2588 779 2592
rect 1522 2588 1523 2592
rect 1701 2588 1702 2592
rect 3741 2588 3742 2592
rect 4866 2588 4867 2592
rect 1805 2578 1806 2582
rect 510 2568 526 2571
rect 1346 2568 1353 2571
rect 2646 2568 2654 2571
rect 3090 2568 3093 2572
rect 3966 2568 3977 2571
rect 4650 2568 4657 2571
rect 5102 2568 5110 2571
rect 3966 2566 3970 2568
rect 482 2558 486 2562
rect 102 2542 105 2551
rect 486 2548 494 2551
rect 538 2548 553 2551
rect 790 2551 793 2561
rect 1042 2558 1046 2562
rect 1142 2558 1150 2561
rect 1370 2558 1374 2562
rect 790 2548 798 2551
rect 1074 2548 1081 2551
rect 1382 2551 1385 2561
rect 1382 2548 1401 2551
rect 1470 2551 1473 2561
rect 1482 2558 1486 2562
rect 1454 2548 1473 2551
rect 1686 2551 1689 2561
rect 2450 2558 2454 2562
rect 1670 2548 1689 2551
rect 1774 2548 1782 2551
rect 2138 2548 2145 2551
rect 2274 2548 2281 2551
rect 2326 2548 2334 2551
rect 2502 2548 2510 2551
rect 2734 2548 2742 2551
rect 2758 2551 2761 2558
rect 2750 2548 2761 2551
rect 2974 2551 2977 2561
rect 2974 2548 2993 2551
rect 3190 2551 3193 2561
rect 3438 2558 3449 2561
rect 3438 2556 3442 2558
rect 3190 2548 3209 2551
rect 3494 2551 3497 2561
rect 3506 2558 3510 2562
rect 3478 2548 3497 2551
rect 3742 2548 3750 2551
rect 3806 2551 3809 2561
rect 4310 2558 4321 2561
rect 4310 2556 4314 2558
rect 3806 2548 3825 2551
rect 4006 2548 4014 2551
rect 118 2538 134 2541
rect 406 2538 425 2541
rect 1066 2538 1078 2541
rect 1082 2538 1089 2541
rect 1094 2538 1102 2541
rect 1350 2538 1361 2541
rect 1862 2538 1870 2541
rect 2006 2538 2014 2541
rect 2038 2538 2046 2541
rect 2062 2538 2094 2541
rect 2262 2538 2281 2541
rect 2590 2538 2625 2541
rect 2666 2538 2673 2541
rect 2698 2538 2713 2541
rect 3302 2538 3321 2541
rect 3646 2538 3654 2541
rect 3774 2541 3777 2548
rect 4190 2542 4193 2551
rect 4398 2548 4406 2551
rect 3774 2538 3785 2541
rect 3806 2538 3814 2541
rect 3838 2538 3846 2541
rect 4114 2538 4129 2541
rect 4358 2538 4366 2541
rect 4406 2541 4409 2548
rect 4630 2548 4638 2551
rect 4806 2542 4809 2551
rect 5166 2548 5190 2551
rect 4406 2538 4417 2541
rect 4846 2538 4857 2541
rect 5006 2538 5018 2541
rect 406 2528 409 2538
rect 866 2528 873 2531
rect 878 2528 881 2538
rect 934 2531 938 2533
rect 926 2528 938 2531
rect 1102 2528 1121 2531
rect 1218 2528 1219 2532
rect 1334 2531 1338 2533
rect 2278 2532 2281 2538
rect 1334 2528 1345 2531
rect 2590 2528 2593 2538
rect 2602 2528 2617 2531
rect 3046 2528 3065 2531
rect 3318 2528 3321 2538
rect 3622 2528 3641 2531
rect 4190 2528 4209 2531
rect 4214 2528 4217 2538
rect 4590 2528 4609 2531
rect 4806 2528 4825 2531
rect 565 2518 566 2522
rect 629 2518 630 2522
rect 1890 2518 1891 2522
rect 1925 2518 1926 2522
rect 2714 2518 2715 2522
rect 2774 2518 2782 2521
rect 3062 2521 3065 2528
rect 3062 2518 3073 2521
rect 3453 2518 3454 2522
rect 3622 2521 3625 2528
rect 3614 2518 3625 2521
rect 3666 2518 3667 2522
rect 3770 2518 3771 2522
rect 3962 2518 3963 2522
rect 4570 2518 4571 2522
rect 5122 2518 5123 2522
rect 5146 2518 5147 2522
rect 1048 2503 1050 2507
rect 1054 2503 1057 2507
rect 1061 2503 1064 2507
rect 2072 2503 2074 2507
rect 2078 2503 2081 2507
rect 2085 2503 2088 2507
rect 3096 2503 3098 2507
rect 3102 2503 3105 2507
rect 3109 2503 3112 2507
rect 4112 2503 4114 2507
rect 4118 2503 4121 2507
rect 4125 2503 4128 2507
rect 1810 2488 1811 2492
rect 2005 2488 2006 2492
rect 2029 2488 2030 2492
rect 2141 2488 2142 2492
rect 4077 2488 4078 2492
rect 262 2478 274 2481
rect 478 2478 489 2481
rect 270 2477 274 2478
rect 478 2477 482 2478
rect 862 2468 873 2471
rect 926 2471 929 2481
rect 906 2468 913 2471
rect 926 2468 945 2471
rect 1250 2468 1257 2471
rect 46 2458 58 2461
rect 314 2458 329 2461
rect 518 2458 526 2461
rect 614 2458 633 2461
rect 662 2458 670 2461
rect 874 2458 881 2461
rect 1294 2462 1297 2471
rect 1518 2471 1521 2481
rect 1630 2478 1641 2481
rect 1646 2478 1657 2481
rect 2578 2478 2582 2482
rect 2794 2478 2795 2482
rect 3446 2478 3454 2482
rect 4162 2478 4166 2482
rect 4630 2478 4646 2481
rect 4790 2478 4809 2481
rect 1654 2472 1657 2478
rect 3446 2472 3449 2478
rect 4886 2472 4889 2481
rect 5110 2478 5129 2481
rect 1518 2468 1537 2471
rect 1662 2468 1670 2471
rect 1846 2468 1854 2471
rect 2074 2468 2097 2471
rect 2142 2468 2158 2471
rect 2390 2468 2417 2471
rect 2454 2468 2481 2471
rect 2494 2468 2502 2471
rect 2550 2468 2566 2471
rect 2746 2468 2753 2471
rect 2910 2468 2937 2471
rect 2962 2468 2969 2471
rect 2974 2468 3001 2471
rect 3150 2468 3158 2471
rect 3350 2468 3358 2471
rect 3370 2468 3377 2471
rect 3494 2468 3521 2471
rect 3838 2468 3862 2471
rect 3878 2468 3894 2471
rect 3950 2468 3958 2471
rect 4146 2468 4161 2471
rect 4342 2468 4369 2471
rect 4438 2468 4449 2471
rect 4554 2468 4561 2471
rect 4614 2468 4625 2471
rect 1270 2458 1278 2461
rect 1362 2458 1369 2461
rect 1606 2458 1614 2461
rect 1638 2458 1657 2461
rect 1978 2458 1985 2461
rect 2118 2458 2121 2468
rect 2562 2458 2569 2461
rect 2650 2458 2665 2461
rect 2806 2458 2814 2461
rect 2854 2458 2881 2461
rect 2958 2458 2966 2461
rect 3122 2458 3129 2461
rect 3158 2458 3166 2461
rect 3226 2458 3233 2461
rect 3438 2458 3446 2461
rect 3486 2458 3494 2461
rect 3542 2458 3561 2461
rect 3602 2458 3609 2461
rect 4446 2462 4449 2468
rect 3850 2458 3857 2461
rect 3890 2458 3897 2461
rect 3926 2458 3934 2461
rect 4062 2458 4070 2461
rect 4090 2458 4097 2461
rect 4182 2458 4190 2461
rect 4254 2458 4262 2461
rect 4390 2458 4409 2461
rect 4518 2458 4526 2461
rect 54 2457 58 2458
rect 286 2452 290 2457
rect 602 2448 606 2452
rect 614 2448 617 2458
rect 1142 2452 1146 2457
rect 2062 2448 2078 2451
rect 2634 2448 2638 2452
rect 3306 2448 3310 2452
rect 3466 2448 3473 2451
rect 3542 2448 3545 2458
rect 3606 2451 3609 2458
rect 3606 2448 3617 2451
rect 4330 2448 4334 2452
rect 4378 2448 4382 2452
rect 4390 2448 4393 2458
rect 4602 2448 4606 2452
rect 4846 2448 4854 2451
rect 2214 2442 2218 2444
rect 1926 2438 1934 2441
rect 4506 2428 4507 2432
rect 786 2418 787 2422
rect 2842 2418 2843 2422
rect 4762 2418 4763 2422
rect 536 2403 538 2407
rect 542 2403 545 2407
rect 549 2403 552 2407
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1573 2403 1576 2407
rect 2584 2403 2586 2407
rect 2590 2403 2593 2407
rect 2597 2403 2600 2407
rect 3608 2403 3610 2407
rect 3614 2403 3617 2407
rect 3621 2403 3624 2407
rect 4632 2403 4634 2407
rect 4638 2403 4641 2407
rect 4645 2403 4648 2407
rect 1189 2388 1190 2392
rect 1293 2388 1294 2392
rect 2677 2388 2678 2392
rect 2786 2388 2787 2392
rect 4181 2388 4182 2392
rect 4370 2388 4371 2392
rect 4858 2388 4859 2392
rect 4770 2378 4771 2382
rect 378 2368 379 2372
rect 538 2368 546 2371
rect 837 2368 838 2372
rect 1910 2368 1918 2371
rect 170 2358 174 2362
rect 506 2358 510 2362
rect 30 2351 34 2353
rect 22 2348 34 2351
rect 142 2348 150 2351
rect 290 2348 297 2351
rect 518 2351 521 2361
rect 646 2352 649 2361
rect 518 2348 553 2351
rect 578 2348 585 2351
rect 686 2348 694 2351
rect 774 2348 790 2351
rect 918 2341 921 2348
rect 1110 2342 1113 2351
rect 1262 2348 1270 2351
rect 1322 2348 1329 2351
rect 1598 2351 1601 2361
rect 1598 2348 1617 2351
rect 1790 2348 1798 2351
rect 910 2338 921 2341
rect 1138 2338 1153 2341
rect 1242 2338 1249 2341
rect 1390 2341 1393 2348
rect 1902 2348 1913 2351
rect 1934 2348 1945 2351
rect 1962 2348 1969 2351
rect 2062 2348 2070 2351
rect 2210 2348 2217 2351
rect 2246 2348 2254 2351
rect 2350 2351 2353 2361
rect 2954 2358 2958 2362
rect 2350 2348 2369 2351
rect 2426 2348 2441 2351
rect 2586 2348 2593 2351
rect 2730 2348 2737 2351
rect 2966 2351 2969 2361
rect 2966 2348 2985 2351
rect 3134 2348 3142 2351
rect 1942 2342 1945 2348
rect 3302 2342 3305 2351
rect 3406 2351 3409 2361
rect 3402 2348 3409 2351
rect 3822 2348 3830 2351
rect 3854 2351 3857 2361
rect 3866 2358 3870 2362
rect 4810 2358 4814 2362
rect 4886 2358 4894 2361
rect 4918 2358 4930 2361
rect 4926 2356 4930 2358
rect 5070 2358 5081 2361
rect 5134 2361 5137 2368
rect 5150 2366 5154 2368
rect 5134 2358 5145 2361
rect 5070 2352 5073 2358
rect 3838 2348 3857 2351
rect 3938 2348 3945 2351
rect 4078 2348 4086 2351
rect 4110 2348 4134 2351
rect 5154 2348 5161 2351
rect 1382 2338 1393 2341
rect 1562 2338 1577 2341
rect 1714 2338 1729 2341
rect 2014 2338 2022 2341
rect 2090 2338 2097 2341
rect 2154 2338 2161 2341
rect 2218 2338 2225 2341
rect 2238 2338 2246 2341
rect 2250 2338 2265 2341
rect 2350 2338 2358 2341
rect 2606 2338 2614 2341
rect 3190 2338 3198 2341
rect 3582 2338 3617 2341
rect 3774 2338 3801 2341
rect 4050 2338 4057 2341
rect 4458 2338 4465 2341
rect 4910 2338 4918 2341
rect 5162 2338 5169 2341
rect 742 2331 746 2333
rect 742 2328 753 2331
rect 1462 2331 1466 2333
rect 1070 2328 1089 2331
rect 1094 2328 1113 2331
rect 1454 2328 1466 2331
rect 2298 2328 2302 2332
rect 3374 2328 3393 2331
rect 3546 2328 3547 2332
rect 3590 2328 3598 2331
rect 3614 2328 3617 2338
rect 4022 2332 4025 2338
rect 4022 2328 4030 2332
rect 4438 2328 4457 2331
rect 5046 2328 5054 2331
rect 1070 2322 1073 2328
rect 309 2318 310 2322
rect 1062 2318 1070 2321
rect 1741 2318 1742 2322
rect 2197 2318 2198 2322
rect 3802 2318 3803 2322
rect 1048 2303 1050 2307
rect 1054 2303 1057 2307
rect 1061 2303 1064 2307
rect 2072 2303 2074 2307
rect 2078 2303 2081 2307
rect 2085 2303 2088 2307
rect 3096 2303 3098 2307
rect 3102 2303 3105 2307
rect 3109 2303 3112 2307
rect 4112 2303 4114 2307
rect 4118 2303 4121 2307
rect 4125 2303 4128 2307
rect 1566 2288 1574 2291
rect 1645 2288 1646 2292
rect 1470 2278 1478 2281
rect 1970 2278 1982 2281
rect 2906 2278 2913 2281
rect 2978 2278 2985 2281
rect 3190 2278 3202 2281
rect 3578 2278 3585 2281
rect 1470 2277 1474 2278
rect 3198 2277 3202 2278
rect 3590 2272 3593 2281
rect 3854 2278 3873 2281
rect 4518 2278 4530 2281
rect 4526 2277 4530 2278
rect 5054 2272 5058 2274
rect 170 2268 177 2271
rect 410 2268 411 2272
rect 462 2268 473 2271
rect 586 2268 593 2271
rect 1306 2268 1313 2271
rect 1330 2268 1353 2271
rect 1762 2268 1769 2271
rect 1830 2268 1838 2271
rect 1874 2268 1889 2271
rect 1998 2268 2009 2271
rect 2018 2268 2033 2271
rect 2082 2268 2105 2271
rect 2170 2268 2177 2271
rect 2330 2268 2337 2271
rect 2534 2268 2561 2271
rect 2622 2268 2633 2271
rect 2818 2268 2825 2271
rect 2934 2268 2942 2271
rect 2946 2268 2953 2271
rect 3174 2268 3182 2271
rect 3374 2268 3393 2271
rect 3594 2268 3625 2271
rect 4142 2268 4158 2271
rect 4326 2268 4337 2271
rect 4470 2268 4478 2271
rect 4494 2268 4502 2271
rect 4946 2268 4953 2271
rect 166 2261 169 2268
rect 126 2258 145 2261
rect 150 2258 169 2261
rect 318 2258 337 2261
rect 470 2262 473 2268
rect 766 2258 782 2261
rect 862 2258 881 2261
rect 1010 2258 1017 2261
rect 1122 2258 1129 2261
rect 1242 2258 1249 2261
rect 1254 2258 1273 2261
rect 1286 2258 1294 2261
rect 1998 2262 2001 2268
rect 1434 2258 1441 2261
rect 1534 2258 1550 2261
rect 2046 2258 2054 2261
rect 2162 2258 2177 2261
rect 2410 2258 2417 2261
rect 2622 2261 2625 2268
rect 2614 2258 2625 2261
rect 2714 2258 2721 2261
rect 3106 2258 3121 2261
rect 3166 2258 3174 2261
rect 3298 2258 3305 2261
rect 3318 2258 3337 2261
rect 3518 2258 3537 2261
rect 3786 2258 3801 2261
rect 4038 2258 4046 2261
rect 4190 2258 4198 2261
rect 4358 2258 4377 2261
rect 4430 2258 4449 2261
rect 4694 2258 4713 2261
rect 126 2248 129 2258
rect 306 2248 310 2252
rect 318 2248 321 2258
rect 714 2248 718 2252
rect 878 2248 881 2258
rect 890 2248 894 2252
rect 1162 2248 1166 2252
rect 1270 2248 1273 2258
rect 1282 2248 1286 2252
rect 1566 2248 1582 2251
rect 2222 2248 2241 2251
rect 3306 2248 3310 2252
rect 3318 2248 3321 2258
rect 3518 2248 3521 2258
rect 4310 2248 4318 2251
rect 4358 2248 4361 2258
rect 4446 2248 4449 2258
rect 4710 2248 4713 2258
rect 1451 2238 1454 2242
rect 1742 2238 1750 2241
rect 3506 2238 3507 2242
rect 3938 2238 3941 2242
rect 4294 2241 4297 2248
rect 4294 2238 4305 2241
rect 4461 2238 4462 2242
rect 3562 2228 3563 2232
rect 602 2218 603 2222
rect 1130 2218 1131 2222
rect 1962 2218 1963 2222
rect 2066 2218 2067 2222
rect 4277 2218 4278 2222
rect 4725 2218 4726 2222
rect 536 2203 538 2207
rect 542 2203 545 2207
rect 549 2203 552 2207
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1573 2203 1576 2207
rect 2584 2203 2586 2207
rect 2590 2203 2593 2207
rect 2597 2203 2600 2207
rect 3608 2203 3610 2207
rect 3614 2203 3617 2207
rect 3621 2203 3624 2207
rect 4632 2203 4634 2207
rect 4638 2203 4641 2207
rect 4645 2203 4648 2207
rect 685 2188 686 2192
rect 2349 2188 2350 2192
rect 3741 2188 3742 2192
rect 4205 2188 4206 2192
rect 4810 2188 4811 2192
rect 3634 2178 3635 2182
rect 2838 2168 2850 2171
rect 3682 2168 3683 2172
rect 3885 2168 3886 2172
rect 2846 2166 2850 2168
rect 4062 2166 4066 2168
rect 4374 2168 4385 2171
rect 4890 2168 4893 2172
rect 4986 2168 4989 2172
rect 4374 2166 4378 2168
rect 30 2151 34 2153
rect 22 2148 34 2151
rect 246 2151 249 2161
rect 246 2148 265 2151
rect 502 2151 505 2161
rect 502 2148 521 2151
rect 530 2148 569 2151
rect 830 2151 833 2161
rect 830 2148 849 2151
rect 910 2151 913 2158
rect 958 2152 961 2161
rect 1430 2158 1449 2161
rect 902 2148 913 2151
rect 1518 2151 1521 2161
rect 1906 2158 1910 2162
rect 1518 2148 1537 2151
rect 1702 2148 1710 2151
rect 118 2138 130 2141
rect 182 2132 185 2142
rect 534 2138 558 2141
rect 1446 2138 1449 2148
rect 1470 2138 1497 2141
rect 1518 2138 1526 2141
rect 1702 2138 1705 2148
rect 1918 2151 1921 2161
rect 1918 2148 1926 2151
rect 2106 2148 2113 2151
rect 2262 2148 2270 2151
rect 2482 2148 2489 2151
rect 2502 2151 2505 2161
rect 3158 2158 3170 2161
rect 3166 2156 3170 2158
rect 2502 2148 2521 2151
rect 2650 2148 2657 2151
rect 2678 2148 2689 2151
rect 1782 2138 1790 2141
rect 2062 2138 2070 2141
rect 2102 2138 2105 2148
rect 2158 2138 2185 2141
rect 2358 2138 2369 2141
rect 2678 2141 2681 2148
rect 2894 2142 2897 2151
rect 2962 2148 2969 2151
rect 3026 2148 3033 2151
rect 3390 2151 3394 2154
rect 3374 2148 3394 2151
rect 3422 2151 3425 2158
rect 3422 2148 3433 2151
rect 3494 2151 3497 2161
rect 3490 2148 3497 2151
rect 3566 2151 3569 2161
rect 3566 2148 3585 2151
rect 3658 2148 3665 2151
rect 3782 2151 3785 2161
rect 3782 2148 3801 2151
rect 3830 2148 3838 2151
rect 3870 2151 3873 2161
rect 3902 2158 3910 2161
rect 4038 2158 4057 2161
rect 4642 2158 4649 2161
rect 3854 2148 3873 2151
rect 4246 2148 4254 2151
rect 4294 2148 4321 2151
rect 2670 2138 2681 2141
rect 2910 2138 2926 2141
rect 3058 2138 3073 2141
rect 3090 2138 3113 2141
rect 3126 2138 3134 2141
rect 3286 2138 3305 2141
rect 3518 2138 3545 2141
rect 3754 2138 3761 2141
rect 3894 2138 3905 2141
rect 4038 2138 4041 2148
rect 4586 2148 4593 2151
rect 4666 2148 4681 2151
rect 4742 2151 4745 2161
rect 4822 2158 4841 2161
rect 4726 2148 4745 2151
rect 4922 2148 4929 2151
rect 5126 2148 5134 2151
rect 4254 2138 4281 2141
rect 4366 2138 4374 2141
rect 4502 2138 4521 2141
rect 4766 2138 4769 2148
rect 4846 2138 4854 2141
rect 374 2132 378 2133
rect 1798 2131 1802 2133
rect 1790 2128 1802 2131
rect 2382 2131 2386 2133
rect 2374 2128 2386 2131
rect 2838 2132 2842 2133
rect 2878 2128 2897 2131
rect 3114 2128 3118 2132
rect 3286 2128 3289 2138
rect 3918 2131 3922 2133
rect 3910 2128 3922 2131
rect 4398 2131 4402 2136
rect 4398 2128 4414 2131
rect 4502 2128 4505 2138
rect 4870 2131 4874 2133
rect 4862 2128 4874 2131
rect 597 2118 598 2122
rect 1106 2118 1113 2121
rect 1562 2118 1569 2121
rect 1693 2118 1694 2122
rect 1754 2118 1755 2122
rect 3330 2118 3331 2122
rect 1048 2103 1050 2107
rect 1054 2103 1057 2107
rect 1061 2103 1064 2107
rect 2072 2103 2074 2107
rect 2078 2103 2081 2107
rect 2085 2103 2088 2107
rect 3096 2103 3098 2107
rect 3102 2103 3105 2107
rect 3109 2103 3112 2107
rect 4112 2103 4114 2107
rect 4118 2103 4121 2107
rect 4125 2103 4128 2107
rect 813 2088 814 2092
rect 1586 2088 1587 2092
rect 1698 2088 1699 2092
rect 2098 2088 2099 2092
rect 2522 2088 2523 2092
rect 2562 2088 2563 2092
rect 3450 2088 3451 2092
rect 3490 2088 3491 2092
rect 4618 2088 4619 2092
rect 126 2078 145 2081
rect 1634 2078 1635 2082
rect 2694 2078 2705 2081
rect 2974 2078 2985 2081
rect 3238 2078 3249 2081
rect 3390 2078 3409 2081
rect 3822 2078 3833 2081
rect 3838 2078 3857 2081
rect 3918 2078 3937 2081
rect 4102 2078 4121 2081
rect 4358 2078 4369 2081
rect 2694 2077 2698 2078
rect 2974 2077 2978 2078
rect 3238 2077 3242 2078
rect 3822 2077 3826 2078
rect 4358 2077 4362 2078
rect 534 2068 561 2071
rect 742 2068 750 2071
rect 874 2068 882 2071
rect 1142 2068 1150 2071
rect 1222 2068 1233 2071
rect 1670 2068 1697 2071
rect 1754 2068 1761 2071
rect 1774 2068 1782 2071
rect 1938 2068 1953 2071
rect 2054 2068 2086 2071
rect 2374 2068 2382 2071
rect 2446 2068 2457 2071
rect 2546 2068 2561 2071
rect 2574 2068 2590 2071
rect 2986 2068 2993 2071
rect 3014 2068 3030 2071
rect 3590 2068 3618 2071
rect 3730 2068 3738 2071
rect 4138 2068 4153 2071
rect 4262 2068 4274 2071
rect 4374 2068 4382 2071
rect 4550 2071 4553 2081
rect 4558 2078 4577 2081
rect 4766 2078 4777 2081
rect 4830 2078 4842 2081
rect 4966 2078 4985 2081
rect 5062 2078 5081 2081
rect 4766 2077 4770 2078
rect 4838 2077 4842 2078
rect 4546 2068 4553 2071
rect 4814 2068 4825 2071
rect 5178 2068 5185 2071
rect 206 2058 222 2061
rect 790 2058 798 2061
rect 998 2058 1017 2061
rect 1230 2061 1233 2068
rect 1230 2058 1238 2061
rect 1242 2058 1249 2061
rect 1254 2058 1262 2061
rect 1314 2058 1321 2061
rect 1526 2058 1534 2061
rect 1718 2058 1737 2061
rect 1746 2058 1753 2061
rect 1902 2058 1910 2061
rect 1966 2058 1974 2061
rect 2030 2058 2038 2061
rect 2066 2058 2089 2061
rect 2386 2058 2393 2061
rect 2422 2058 2438 2061
rect 2478 2058 2497 2061
rect 2638 2058 2654 2061
rect 2726 2058 2745 2061
rect 2806 2058 2822 2061
rect 3086 2058 3121 2061
rect 3134 2058 3142 2061
rect 3766 2058 3782 2061
rect 4406 2058 4425 2061
rect 4662 2058 4670 2061
rect 5102 2058 5121 2061
rect 5146 2058 5161 2061
rect 5166 2058 5174 2061
rect 474 2048 478 2052
rect 506 2048 510 2052
rect 518 2048 526 2051
rect 718 2048 721 2058
rect 766 2051 769 2058
rect 758 2048 769 2051
rect 998 2048 1001 2058
rect 1046 2048 1081 2051
rect 1262 2048 1273 2051
rect 2742 2048 2745 2058
rect 2866 2048 2870 2052
rect 3118 2048 3121 2058
rect 4406 2048 4409 2058
rect 4462 2048 4481 2051
rect 4518 2048 4537 2051
rect 4658 2048 4662 2052
rect 4802 2048 4806 2052
rect 5118 2048 5121 2058
rect 1270 2042 1273 2048
rect 5030 2042 5034 2044
rect 205 2038 206 2042
rect 442 2038 443 2042
rect 1093 2038 1094 2042
rect 1427 2038 1430 2042
rect 3986 2038 3989 2042
rect 4450 2038 4451 2042
rect 986 2028 987 2032
rect 570 2018 571 2022
rect 2757 2018 2758 2022
rect 2834 2018 2835 2022
rect 3053 2018 3054 2022
rect 536 2003 538 2007
rect 542 2003 545 2007
rect 549 2003 552 2007
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1573 2003 1576 2007
rect 2584 2003 2586 2007
rect 2590 2003 2593 2007
rect 2597 2003 2600 2007
rect 3608 2003 3610 2007
rect 3614 2003 3617 2007
rect 3621 2003 3624 2007
rect 4632 2003 4634 2007
rect 4638 2003 4641 2007
rect 4645 2003 4648 2007
rect 1794 1988 1795 1992
rect 2042 1988 2043 1992
rect 2106 1988 2107 1992
rect 3802 1988 3803 1992
rect 4722 1988 4723 1992
rect 258 1978 259 1982
rect 802 1968 803 1972
rect 1314 1968 1315 1972
rect 2314 1968 2317 1972
rect 3770 1968 3771 1972
rect 4474 1968 4475 1972
rect 4786 1968 4787 1972
rect 3814 1966 3818 1968
rect 270 1951 273 1961
rect 618 1958 622 1962
rect 250 1948 257 1951
rect 270 1948 289 1951
rect 478 1948 494 1951
rect 630 1951 633 1961
rect 630 1948 649 1951
rect 814 1951 817 1961
rect 794 1948 801 1951
rect 814 1948 833 1951
rect 1022 1948 1030 1951
rect 1238 1948 1265 1951
rect 1326 1951 1329 1961
rect 1326 1948 1345 1951
rect 1446 1951 1449 1961
rect 1446 1948 1465 1951
rect 1654 1948 1662 1951
rect 1742 1951 1745 1961
rect 1742 1948 1761 1951
rect 1806 1948 1833 1951
rect 1878 1951 1881 1961
rect 1890 1958 1894 1962
rect 2766 1958 2778 1961
rect 3114 1958 3121 1961
rect 2774 1956 2778 1958
rect 1862 1948 1881 1951
rect 1894 1948 1902 1951
rect 2074 1948 2089 1951
rect 2118 1948 2126 1951
rect 2190 1948 2198 1951
rect 2414 1942 2417 1951
rect 2630 1948 2638 1951
rect 2670 1948 2681 1951
rect 566 1932 569 1942
rect 938 1938 945 1941
rect 1214 1938 1225 1941
rect 1406 1938 1425 1941
rect 1446 1938 1454 1941
rect 1906 1938 1913 1941
rect 2670 1941 2673 1948
rect 2894 1942 2897 1951
rect 3106 1948 3129 1951
rect 3178 1948 3185 1951
rect 2662 1938 2673 1941
rect 3142 1938 3150 1941
rect 3230 1941 3233 1948
rect 3398 1951 3401 1961
rect 3822 1958 3830 1961
rect 3906 1958 3910 1962
rect 3398 1948 3417 1951
rect 3522 1948 3529 1951
rect 3562 1948 3569 1951
rect 3598 1948 3622 1951
rect 3694 1948 3705 1951
rect 3754 1948 3761 1951
rect 3910 1948 3918 1951
rect 3230 1938 3241 1941
rect 3702 1941 3705 1948
rect 4022 1951 4025 1958
rect 4022 1948 4033 1951
rect 4210 1948 4217 1951
rect 4230 1951 4233 1961
rect 4230 1948 4249 1951
rect 4438 1951 4441 1958
rect 4438 1948 4449 1951
rect 4486 1951 4489 1961
rect 4658 1958 4662 1962
rect 4486 1948 4505 1951
rect 4670 1951 4673 1961
rect 4798 1958 4817 1961
rect 4670 1948 4689 1951
rect 4854 1951 4857 1961
rect 4866 1958 4870 1962
rect 4838 1948 4857 1951
rect 3702 1938 3721 1941
rect 4062 1938 4081 1941
rect 4202 1938 4209 1941
rect 4642 1938 4649 1941
rect 4878 1938 4889 1941
rect 414 1928 433 1931
rect 2398 1928 2417 1931
rect 2469 1928 2470 1932
rect 2878 1928 2897 1931
rect 2934 1928 2953 1931
rect 3254 1931 3258 1933
rect 3246 1928 3258 1931
rect 3558 1928 3561 1938
rect 4014 1931 4018 1933
rect 4014 1928 4025 1931
rect 4062 1928 4065 1938
rect 4178 1928 4179 1932
rect 4534 1931 4538 1933
rect 4902 1931 4906 1933
rect 5022 1931 5026 1933
rect 4526 1928 4538 1931
rect 4894 1928 4906 1931
rect 5014 1928 5026 1931
rect 5142 1928 5161 1931
rect 973 1918 974 1922
rect 1277 1918 1278 1922
rect 1618 1918 1625 1921
rect 2573 1918 2574 1922
rect 2989 1918 2990 1922
rect 1048 1903 1050 1907
rect 1054 1903 1057 1907
rect 1061 1903 1064 1907
rect 2072 1903 2074 1907
rect 2078 1903 2081 1907
rect 2085 1903 2088 1907
rect 3096 1903 3098 1907
rect 3102 1903 3105 1907
rect 3109 1903 3112 1907
rect 4112 1903 4114 1907
rect 4118 1903 4121 1907
rect 4125 1903 4128 1907
rect 1834 1888 1835 1892
rect 1901 1888 1902 1892
rect 3605 1888 3606 1892
rect 4546 1888 4547 1892
rect 4638 1888 4649 1891
rect 5182 1888 5190 1891
rect 598 1878 610 1881
rect 934 1878 945 1881
rect 1694 1878 1705 1881
rect 2326 1878 2337 1881
rect 2502 1878 2514 1881
rect 2878 1878 2897 1881
rect 3294 1878 3305 1881
rect 3550 1878 3569 1881
rect 3678 1878 3690 1881
rect 4638 1881 4641 1888
rect 4622 1878 4641 1881
rect 4806 1878 4825 1881
rect 5070 1878 5081 1881
rect 606 1877 610 1878
rect 934 1877 938 1878
rect 1694 1877 1698 1878
rect 2326 1877 2330 1878
rect 2510 1877 2514 1878
rect 3294 1877 3298 1878
rect 3686 1877 3690 1878
rect 5070 1877 5074 1878
rect 5166 1874 5170 1878
rect 230 1858 249 1861
rect 414 1858 433 1861
rect 566 1858 574 1861
rect 702 1862 705 1871
rect 950 1868 961 1871
rect 1454 1868 1465 1871
rect 1710 1868 1721 1871
rect 2342 1868 2353 1871
rect 2486 1868 2497 1871
rect 3114 1868 3121 1871
rect 3146 1868 3153 1871
rect 3310 1868 3321 1871
rect 4106 1868 4113 1871
rect 718 1858 726 1861
rect 754 1858 761 1861
rect 974 1858 982 1861
rect 1038 1858 1073 1861
rect 1154 1858 1161 1861
rect 1214 1858 1222 1861
rect 2350 1862 2353 1868
rect 1510 1858 1518 1861
rect 1742 1858 1761 1861
rect 1862 1858 1889 1861
rect 2046 1858 2054 1861
rect 2078 1858 2102 1861
rect 2206 1858 2225 1861
rect 2374 1858 2393 1861
rect 2446 1858 2465 1861
rect 2478 1858 2486 1861
rect 2942 1858 2950 1861
rect 3014 1858 3022 1861
rect 3086 1858 3121 1861
rect 3310 1858 3318 1861
rect 3642 1858 3649 1861
rect 3654 1858 3662 1861
rect 4014 1858 4022 1861
rect 4078 1858 4086 1861
rect 4386 1858 4393 1861
rect 4434 1858 4441 1861
rect 4454 1858 4473 1861
rect 5126 1858 5134 1861
rect 246 1848 249 1858
rect 414 1848 417 1858
rect 1046 1848 1062 1851
rect 1070 1848 1073 1858
rect 1242 1848 1246 1852
rect 1742 1848 1745 1858
rect 2206 1848 2209 1858
rect 2374 1848 2377 1858
rect 2462 1848 2465 1858
rect 2474 1848 2478 1852
rect 2782 1851 2786 1854
rect 2782 1848 2793 1851
rect 3070 1848 3078 1851
rect 3118 1848 3121 1858
rect 3174 1848 3193 1851
rect 4126 1848 4145 1851
rect 4454 1848 4457 1858
rect 1838 1842 1842 1844
rect 3038 1842 3042 1844
rect 3198 1842 3202 1844
rect 4142 1842 4145 1848
rect 946 1838 953 1841
rect 2307 1838 2310 1842
rect 4114 1838 4121 1841
rect 4573 1838 4574 1842
rect 4754 1838 4755 1842
rect 5051 1838 5054 1842
rect 762 1818 763 1822
rect 1005 1818 1006 1822
rect 4506 1818 4507 1822
rect 536 1803 538 1807
rect 542 1803 545 1807
rect 549 1803 552 1807
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1573 1803 1576 1807
rect 2584 1803 2586 1807
rect 2590 1803 2593 1807
rect 2597 1803 2600 1807
rect 3608 1803 3610 1807
rect 3614 1803 3617 1807
rect 3621 1803 3624 1807
rect 4632 1803 4634 1807
rect 4638 1803 4641 1807
rect 4645 1803 4648 1807
rect 1173 1788 1174 1792
rect 1221 1788 1222 1792
rect 1938 1788 1939 1792
rect 2250 1788 2251 1792
rect 2450 1788 2451 1792
rect 2746 1788 2747 1792
rect 2933 1788 2934 1792
rect 3581 1788 3582 1792
rect 4282 1788 4283 1792
rect 4322 1788 4323 1792
rect 5101 1788 5102 1792
rect 5186 1788 5187 1792
rect 3418 1778 3419 1782
rect 4642 1778 4649 1781
rect 299 1768 302 1772
rect 1322 1768 1325 1772
rect 1486 1768 1497 1771
rect 3053 1768 3054 1772
rect 4773 1768 4774 1772
rect 338 1758 342 1762
rect 206 1741 209 1751
rect 350 1751 353 1761
rect 546 1758 561 1761
rect 710 1761 713 1768
rect 1486 1766 1490 1768
rect 702 1758 713 1761
rect 330 1748 337 1751
rect 350 1748 369 1751
rect 422 1748 430 1751
rect 614 1748 622 1751
rect 194 1738 209 1741
rect 686 1741 689 1748
rect 678 1738 689 1741
rect 742 1738 745 1748
rect 1074 1748 1097 1751
rect 1190 1748 1198 1751
rect 1774 1751 1777 1761
rect 2410 1758 2414 1762
rect 1758 1748 1777 1751
rect 1866 1748 1881 1751
rect 1950 1748 1958 1751
rect 2166 1748 2177 1751
rect 2226 1748 2233 1751
rect 2322 1748 2337 1751
rect 2478 1751 2481 1761
rect 2786 1758 2790 1762
rect 2906 1758 2913 1761
rect 3442 1758 3446 1762
rect 2474 1748 2481 1751
rect 2758 1748 2774 1751
rect 2838 1748 2854 1751
rect 3150 1748 3161 1751
rect 3178 1748 3185 1751
rect 854 1738 865 1741
rect 1274 1738 1281 1741
rect 1490 1738 1498 1741
rect 1718 1738 1721 1748
rect 1802 1738 1809 1741
rect 2166 1741 2169 1748
rect 3374 1742 3377 1751
rect 3582 1748 3590 1751
rect 3774 1751 3777 1761
rect 4038 1752 4041 1761
rect 3774 1748 3793 1751
rect 4226 1748 4233 1751
rect 4274 1748 4281 1751
rect 4446 1751 4449 1761
rect 4458 1758 4462 1762
rect 4430 1748 4449 1751
rect 4598 1751 4601 1761
rect 4802 1758 4806 1762
rect 4582 1748 4601 1751
rect 4774 1748 4790 1751
rect 5086 1751 5089 1761
rect 5070 1748 5089 1751
rect 2162 1738 2169 1741
rect 2946 1738 2953 1741
rect 2986 1738 2993 1741
rect 3102 1738 3134 1741
rect 3250 1738 3257 1741
rect 3590 1738 3601 1741
rect 3842 1738 3849 1741
rect 4006 1738 4025 1741
rect 4262 1738 4273 1741
rect 4398 1738 4406 1741
rect 4622 1738 4649 1741
rect 4934 1738 4937 1748
rect 5110 1738 5118 1741
rect 210 1728 217 1731
rect 510 1728 529 1731
rect 534 1728 542 1731
rect 838 1731 842 1733
rect 838 1728 849 1731
rect 1278 1728 1281 1738
rect 1494 1736 1498 1738
rect 1286 1728 1294 1731
rect 1422 1728 1441 1731
rect 1622 1731 1626 1733
rect 1822 1731 1826 1733
rect 1614 1728 1626 1731
rect 1814 1728 1826 1731
rect 2582 1728 2601 1731
rect 2894 1731 2898 1733
rect 2894 1728 2905 1731
rect 3006 1728 3025 1731
rect 3130 1728 3137 1731
rect 3230 1728 3249 1731
rect 4006 1728 4009 1738
rect 4198 1731 4202 1733
rect 4034 1728 4046 1731
rect 4198 1728 4209 1731
rect 4662 1731 4666 1733
rect 4654 1728 4666 1731
rect 5126 1728 5145 1731
rect 565 1718 566 1722
rect 1062 1718 1070 1721
rect 2598 1721 2601 1728
rect 2598 1718 2609 1721
rect 1048 1703 1050 1707
rect 1054 1703 1057 1707
rect 1061 1703 1064 1707
rect 2072 1703 2074 1707
rect 2078 1703 2081 1707
rect 2085 1703 2088 1707
rect 3096 1703 3098 1707
rect 3102 1703 3105 1707
rect 3109 1703 3112 1707
rect 4112 1703 4114 1707
rect 4118 1703 4121 1707
rect 4125 1703 4128 1707
rect 765 1688 766 1692
rect 1029 1688 1030 1692
rect 1525 1688 1526 1692
rect 1834 1688 1835 1692
rect 2861 1688 2862 1692
rect 3037 1688 3038 1692
rect 3397 1688 3398 1692
rect 3981 1688 3982 1692
rect 4474 1688 4475 1692
rect 4898 1688 4899 1692
rect 102 1678 121 1681
rect 318 1678 329 1681
rect 806 1678 825 1681
rect 1278 1678 1297 1681
rect 1654 1678 1665 1681
rect 318 1677 322 1678
rect 1654 1677 1658 1678
rect 330 1668 337 1671
rect 526 1668 553 1671
rect 606 1662 609 1671
rect 774 1668 782 1671
rect 834 1668 842 1671
rect 1058 1668 1073 1671
rect 1194 1668 1201 1671
rect 1466 1668 1473 1671
rect 1730 1668 1737 1671
rect 1798 1668 1806 1671
rect 1910 1671 1913 1681
rect 1894 1668 1913 1671
rect 1990 1668 1998 1671
rect 2070 1668 2086 1671
rect 2118 1668 2129 1671
rect 2206 1671 2209 1681
rect 2246 1678 2258 1681
rect 4650 1678 4657 1681
rect 4782 1678 4794 1681
rect 5086 1678 5098 1681
rect 2254 1677 2258 1678
rect 4790 1677 4794 1678
rect 4974 1674 4978 1678
rect 5094 1677 5098 1678
rect 2190 1668 2209 1671
rect 2758 1668 2777 1671
rect 3382 1668 3390 1671
rect 3422 1668 3433 1671
rect 3710 1668 3721 1671
rect 4026 1668 4033 1671
rect 4054 1668 4062 1671
rect 4334 1668 4345 1671
rect 4766 1668 4777 1671
rect 166 1658 182 1661
rect 462 1658 481 1661
rect 630 1658 646 1661
rect 806 1658 809 1668
rect 2126 1662 2129 1668
rect 1006 1658 1014 1661
rect 1442 1658 1449 1661
rect 1486 1658 1494 1661
rect 1686 1658 1705 1661
rect 1762 1658 1769 1661
rect 1966 1658 1974 1661
rect 2082 1658 2105 1661
rect 2178 1658 2185 1661
rect 2354 1658 2361 1661
rect 2670 1658 2678 1661
rect 2982 1658 3001 1661
rect 3122 1658 3145 1661
rect 3150 1658 3166 1661
rect 3578 1658 3585 1661
rect 3598 1658 3633 1661
rect 3738 1658 3745 1661
rect 3830 1658 3849 1661
rect 4174 1658 4201 1661
rect 4238 1658 4257 1661
rect 4270 1658 4286 1661
rect 4342 1661 4345 1668
rect 4766 1662 4769 1668
rect 4342 1658 4350 1661
rect 4578 1658 4585 1661
rect 4622 1658 4646 1661
rect 4650 1658 4654 1661
rect 4726 1658 4745 1661
rect 450 1648 454 1652
rect 462 1648 465 1658
rect 1222 1648 1241 1651
rect 1702 1648 1705 1658
rect 2998 1648 3001 1658
rect 3190 1651 3194 1654
rect 3182 1648 3194 1651
rect 3586 1648 3590 1652
rect 3598 1648 3601 1658
rect 3610 1648 3625 1651
rect 3846 1648 3849 1658
rect 3966 1651 3970 1654
rect 3966 1648 3977 1651
rect 4254 1648 4257 1658
rect 4742 1648 4745 1658
rect 4754 1648 4758 1652
rect 2854 1642 2858 1644
rect 1147 1638 1150 1642
rect 2362 1638 2363 1642
rect 3301 1638 3302 1642
rect 3730 1638 3738 1641
rect 4162 1638 4163 1642
rect 4941 1638 4942 1642
rect 3013 1618 3014 1622
rect 3789 1618 3790 1622
rect 4269 1618 4270 1622
rect 536 1603 538 1607
rect 542 1603 545 1607
rect 549 1603 552 1607
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1573 1603 1576 1607
rect 2584 1603 2586 1607
rect 2590 1603 2593 1607
rect 2597 1603 2600 1607
rect 3608 1603 3610 1607
rect 3614 1603 3617 1607
rect 3621 1603 3624 1607
rect 4632 1603 4634 1607
rect 4638 1603 4641 1607
rect 4645 1603 4648 1607
rect 290 1588 291 1592
rect 370 1588 371 1592
rect 1173 1588 1174 1592
rect 1773 1588 1774 1592
rect 1922 1588 1923 1592
rect 2021 1588 2022 1592
rect 2069 1588 2070 1592
rect 2181 1588 2182 1592
rect 2941 1588 2942 1592
rect 2989 1588 2990 1592
rect 3205 1588 3206 1592
rect 3837 1588 3838 1592
rect 4109 1588 4110 1592
rect 4378 1588 4379 1592
rect 1434 1578 1435 1582
rect 2290 1578 2291 1582
rect 3333 1578 3334 1582
rect 3573 1578 3574 1582
rect 547 1568 550 1572
rect 1214 1566 1218 1568
rect 4898 1568 4901 1572
rect 1334 1566 1338 1568
rect 302 1551 305 1561
rect 566 1558 593 1561
rect 1334 1558 1345 1561
rect 1354 1558 1358 1562
rect 1490 1558 1494 1562
rect 1966 1558 1985 1561
rect 3362 1558 3366 1562
rect 566 1556 570 1558
rect 282 1548 289 1551
rect 302 1548 321 1551
rect 1254 1548 1262 1551
rect 1390 1548 1398 1551
rect 1426 1548 1433 1551
rect 1494 1548 1502 1551
rect 1686 1548 1694 1551
rect 1958 1548 1966 1551
rect 2114 1548 2121 1551
rect 2162 1548 2169 1551
rect 2210 1548 2217 1551
rect 2638 1548 2646 1551
rect 2798 1548 2825 1551
rect 2854 1548 2862 1551
rect 2870 1548 2889 1551
rect 2974 1548 2982 1551
rect 3022 1548 3041 1551
rect 3090 1548 3105 1551
rect 3334 1548 3342 1551
rect 3374 1551 3377 1561
rect 3526 1552 3529 1561
rect 3538 1558 3542 1562
rect 3794 1558 3798 1562
rect 3878 1558 3905 1561
rect 3374 1548 3393 1551
rect 350 1538 361 1541
rect 394 1538 401 1541
rect 426 1538 433 1541
rect 886 1538 894 1541
rect 918 1538 926 1541
rect 1122 1538 1129 1541
rect 1374 1538 1377 1548
rect 1414 1538 1425 1541
rect 1502 1538 1513 1541
rect 1642 1538 1649 1541
rect 1802 1538 1809 1541
rect 1902 1541 1905 1548
rect 3574 1548 3582 1551
rect 3786 1548 3793 1551
rect 4070 1548 4078 1551
rect 4126 1548 4134 1551
rect 4142 1548 4161 1551
rect 1902 1538 1913 1541
rect 2378 1538 2385 1541
rect 3590 1541 3593 1548
rect 3590 1538 3601 1541
rect 3774 1538 3785 1541
rect 3862 1538 3865 1548
rect 3918 1538 3921 1548
rect 4142 1542 4145 1548
rect 4294 1548 4310 1551
rect 4342 1548 4350 1551
rect 4654 1551 4657 1561
rect 4666 1558 4670 1562
rect 4622 1548 4657 1551
rect 5030 1551 5033 1561
rect 5026 1548 5033 1551
rect 5058 1548 5065 1551
rect 5070 1548 5078 1551
rect 5154 1548 5161 1551
rect 3930 1538 3937 1541
rect 4318 1538 4329 1541
rect 4790 1538 4801 1541
rect 5086 1538 5094 1541
rect 126 1528 145 1531
rect 246 1531 250 1533
rect 246 1528 257 1531
rect 446 1528 465 1531
rect 894 1528 913 1531
rect 918 1528 921 1538
rect 973 1528 974 1532
rect 1549 1528 1550 1532
rect 2133 1528 2134 1532
rect 2590 1528 2609 1531
rect 4518 1531 4522 1533
rect 4510 1528 4522 1531
rect 4774 1531 4778 1533
rect 4878 1531 4882 1533
rect 4774 1528 4785 1531
rect 4870 1528 4882 1531
rect 4998 1528 5017 1531
rect 5102 1531 5106 1533
rect 5094 1528 5106 1531
rect 2590 1521 2593 1528
rect 2582 1518 2593 1521
rect 2869 1518 2870 1522
rect 3909 1518 3910 1522
rect 1048 1503 1050 1507
rect 1054 1503 1057 1507
rect 1061 1503 1064 1507
rect 2072 1503 2074 1507
rect 2078 1503 2081 1507
rect 2085 1503 2088 1507
rect 3096 1503 3098 1507
rect 3102 1503 3105 1507
rect 3109 1503 3112 1507
rect 4112 1503 4114 1507
rect 4118 1503 4121 1507
rect 4125 1503 4128 1507
rect 669 1488 670 1492
rect 749 1488 750 1492
rect 778 1488 779 1492
rect 1690 1488 1691 1492
rect 1938 1488 1939 1492
rect 2642 1488 2643 1492
rect 3029 1488 3030 1492
rect 3086 1488 3105 1491
rect 3450 1488 3451 1492
rect 3674 1488 3675 1492
rect 3698 1488 3699 1492
rect 3850 1488 3851 1492
rect 3970 1488 3971 1492
rect 4106 1488 4107 1492
rect 4770 1488 4771 1492
rect 3102 1482 3105 1488
rect 222 1471 225 1481
rect 710 1478 729 1481
rect 2286 1478 2298 1481
rect 2942 1478 2961 1481
rect 3990 1478 4002 1481
rect 574 1477 578 1478
rect 2294 1477 2298 1478
rect 3998 1477 4002 1478
rect 4222 1478 4233 1481
rect 4222 1477 4226 1478
rect 206 1468 225 1471
rect 414 1468 425 1471
rect 1142 1468 1150 1471
rect 2070 1468 2086 1471
rect 2238 1468 2246 1471
rect 3098 1468 3110 1471
rect 3142 1468 3150 1471
rect 126 1458 145 1461
rect 622 1458 641 1461
rect 806 1458 814 1461
rect 1102 1458 1121 1461
rect 1190 1458 1198 1461
rect 1326 1458 1334 1461
rect 1450 1458 1457 1461
rect 1614 1458 1630 1461
rect 1706 1458 1713 1461
rect 2142 1458 2150 1461
rect 2174 1458 2190 1461
rect 2230 1458 2246 1461
rect 2338 1458 2353 1461
rect 2750 1458 2766 1461
rect 3014 1458 3022 1461
rect 3062 1458 3081 1461
rect 3126 1458 3145 1461
rect 3162 1458 3169 1461
rect 3406 1462 3409 1471
rect 4374 1471 4377 1481
rect 4702 1478 4721 1481
rect 4358 1468 4377 1471
rect 4962 1468 4970 1471
rect 5018 1468 5019 1472
rect 3486 1458 3505 1461
rect 3598 1458 3622 1461
rect 3898 1458 3905 1461
rect 4526 1458 4545 1461
rect 5146 1458 5153 1461
rect 126 1448 129 1458
rect 622 1448 625 1458
rect 910 1451 914 1454
rect 910 1448 921 1451
rect 1118 1448 1121 1458
rect 1158 1448 1177 1451
rect 1438 1448 1449 1451
rect 2138 1448 2142 1452
rect 3086 1448 3094 1451
rect 3254 1451 3258 1454
rect 3246 1448 3258 1451
rect 3386 1448 3390 1452
rect 3486 1448 3489 1458
rect 3562 1448 3566 1452
rect 3734 1448 3737 1458
rect 3918 1448 3921 1458
rect 4110 1448 4118 1451
rect 4330 1448 4334 1452
rect 4526 1448 4529 1458
rect 4810 1448 4814 1452
rect 4858 1448 4865 1451
rect 934 1441 937 1448
rect 1238 1442 1242 1444
rect 1438 1442 1442 1444
rect 3366 1442 3370 1444
rect 4870 1442 4874 1444
rect 926 1438 937 1441
rect 2314 1438 2317 1442
rect 3734 1438 3745 1441
rect 3906 1438 3907 1442
rect 4578 1438 4581 1442
rect 466 1418 467 1422
rect 1514 1418 1515 1422
rect 3213 1418 3214 1422
rect 3474 1418 3475 1422
rect 3597 1418 3598 1422
rect 3722 1418 3723 1422
rect 3941 1418 3942 1422
rect 536 1403 538 1407
rect 542 1403 545 1407
rect 549 1403 552 1407
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1573 1403 1576 1407
rect 2584 1403 2586 1407
rect 2590 1403 2593 1407
rect 2597 1403 2600 1407
rect 3608 1403 3610 1407
rect 3614 1403 3617 1407
rect 3621 1403 3624 1407
rect 4632 1403 4634 1407
rect 4638 1403 4641 1407
rect 4645 1403 4648 1407
rect 565 1388 566 1392
rect 810 1388 811 1392
rect 1013 1388 1014 1392
rect 1365 1388 1366 1392
rect 1642 1388 1643 1392
rect 2658 1388 2659 1392
rect 3813 1388 3814 1392
rect 290 1368 291 1372
rect 822 1368 830 1371
rect 1098 1368 1099 1372
rect 2478 1368 2486 1371
rect 3930 1368 3933 1372
rect 4619 1368 4622 1372
rect 38 1348 46 1351
rect 106 1348 113 1351
rect 138 1348 145 1351
rect 214 1348 222 1351
rect 302 1351 305 1361
rect 302 1348 321 1351
rect 366 1351 369 1361
rect 594 1358 598 1362
rect 366 1348 385 1351
rect 422 1348 430 1351
rect 622 1351 625 1358
rect 614 1348 625 1351
rect 662 1348 670 1351
rect 750 1351 753 1361
rect 870 1361 873 1368
rect 862 1358 873 1361
rect 1534 1358 1545 1361
rect 1842 1358 1846 1362
rect 2306 1358 2310 1362
rect 1534 1356 1538 1358
rect 3438 1352 3441 1361
rect 3666 1358 3670 1362
rect 3890 1358 3894 1362
rect 750 1348 769 1351
rect 1058 1348 1065 1351
rect 158 1338 166 1341
rect 606 1338 617 1341
rect 882 1338 889 1341
rect 1078 1338 1081 1348
rect 1430 1348 1438 1351
rect 1498 1348 1505 1351
rect 1658 1348 1673 1351
rect 1714 1348 1721 1351
rect 1730 1348 1742 1351
rect 2074 1348 2097 1351
rect 2102 1348 2110 1351
rect 2150 1348 2158 1351
rect 2218 1348 2225 1351
rect 2230 1348 2238 1351
rect 2310 1348 2318 1351
rect 2582 1348 2590 1351
rect 2786 1348 2801 1351
rect 2854 1348 2862 1351
rect 3158 1348 3169 1351
rect 3254 1348 3273 1351
rect 1782 1338 1790 1341
rect 1798 1338 1801 1348
rect 2238 1338 2265 1341
rect 2350 1341 2353 1348
rect 3814 1348 3822 1351
rect 3894 1348 3902 1351
rect 4174 1351 4177 1361
rect 4186 1358 4190 1362
rect 4158 1348 4177 1351
rect 4246 1351 4249 1361
rect 4674 1358 4678 1362
rect 4246 1348 4265 1351
rect 2350 1338 2361 1341
rect 2582 1338 2606 1341
rect 3138 1338 3145 1341
rect 3222 1338 3241 1341
rect 3630 1338 3646 1341
rect 3678 1338 3689 1341
rect 4206 1341 4209 1348
rect 4822 1348 4830 1351
rect 4898 1348 4913 1351
rect 5038 1351 5041 1358
rect 5030 1348 5041 1351
rect 5058 1348 5065 1351
rect 5118 1348 5126 1351
rect 4206 1338 4225 1341
rect 4658 1338 4665 1341
rect 4806 1338 4809 1348
rect 4954 1338 4961 1341
rect 4974 1338 4993 1341
rect 5034 1338 5041 1341
rect 1942 1336 1946 1338
rect 630 1331 634 1333
rect 622 1328 634 1331
rect 2374 1331 2378 1333
rect 2366 1328 2378 1331
rect 2502 1328 2521 1331
rect 2694 1328 2713 1331
rect 3158 1328 3166 1331
rect 3238 1328 3241 1338
rect 3438 1332 3441 1338
rect 3434 1328 3441 1332
rect 3702 1331 3706 1333
rect 3694 1328 3706 1331
rect 4478 1328 4497 1331
rect 4854 1331 4858 1333
rect 4846 1328 4858 1331
rect 4974 1328 4977 1338
rect 5062 1331 5065 1338
rect 5086 1331 5090 1333
rect 5062 1328 5073 1331
rect 5078 1328 5090 1331
rect 1325 1318 1326 1322
rect 2621 1318 2622 1322
rect 5050 1318 5051 1322
rect 1048 1303 1050 1307
rect 1054 1303 1057 1307
rect 1061 1303 1064 1307
rect 2072 1303 2074 1307
rect 2078 1303 2081 1307
rect 2085 1303 2088 1307
rect 3096 1303 3098 1307
rect 3102 1303 3105 1307
rect 3109 1303 3112 1307
rect 4112 1303 4114 1307
rect 4118 1303 4121 1307
rect 4125 1303 4128 1307
rect 437 1288 438 1292
rect 1189 1288 1190 1292
rect 1994 1288 1995 1292
rect 2202 1288 2203 1292
rect 3086 1288 3097 1291
rect 4274 1288 4275 1292
rect 4714 1288 4715 1292
rect 4738 1288 4739 1292
rect 4762 1288 4763 1292
rect 4786 1288 4787 1292
rect 458 1278 462 1282
rect 670 1271 673 1281
rect 1578 1278 1593 1281
rect 1598 1278 1617 1281
rect 894 1276 898 1278
rect 670 1268 689 1271
rect 126 1258 145 1261
rect 222 1261 225 1268
rect 206 1258 225 1261
rect 394 1258 409 1261
rect 614 1258 633 1261
rect 822 1262 825 1271
rect 1074 1268 1081 1271
rect 1618 1268 1625 1271
rect 1702 1271 1705 1281
rect 1702 1268 1721 1271
rect 1822 1268 1834 1271
rect 1950 1271 1953 1281
rect 3094 1281 3097 1288
rect 1930 1268 1937 1271
rect 1950 1268 1969 1271
rect 2349 1268 2350 1272
rect 2614 1271 2617 1281
rect 3094 1278 3113 1281
rect 3350 1278 3369 1281
rect 4310 1278 4329 1281
rect 4642 1278 4657 1281
rect 2582 1268 2617 1271
rect 3106 1268 3121 1271
rect 3238 1268 3246 1271
rect 3398 1268 3409 1271
rect 4029 1268 4030 1272
rect 4382 1268 4409 1271
rect 4630 1268 4673 1271
rect 4770 1268 4777 1271
rect 4933 1268 4934 1272
rect 5070 1268 5081 1271
rect 1138 1258 1145 1261
rect 1150 1258 1166 1261
rect 1182 1261 1185 1268
rect 1174 1258 1185 1261
rect 1290 1258 1297 1261
rect 1366 1258 1382 1261
rect 1702 1258 1710 1261
rect 2270 1258 2289 1261
rect 2530 1258 2537 1261
rect 2906 1258 2913 1261
rect 2950 1258 2969 1261
rect 2982 1258 2990 1261
rect 3406 1262 3409 1268
rect 3118 1258 3137 1261
rect 3194 1258 3201 1261
rect 3446 1258 3457 1261
rect 3526 1258 3534 1261
rect 3890 1258 3905 1261
rect 3954 1258 3961 1261
rect 4286 1258 4294 1261
rect 4590 1258 4609 1261
rect 5074 1258 5081 1261
rect 114 1248 118 1252
rect 126 1248 129 1258
rect 174 1248 193 1251
rect 422 1248 433 1251
rect 614 1248 617 1258
rect 834 1248 838 1252
rect 1114 1248 1118 1252
rect 1374 1248 1393 1251
rect 2014 1248 2033 1251
rect 2162 1248 2169 1251
rect 2270 1248 2273 1258
rect 2610 1248 2617 1251
rect 2966 1248 2969 1258
rect 3446 1252 3449 1258
rect 3242 1248 3249 1251
rect 3474 1248 3481 1251
rect 3602 1248 3606 1252
rect 3694 1248 3713 1251
rect 4430 1248 4449 1251
rect 4606 1248 4609 1258
rect 5058 1248 5062 1252
rect 430 1242 434 1244
rect 410 1238 411 1242
rect 1454 1242 1458 1244
rect 3462 1242 3466 1244
rect 2453 1238 2454 1242
rect 3181 1238 3182 1242
rect 3205 1238 3206 1242
rect 3486 1241 3490 1244
rect 3686 1242 3690 1244
rect 4478 1242 4482 1244
rect 3486 1238 3497 1241
rect 3725 1238 3726 1242
rect 4010 1238 4013 1242
rect 4718 1241 4722 1244
rect 4718 1238 4726 1241
rect 4766 1241 4770 1244
rect 4790 1242 4794 1244
rect 4766 1238 4774 1241
rect 4818 1238 4821 1242
rect 378 1218 379 1222
rect 4682 1218 4683 1222
rect 536 1203 538 1207
rect 542 1203 545 1207
rect 549 1203 552 1207
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1573 1203 1576 1207
rect 2584 1203 2586 1207
rect 2590 1203 2593 1207
rect 2597 1203 2600 1207
rect 3608 1203 3610 1207
rect 3614 1203 3617 1207
rect 3621 1203 3624 1207
rect 4632 1203 4634 1207
rect 4638 1203 4641 1207
rect 4645 1203 4648 1207
rect 877 1188 878 1192
rect 1010 1188 1011 1192
rect 1242 1188 1243 1192
rect 1426 1188 1427 1192
rect 1698 1188 1699 1192
rect 2714 1188 2715 1192
rect 3197 1188 3198 1192
rect 3685 1188 3686 1192
rect 3853 1188 3854 1192
rect 4082 1188 4083 1192
rect 4386 1188 4387 1192
rect 4666 1188 4667 1192
rect 166 1168 178 1171
rect 606 1168 614 1171
rect 746 1168 747 1172
rect 781 1168 782 1172
rect 1805 1168 1806 1172
rect 2134 1168 2145 1171
rect 2462 1168 2473 1171
rect 3078 1168 3090 1171
rect 186 1158 190 1162
rect 594 1158 598 1162
rect 766 1152 769 1161
rect 1458 1158 1462 1162
rect 578 1148 593 1151
rect 610 1148 617 1151
rect 670 1148 678 1151
rect 690 1148 697 1151
rect 782 1148 798 1151
rect 858 1148 865 1151
rect 926 1148 934 1151
rect 1542 1151 1545 1161
rect 1554 1158 1558 1162
rect 1710 1158 1729 1161
rect 1526 1148 1545 1151
rect 1862 1151 1865 1161
rect 2122 1158 2126 1162
rect 2426 1158 2430 1162
rect 2446 1161 2449 1168
rect 2462 1166 2466 1168
rect 3086 1166 3090 1168
rect 2438 1158 2449 1161
rect 3094 1158 3129 1161
rect 3506 1158 3510 1162
rect 2158 1153 2162 1158
rect 1862 1148 1881 1151
rect 1886 1148 1902 1151
rect 2194 1148 2201 1151
rect 2502 1148 2510 1151
rect 2850 1148 2865 1151
rect 250 1138 265 1141
rect 614 1138 617 1148
rect 826 1138 833 1141
rect 1406 1138 1417 1141
rect 1478 1138 1481 1148
rect 1814 1138 1825 1141
rect 2102 1138 2105 1148
rect 2278 1141 2281 1148
rect 3142 1148 3150 1151
rect 3178 1148 3185 1151
rect 3226 1148 3233 1151
rect 3518 1151 3521 1161
rect 3742 1161 3745 1168
rect 3734 1158 3745 1161
rect 4210 1158 4214 1162
rect 3518 1148 3537 1151
rect 3702 1148 3710 1151
rect 3766 1148 3774 1151
rect 3894 1148 3902 1151
rect 3986 1148 4001 1151
rect 4058 1148 4065 1151
rect 4146 1148 4153 1151
rect 4182 1148 4190 1151
rect 4410 1148 4417 1151
rect 4498 1148 4505 1151
rect 4522 1148 4529 1151
rect 4558 1148 4585 1151
rect 4614 1148 4638 1151
rect 2270 1138 2281 1141
rect 2598 1138 2606 1141
rect 2646 1138 2654 1141
rect 2894 1138 2902 1141
rect 3646 1138 3662 1141
rect 3786 1138 3793 1141
rect 4106 1138 4121 1141
rect 4226 1138 4233 1141
rect 4598 1138 4601 1148
rect 4918 1142 4921 1151
rect 4998 1148 5006 1151
rect 4718 1138 4729 1141
rect 4950 1138 4969 1141
rect 4982 1138 4985 1148
rect 2758 1128 2777 1131
rect 2958 1128 2977 1131
rect 3062 1131 3066 1136
rect 3050 1128 3066 1131
rect 3566 1128 3585 1131
rect 4170 1128 4171 1132
rect 4246 1131 4250 1133
rect 4238 1128 4250 1131
rect 4438 1128 4457 1131
rect 4546 1128 4547 1132
rect 4742 1131 4746 1133
rect 4734 1128 4746 1131
rect 4846 1128 4865 1131
rect 4950 1128 4953 1138
rect 5030 1131 5034 1133
rect 5022 1128 5034 1131
rect 805 1118 806 1122
rect 4349 1118 4350 1122
rect 4477 1118 4478 1122
rect 1048 1103 1050 1107
rect 1054 1103 1057 1107
rect 1061 1103 1064 1107
rect 2072 1103 2074 1107
rect 2078 1103 2081 1107
rect 2085 1103 2088 1107
rect 3096 1103 3098 1107
rect 3102 1103 3105 1107
rect 3109 1103 3112 1107
rect 4112 1103 4114 1107
rect 4118 1103 4121 1107
rect 4125 1103 4128 1107
rect 1013 1088 1014 1092
rect 1458 1088 1459 1092
rect 2061 1088 2062 1092
rect 2605 1088 2606 1092
rect 2717 1088 2718 1092
rect 3614 1088 3622 1091
rect 3890 1088 3891 1092
rect 4086 1088 4097 1091
rect 4578 1088 4579 1092
rect 4834 1088 4835 1092
rect 766 1078 774 1081
rect 782 1078 801 1081
rect 2541 1078 2542 1082
rect 2854 1078 2873 1081
rect 2882 1078 2890 1081
rect 766 1077 770 1078
rect 2886 1077 2890 1078
rect 3302 1074 3306 1078
rect 3382 1072 3385 1081
rect 3390 1078 3409 1081
rect 3626 1078 3633 1081
rect 4086 1081 4089 1088
rect 134 1062 137 1071
rect 1126 1068 1134 1071
rect 106 1058 113 1061
rect 230 1058 238 1061
rect 378 1058 385 1061
rect 538 1058 561 1061
rect 730 1058 737 1061
rect 1074 1058 1081 1061
rect 1094 1058 1113 1061
rect 1122 1058 1145 1061
rect 1182 1058 1190 1061
rect 1614 1062 1617 1071
rect 1854 1068 1862 1071
rect 2478 1068 2489 1071
rect 2634 1068 2641 1071
rect 2773 1068 2774 1072
rect 2834 1068 2841 1071
rect 3114 1068 3137 1071
rect 3226 1068 3233 1071
rect 3410 1068 3417 1071
rect 3630 1071 3633 1078
rect 3630 1068 3641 1071
rect 3718 1071 3721 1081
rect 4070 1078 4089 1081
rect 4366 1078 4378 1081
rect 4374 1077 4378 1078
rect 3702 1068 3721 1071
rect 4022 1068 4030 1071
rect 4062 1068 4070 1071
rect 1630 1058 1646 1061
rect 1814 1058 1830 1061
rect 1846 1058 1854 1061
rect 1926 1058 1953 1061
rect 2110 1058 2118 1061
rect 2282 1058 2289 1061
rect 2410 1058 2417 1061
rect 2434 1058 2449 1061
rect 2502 1058 2529 1061
rect 2558 1058 2566 1061
rect 2634 1058 2641 1061
rect 2682 1058 2689 1061
rect 2854 1058 2857 1068
rect 2918 1058 2926 1061
rect 3154 1058 3161 1061
rect 3442 1058 3449 1061
rect 3462 1058 3481 1061
rect 3546 1058 3553 1061
rect 3642 1058 3649 1061
rect 4222 1062 4225 1071
rect 4358 1068 4366 1071
rect 4614 1071 4617 1081
rect 4614 1068 4633 1071
rect 5046 1068 5049 1078
rect 3866 1058 3873 1061
rect 4026 1058 4041 1061
rect 4046 1058 4054 1061
rect 4146 1058 4153 1061
rect 4426 1058 4433 1061
rect 4522 1058 4529 1061
rect 4586 1058 4593 1061
rect 4986 1058 4993 1061
rect 5058 1058 5073 1061
rect 182 1048 185 1058
rect 546 1048 553 1051
rect 1026 1048 1033 1051
rect 1094 1048 1097 1058
rect 1158 1048 1161 1058
rect 1570 1048 1585 1051
rect 1594 1048 1598 1052
rect 1702 1051 1706 1054
rect 1670 1048 1689 1051
rect 1694 1048 1706 1051
rect 1810 1048 1814 1052
rect 1882 1048 1889 1051
rect 1894 1048 1905 1051
rect 2034 1048 2038 1052
rect 2106 1048 2110 1052
rect 2258 1048 2262 1052
rect 2450 1048 2454 1052
rect 2462 1048 2470 1051
rect 3254 1048 3273 1051
rect 3462 1048 3465 1058
rect 3650 1048 3654 1052
rect 3982 1048 4001 1051
rect 1902 1042 1905 1048
rect 197 1038 198 1042
rect 354 1038 355 1042
rect 386 1038 387 1042
rect 526 1038 554 1041
rect 1146 1038 1147 1042
rect 1181 1038 1182 1042
rect 3278 1041 3282 1044
rect 3470 1042 3474 1044
rect 3686 1042 3690 1044
rect 3278 1038 3289 1041
rect 3862 1042 3866 1044
rect 3974 1042 3978 1044
rect 536 1003 538 1007
rect 542 1003 545 1007
rect 549 1003 552 1007
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1573 1003 1576 1007
rect 2584 1003 2586 1007
rect 2590 1003 2593 1007
rect 2597 1003 2600 1007
rect 3608 1003 3610 1007
rect 3614 1003 3617 1007
rect 3621 1003 3624 1007
rect 4632 1003 4634 1007
rect 4638 1003 4641 1007
rect 4645 1003 4648 1007
rect 370 988 371 992
rect 1778 988 1779 992
rect 2030 988 2038 991
rect 2226 988 2227 992
rect 2941 988 2942 992
rect 2986 988 2987 992
rect 3397 988 3398 992
rect 3738 988 3739 992
rect 3818 988 3819 992
rect 3997 988 3998 992
rect 4413 988 4414 992
rect 1130 968 1131 972
rect 1358 968 1370 971
rect 1550 968 1558 971
rect 1854 968 1865 971
rect 2835 968 2838 972
rect 4098 968 4113 971
rect 210 958 214 962
rect 38 948 46 951
rect 222 951 225 961
rect 222 948 241 951
rect 382 951 385 961
rect 382 948 401 951
rect 494 948 502 951
rect 846 951 849 961
rect 830 948 849 951
rect 62 932 65 942
rect 694 941 697 948
rect 990 948 1006 951
rect 1054 948 1062 951
rect 1142 951 1145 961
rect 1494 958 1502 961
rect 1142 948 1161 951
rect 1254 948 1262 951
rect 1370 948 1377 951
rect 1486 948 1497 951
rect 1574 951 1577 961
rect 1586 958 1590 962
rect 1842 958 1846 962
rect 1542 948 1577 951
rect 1814 948 1822 951
rect 1990 951 1993 961
rect 2002 958 2006 962
rect 2162 958 2166 962
rect 1974 948 1993 951
rect 2006 948 2022 951
rect 2298 948 2305 951
rect 1494 942 1497 948
rect 686 938 697 941
rect 1414 938 1422 941
rect 2350 941 2353 948
rect 2910 948 2918 951
rect 3266 948 3273 951
rect 3286 951 3289 961
rect 3286 948 3305 951
rect 3358 948 3385 951
rect 3446 948 3462 951
rect 3486 951 3489 961
rect 3470 948 3489 951
rect 3730 948 3737 951
rect 3790 948 3798 951
rect 3998 948 4006 951
rect 2350 938 2362 941
rect 2526 938 2534 941
rect 2678 938 2686 941
rect 2690 938 2697 941
rect 2886 938 2905 941
rect 2478 928 2497 931
rect 2886 928 2889 938
rect 3094 932 3097 942
rect 3446 941 3449 948
rect 3334 938 3345 941
rect 3438 938 3449 941
rect 3758 938 3774 941
rect 4006 938 4014 941
rect 4214 941 4217 948
rect 4342 951 4345 961
rect 4754 958 4758 962
rect 4974 952 4977 961
rect 5158 958 5177 961
rect 4342 948 4361 951
rect 4462 948 4470 951
rect 4522 948 4537 951
rect 4726 948 4734 951
rect 4970 948 4974 951
rect 4206 938 4217 941
rect 4422 938 4449 941
rect 4770 938 4777 941
rect 4886 938 4889 948
rect 5150 948 5158 951
rect 5022 938 5030 941
rect 5134 938 5137 948
rect 3158 928 3161 938
rect 4018 928 4022 932
rect 4222 931 4226 933
rect 4046 928 4065 931
rect 4214 928 4226 931
rect 4942 928 4961 931
rect 5038 931 5042 933
rect 5030 928 5042 931
rect 517 918 518 922
rect 1434 918 1435 922
rect 3021 918 3022 922
rect 3126 918 3134 921
rect 5005 918 5006 922
rect 1048 903 1050 907
rect 1054 903 1057 907
rect 1061 903 1064 907
rect 2072 903 2074 907
rect 2078 903 2081 907
rect 2085 903 2088 907
rect 3096 903 3098 907
rect 3102 903 3105 907
rect 3109 903 3112 907
rect 4112 903 4114 907
rect 4118 903 4121 907
rect 4125 903 4128 907
rect 882 888 883 892
rect 973 888 974 892
rect 1634 888 1635 892
rect 1658 888 1659 892
rect 1810 888 1811 892
rect 3818 888 3819 892
rect 4242 888 4243 892
rect 4266 888 4267 892
rect 4546 888 4547 892
rect 4874 888 4875 892
rect 318 878 337 881
rect 554 878 561 881
rect 2270 878 2289 881
rect 2342 878 2361 881
rect 2654 878 2673 881
rect 3726 878 3745 881
rect 3950 878 3969 881
rect 4430 878 4449 881
rect 4578 878 4579 882
rect 3670 876 3674 878
rect 814 868 822 871
rect 938 868 945 871
rect 1034 868 1042 871
rect 1190 868 1198 871
rect 1293 868 1294 872
rect 1578 868 1593 871
rect 1922 868 1930 871
rect 2306 868 2329 871
rect 2790 868 2802 871
rect 2966 868 2977 871
rect 3254 868 3265 871
rect 3390 868 3401 871
rect 3410 868 3417 871
rect 3541 868 3542 872
rect 3690 868 3697 871
rect 3942 868 3950 871
rect 4062 868 4089 871
rect 4250 868 4257 871
rect 4530 868 4537 871
rect 4642 868 4657 871
rect 4734 871 4737 881
rect 5022 878 5034 881
rect 5030 877 5034 878
rect 4718 868 4737 871
rect 5014 868 5022 871
rect 5150 868 5158 871
rect 126 858 145 861
rect 198 858 206 861
rect 278 858 286 861
rect 318 858 321 868
rect 402 858 409 861
rect 622 858 641 861
rect 830 861 833 868
rect 830 858 849 861
rect 1158 858 1177 861
rect 1374 858 1393 861
rect 1558 858 1593 861
rect 1726 858 1745 861
rect 1978 858 1985 861
rect 2046 858 2065 861
rect 2186 858 2201 861
rect 2582 858 2617 861
rect 2850 858 2857 861
rect 2918 858 2937 861
rect 3142 858 3161 861
rect 3206 858 3225 861
rect 3350 858 3369 861
rect 3438 858 3457 861
rect 3862 858 3870 861
rect 4090 858 4097 861
rect 4102 858 4118 861
rect 4518 858 4526 861
rect 4678 858 4697 861
rect 4918 858 4934 861
rect 5082 858 5089 861
rect 126 848 129 858
rect 638 848 641 858
rect 986 848 993 851
rect 1158 848 1161 858
rect 1206 848 1225 851
rect 1374 848 1377 858
rect 1590 848 1593 858
rect 1726 848 1729 858
rect 1790 848 1798 851
rect 2046 848 2049 858
rect 2590 848 2598 851
rect 2614 848 2617 858
rect 2918 848 2921 858
rect 3130 848 3134 852
rect 3142 848 3145 858
rect 3206 848 3209 858
rect 3366 848 3369 858
rect 3438 848 3441 858
rect 4022 848 4041 851
rect 4246 848 4254 851
rect 4678 848 4681 858
rect 4994 848 4998 852
rect 3358 842 3362 844
rect 4550 842 4554 844
rect 254 838 266 841
rect 515 838 518 842
rect 862 838 870 841
rect 946 838 953 841
rect 2515 838 2518 842
rect 3426 838 3427 842
rect 277 818 278 822
rect 589 818 590 822
rect 850 818 851 822
rect 1714 818 1715 822
rect 3485 818 3486 822
rect 4053 818 4054 822
rect 4506 818 4507 822
rect 536 803 538 807
rect 542 803 545 807
rect 549 803 552 807
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1573 803 1576 807
rect 2584 803 2586 807
rect 2590 803 2593 807
rect 2597 803 2600 807
rect 3608 803 3610 807
rect 3614 803 3617 807
rect 3621 803 3624 807
rect 4632 803 4634 807
rect 4638 803 4641 807
rect 4645 803 4648 807
rect 181 788 182 792
rect 714 788 715 792
rect 989 788 990 792
rect 1082 788 1083 792
rect 1394 788 1395 792
rect 2285 788 2286 792
rect 2394 788 2395 792
rect 2418 788 2419 792
rect 2613 788 2614 792
rect 3266 788 3267 792
rect 3677 788 3678 792
rect 3786 788 3787 792
rect 3877 788 3878 792
rect 4034 788 4035 792
rect 4530 788 4531 792
rect 4589 788 4590 792
rect 242 768 243 772
rect 675 768 678 772
rect 1250 768 1251 772
rect 1510 768 1518 771
rect 1510 766 1514 768
rect 1550 766 1554 768
rect 2230 768 2238 771
rect 2365 768 2366 772
rect 4658 768 4661 772
rect 1614 766 1618 768
rect 4278 766 4282 768
rect 474 758 478 762
rect 258 748 265 751
rect 486 751 489 761
rect 486 748 505 751
rect 510 748 526 751
rect 574 751 577 761
rect 586 758 590 762
rect 974 752 977 761
rect 530 748 553 751
rect 558 748 577 751
rect 806 748 814 751
rect 1110 751 1113 761
rect 1282 758 1286 762
rect 1106 748 1113 751
rect 1174 748 1182 751
rect 1342 748 1350 751
rect 1358 748 1366 751
rect 1866 748 1881 751
rect 2082 748 2105 751
rect 2110 748 2118 751
rect 2242 748 2249 751
rect 2350 751 2353 761
rect 3018 758 3022 762
rect 2926 753 2930 758
rect 2334 748 2353 751
rect 2398 748 2406 751
rect 2442 748 2449 751
rect 2626 748 2633 751
rect 3030 751 3033 761
rect 3030 748 3049 751
rect 3122 748 3145 751
rect 3318 751 3321 761
rect 3302 748 3321 751
rect 3358 748 3385 751
rect 3398 751 3401 761
rect 3398 748 3417 751
rect 3658 748 3665 751
rect 3706 748 3713 751
rect 3862 751 3865 761
rect 3846 748 3865 751
rect 3954 748 3961 751
rect 3986 748 3993 751
rect 4046 748 4054 751
rect 4066 748 4073 751
rect 4078 748 4086 751
rect 4246 751 4249 761
rect 4246 748 4265 751
rect 4298 748 4305 751
rect 4318 748 4345 751
rect 4386 748 4393 751
rect 278 738 286 741
rect 522 738 545 741
rect 1322 738 1329 741
rect 1374 738 1385 741
rect 1486 738 1494 741
rect 1562 738 1577 741
rect 1594 738 1601 741
rect 1910 738 1922 741
rect 2294 738 2305 741
rect 2402 738 2409 741
rect 2574 738 2590 741
rect 2638 738 2657 741
rect 3062 738 3070 741
rect 3246 738 3257 741
rect 3886 738 3897 741
rect 3918 738 3926 741
rect 4086 738 4102 741
rect 4302 738 4305 748
rect 4542 748 4558 751
rect 4682 748 4697 751
rect 4866 748 4873 751
rect 4998 748 5006 751
rect 4766 738 4785 741
rect 126 728 145 731
rect 206 728 209 738
rect 950 732 953 738
rect 950 728 958 732
rect 2654 728 2657 738
rect 2910 731 2914 733
rect 2902 728 2914 731
rect 3902 728 3910 731
rect 4198 731 4202 733
rect 4198 728 4209 731
rect 4614 728 4633 731
rect 4750 728 4758 731
rect 4782 728 4785 738
rect 5038 732 5042 736
rect 4918 728 4937 731
rect 1458 718 1459 722
rect 1477 718 1478 722
rect 1506 718 1507 722
rect 3165 718 3166 722
rect 3357 718 3358 722
rect 4630 721 4633 728
rect 4630 718 4641 721
rect 5069 718 5070 722
rect 1048 703 1050 707
rect 1054 703 1057 707
rect 1061 703 1064 707
rect 2072 703 2074 707
rect 2078 703 2081 707
rect 2085 703 2088 707
rect 3096 703 3098 707
rect 3102 703 3105 707
rect 3109 703 3112 707
rect 4112 703 4114 707
rect 4118 703 4121 707
rect 4125 703 4128 707
rect 573 688 574 692
rect 901 688 902 692
rect 981 688 982 692
rect 1106 688 1113 691
rect 1149 688 1150 692
rect 1405 688 1406 692
rect 2333 688 2334 692
rect 4378 688 4379 692
rect 4626 688 4627 692
rect 4078 681 4081 688
rect 3910 678 3929 681
rect 4078 678 4098 681
rect 4262 678 4274 681
rect 5014 678 5033 681
rect 5086 678 5098 681
rect 1310 674 1314 678
rect 4094 677 4098 678
rect 4270 677 4274 678
rect 5094 677 5098 678
rect 3726 672 3730 674
rect 542 668 558 671
rect 230 658 249 661
rect 298 658 305 661
rect 374 658 382 661
rect 502 658 521 661
rect 534 658 566 661
rect 854 658 873 661
rect 878 658 886 661
rect 942 658 961 661
rect 1126 658 1134 661
rect 1158 661 1161 671
rect 1158 658 1166 661
rect 1358 658 1377 661
rect 1486 658 1494 661
rect 1638 658 1657 661
rect 1726 658 1745 661
rect 1826 658 1833 661
rect 2158 658 2166 661
rect 2294 662 2297 671
rect 2446 662 2449 671
rect 3038 668 3046 671
rect 3622 668 3650 671
rect 4598 668 4606 671
rect 4758 668 4766 671
rect 5042 668 5049 671
rect 2666 658 2673 661
rect 3038 658 3057 661
rect 3134 658 3153 661
rect 3494 658 3513 661
rect 3746 658 3753 661
rect 3766 658 3785 661
rect 3858 658 3865 661
rect 4126 658 4134 661
rect 4322 658 4329 661
rect 4538 658 4545 661
rect 4662 658 4681 661
rect 4946 658 4953 661
rect 230 648 233 658
rect 306 648 310 652
rect 518 648 521 658
rect 550 648 569 651
rect 854 648 857 658
rect 894 648 897 658
rect 942 648 945 658
rect 1358 648 1361 658
rect 1654 648 1657 658
rect 1742 648 1745 658
rect 1754 648 1758 652
rect 1946 648 1950 652
rect 2010 648 2014 652
rect 2022 648 2030 651
rect 2166 648 2174 651
rect 2286 651 2290 654
rect 2286 648 2297 651
rect 2466 648 2470 652
rect 2886 648 2889 658
rect 2894 648 2913 651
rect 2922 648 2926 652
rect 3038 648 3041 658
rect 3150 648 3153 658
rect 3494 648 3497 658
rect 3754 648 3758 652
rect 3766 648 3769 658
rect 4630 648 4646 651
rect 4678 648 4681 658
rect 550 642 553 648
rect 1398 642 1402 644
rect 2414 642 2418 644
rect 2990 642 2994 644
rect 373 638 374 642
rect 459 638 462 642
rect 1086 638 1114 641
rect 1610 638 1611 642
rect 2115 638 2118 642
rect 2782 638 2794 641
rect 3046 642 3050 644
rect 3278 642 3282 644
rect 3398 642 3402 644
rect 3554 638 3557 642
rect 2674 628 2675 632
rect 274 618 275 622
rect 536 603 538 607
rect 542 603 545 607
rect 549 603 552 607
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1573 603 1576 607
rect 2584 603 2586 607
rect 2590 603 2593 607
rect 2597 603 2600 607
rect 3608 603 3610 607
rect 3614 603 3617 607
rect 3621 603 3624 607
rect 4632 603 4634 607
rect 4638 603 4641 607
rect 4645 603 4648 607
rect 813 588 814 592
rect 845 588 846 592
rect 874 588 875 592
rect 1037 588 1038 592
rect 1194 588 1195 592
rect 3397 588 3398 592
rect 3866 588 3867 592
rect 4018 588 4019 592
rect 4149 588 4150 592
rect 4181 588 4182 592
rect 4413 588 4414 592
rect 1469 578 1470 582
rect 427 568 430 572
rect 925 568 926 572
rect 1803 568 1806 572
rect 1963 568 1966 572
rect 1982 568 1994 571
rect 2005 568 2006 572
rect 2078 568 2086 571
rect 3773 568 3774 572
rect 3834 568 3835 572
rect 4074 568 4075 572
rect 4086 568 4094 571
rect 114 558 118 562
rect 126 551 129 561
rect 126 548 145 551
rect 190 548 198 551
rect 222 551 225 561
rect 222 548 241 551
rect 246 548 254 551
rect 314 548 321 551
rect 598 551 601 561
rect 610 558 614 562
rect 766 558 774 561
rect 582 548 601 551
rect 814 548 830 551
rect 1006 548 1014 551
rect 1142 548 1150 551
rect 1326 551 1329 561
rect 1298 548 1305 551
rect 1310 548 1329 551
rect 1470 548 1478 551
rect 1590 548 1598 551
rect 1698 548 1713 551
rect 1862 551 1865 561
rect 1846 548 1865 551
rect 2006 548 2014 551
rect 2026 548 2033 551
rect 2102 551 2105 561
rect 2982 558 2990 561
rect 3330 558 3334 562
rect 3362 558 3366 562
rect 3546 558 3553 561
rect 2058 548 2065 551
rect 2070 548 2105 551
rect 2274 548 2289 551
rect 2314 548 2321 551
rect 2326 548 2334 551
rect 2390 548 2398 551
rect 2470 548 2478 551
rect 350 538 362 541
rect 506 538 507 542
rect 786 538 793 541
rect 1154 538 1161 541
rect 1218 538 1225 541
rect 1670 538 1673 548
rect 2750 542 2753 551
rect 2774 548 2782 551
rect 2814 548 2830 551
rect 3274 548 3281 551
rect 3366 548 3374 551
rect 3430 548 3438 551
rect 3774 548 3782 551
rect 3826 548 3833 551
rect 3962 548 3969 551
rect 4134 551 4137 561
rect 4450 558 4457 561
rect 4658 558 4662 562
rect 4058 548 4073 551
rect 4102 548 4137 551
rect 4322 548 4337 551
rect 2262 538 2270 541
rect 2790 538 2801 541
rect 3146 538 3153 541
rect 3158 538 3174 541
rect 3542 538 3550 541
rect 3610 538 3617 541
rect 3790 538 3793 548
rect 4446 541 4449 548
rect 4978 548 4993 551
rect 5118 548 5126 551
rect 4438 538 4449 541
rect 4462 538 4478 541
rect 5054 538 5073 541
rect 2734 528 2753 531
rect 2910 528 2929 531
rect 3126 528 3145 531
rect 4230 528 4249 531
rect 4462 528 4465 538
rect 4774 528 4793 531
rect 4830 528 4849 531
rect 4886 528 4905 531
rect 5054 528 5057 538
rect 4386 518 4387 522
rect 1048 503 1050 507
rect 1054 503 1057 507
rect 1061 503 1064 507
rect 2072 503 2074 507
rect 2078 503 2081 507
rect 2085 503 2088 507
rect 3096 503 3098 507
rect 3102 503 3105 507
rect 3109 503 3112 507
rect 4112 503 4114 507
rect 4118 503 4121 507
rect 4125 503 4128 507
rect 477 488 478 492
rect 645 488 646 492
rect 917 488 918 492
rect 1197 488 1198 492
rect 1453 488 1454 492
rect 2389 488 2390 492
rect 2501 488 2502 492
rect 2606 488 2622 491
rect 2821 488 2822 492
rect 3381 488 3382 492
rect 4098 488 4099 492
rect 4410 488 4411 492
rect 4490 488 4491 492
rect 4646 488 4662 491
rect 5106 488 5107 492
rect 286 478 297 481
rect 286 477 290 478
rect 130 468 137 471
rect 506 468 514 471
rect 854 468 865 471
rect 74 458 81 461
rect 162 458 177 461
rect 854 462 857 468
rect 342 458 350 461
rect 430 458 449 461
rect 630 458 638 461
rect 714 458 721 461
rect 842 458 854 461
rect 934 461 937 481
rect 3350 478 3358 481
rect 1630 474 1634 478
rect 3350 477 3354 478
rect 930 458 937 461
rect 974 458 993 461
rect 1502 462 1505 471
rect 1486 458 1494 461
rect 1806 458 1822 461
rect 1838 458 1857 461
rect 1870 458 1878 461
rect 1938 458 1945 461
rect 2030 458 2049 461
rect 2430 461 2433 471
rect 2486 468 2497 471
rect 3070 468 3086 471
rect 3478 471 3481 481
rect 3942 478 3961 481
rect 4198 474 4202 478
rect 3462 468 3481 471
rect 3962 468 3969 471
rect 4246 471 4249 481
rect 4446 478 4465 481
rect 4526 478 4545 481
rect 4658 478 4673 481
rect 4678 478 4697 481
rect 5046 478 5065 481
rect 4878 472 4881 478
rect 4230 468 4249 471
rect 4374 468 4385 471
rect 4438 468 4446 471
rect 4878 468 4882 472
rect 2494 462 2497 468
rect 2426 458 2433 461
rect 2626 458 2641 461
rect 2842 458 2849 461
rect 3118 458 3137 461
rect 3662 458 3670 461
rect 3822 458 3830 461
rect 4374 462 4377 468
rect 4042 458 4049 461
rect 4590 458 4598 461
rect 4802 458 4809 461
rect 5062 458 5065 468
rect 430 448 433 458
rect 618 448 622 452
rect 630 448 633 458
rect 770 448 774 452
rect 802 448 806 452
rect 974 448 977 458
rect 1058 448 1065 451
rect 1482 448 1486 452
rect 1722 448 1726 452
rect 1854 448 1857 458
rect 2046 448 2049 458
rect 2350 448 2353 458
rect 2814 448 2817 458
rect 3134 448 3137 458
rect 3422 448 3441 451
rect 3678 451 3682 454
rect 3670 448 3682 451
rect 1022 442 1026 444
rect 178 438 179 442
rect 267 438 270 442
rect 1190 441 1194 444
rect 2998 442 3002 444
rect 1182 438 1194 441
rect 2606 438 2634 441
rect 3374 442 3378 444
rect 53 418 54 422
rect 1226 418 1227 422
rect 2978 418 2979 422
rect 536 403 538 407
rect 542 403 545 407
rect 549 403 552 407
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1573 403 1576 407
rect 2584 403 2586 407
rect 2590 403 2593 407
rect 2597 403 2600 407
rect 3608 403 3610 407
rect 3614 403 3617 407
rect 3621 403 3624 407
rect 4632 403 4634 407
rect 4638 403 4641 407
rect 4645 403 4648 407
rect 634 388 635 392
rect 1046 388 1062 391
rect 1082 388 1083 392
rect 1421 388 1422 392
rect 1693 388 1694 392
rect 1914 388 1915 392
rect 2362 388 2363 392
rect 2666 388 2667 392
rect 3578 388 3579 392
rect 3642 388 3643 392
rect 3866 388 3867 392
rect 4818 388 4819 392
rect 346 378 347 382
rect 486 368 502 371
rect 1011 368 1014 372
rect 1114 368 1115 372
rect 1453 368 1454 372
rect 1546 368 1547 372
rect 1558 368 1566 371
rect 1782 368 1793 371
rect 2093 368 2094 372
rect 2259 368 2262 372
rect 2330 368 2331 372
rect 2406 368 2417 371
rect 2915 368 2918 372
rect 3501 368 3502 372
rect 3834 368 3835 372
rect 4178 368 4186 371
rect 4434 368 4437 372
rect 4930 368 4933 372
rect 2414 362 2417 368
rect 38 348 54 351
rect 206 351 209 361
rect 378 358 382 362
rect 474 358 478 362
rect 822 358 830 361
rect 190 348 209 351
rect 270 348 278 351
rect 394 348 409 351
rect 422 348 441 351
rect 446 348 454 351
rect 422 342 425 348
rect 626 348 633 351
rect 894 351 897 361
rect 1770 358 1774 362
rect 878 348 897 351
rect 1234 348 1241 351
rect 1506 348 1513 351
rect 1842 348 1849 351
rect 1966 348 1974 351
rect 2078 351 2081 361
rect 2046 348 2081 351
rect 2158 351 2161 361
rect 2394 358 2398 362
rect 2698 358 2702 362
rect 2142 348 2161 351
rect 1486 338 1494 341
rect 1750 338 1753 348
rect 2310 348 2318 351
rect 2346 348 2361 351
rect 2378 348 2393 351
rect 1894 338 1905 341
rect 2310 338 2313 348
rect 2658 348 2665 351
rect 2710 351 2713 361
rect 2810 358 2814 362
rect 2822 358 2830 361
rect 2710 348 2729 351
rect 2962 348 2969 351
rect 3022 351 3025 361
rect 3290 358 3294 362
rect 3006 348 3025 351
rect 3302 351 3305 361
rect 4194 358 4198 362
rect 4522 358 4526 362
rect 3302 348 3321 351
rect 3390 348 3398 351
rect 3458 348 3465 351
rect 3534 348 3542 351
rect 3678 348 3686 351
rect 3738 348 3753 351
rect 3882 348 3889 351
rect 2646 338 2657 341
rect 3050 338 3062 341
rect 1014 332 1018 336
rect 1382 331 1386 333
rect 3126 332 3129 342
rect 3542 338 3550 341
rect 3558 338 3569 341
rect 3814 338 3817 348
rect 3914 338 3929 341
rect 4062 341 4065 348
rect 4210 348 4225 351
rect 4230 348 4238 351
rect 4290 348 4305 351
rect 4390 348 4398 351
rect 4538 348 4553 351
rect 4698 348 4705 351
rect 4054 338 4065 341
rect 4366 338 4385 341
rect 5030 338 5049 341
rect 1382 328 1393 331
rect 4366 328 4369 338
rect 4394 328 4401 331
rect 4582 328 4601 331
rect 4758 328 4761 338
rect 5030 328 5033 338
rect 5086 328 5105 331
rect 4882 318 4883 322
rect 1048 303 1050 307
rect 1054 303 1057 307
rect 1061 303 1064 307
rect 2072 303 2074 307
rect 2078 303 2081 307
rect 2085 303 2088 307
rect 3096 303 3098 307
rect 3102 303 3105 307
rect 3109 303 3112 307
rect 4112 303 4114 307
rect 4118 303 4121 307
rect 4125 303 4128 307
rect 1069 288 1070 292
rect 1517 288 1518 292
rect 1550 288 1566 291
rect 1917 288 1918 292
rect 3437 288 3438 292
rect 1398 274 1402 278
rect 3334 278 3353 281
rect 4038 278 4057 281
rect 4062 278 4074 281
rect 1710 274 1714 278
rect 4070 277 4074 278
rect 126 258 145 261
rect 614 262 617 271
rect 1038 268 1062 271
rect 1302 268 1313 271
rect 1554 268 1577 271
rect 358 258 374 261
rect 570 258 593 261
rect 674 258 681 261
rect 750 258 769 261
rect 1302 262 1305 268
rect 1006 258 1025 261
rect 1354 258 1361 261
rect 1366 258 1374 261
rect 1598 262 1601 271
rect 2110 268 2138 271
rect 2542 268 2550 271
rect 2554 268 2570 271
rect 2750 268 2758 271
rect 2906 268 2913 271
rect 2966 268 2974 271
rect 1610 258 1617 261
rect 1690 258 1697 261
rect 1766 258 1785 261
rect 1982 258 2001 261
rect 2006 258 2014 261
rect 2254 258 2273 261
rect 2278 258 2286 261
rect 2406 258 2425 261
rect 2618 258 2625 261
rect 2678 258 2686 261
rect 2698 258 2705 261
rect 2750 258 2769 261
rect 2906 258 2921 261
rect 2934 258 2942 261
rect 2990 258 2998 261
rect 3166 258 3185 261
rect 3246 258 3254 261
rect 3266 258 3273 261
rect 3370 258 3377 261
rect 3390 258 3409 261
rect 3566 258 3590 261
rect 3694 262 3697 271
rect 3730 258 3737 261
rect 3754 258 3769 261
rect 3774 258 3782 261
rect 3842 258 3849 261
rect 4202 258 4217 261
rect 4390 261 4393 271
rect 4550 268 4562 271
rect 4694 271 4697 281
rect 4810 278 4818 281
rect 4814 277 4818 278
rect 4666 268 4681 271
rect 4694 268 4713 271
rect 4998 268 5010 271
rect 4390 258 4398 261
rect 4414 258 4433 261
rect 4742 258 4761 261
rect 114 248 118 252
rect 126 248 129 258
rect 422 248 425 258
rect 606 248 609 258
rect 666 248 673 251
rect 750 248 753 258
rect 1006 248 1009 258
rect 1282 248 1286 252
rect 1618 248 1622 252
rect 1782 248 1785 258
rect 1794 248 1798 252
rect 1982 248 1985 258
rect 2254 248 2257 258
rect 2422 248 2425 258
rect 2434 248 2438 252
rect 2654 251 2658 254
rect 2654 248 2665 251
rect 2674 248 2678 252
rect 2750 248 2753 258
rect 2934 248 2937 258
rect 3018 248 3022 252
rect 3182 248 3185 258
rect 3390 248 3393 258
rect 3598 251 3602 254
rect 3574 248 3602 251
rect 4218 248 4222 252
rect 4430 248 4433 258
rect 4758 248 4761 258
rect 2758 242 2762 244
rect 414 238 426 241
rect 1082 238 1090 241
rect 1374 238 1385 241
rect 2363 238 2366 242
rect 2851 238 2854 242
rect 3474 238 3477 242
rect 3738 238 3739 242
rect 4834 238 4837 242
rect 181 218 182 222
rect 309 218 310 222
rect 738 218 739 222
rect 2957 218 2958 222
rect 3197 218 3198 222
rect 3378 218 3379 222
rect 4445 218 4446 222
rect 4773 218 4774 222
rect 536 203 538 207
rect 542 203 545 207
rect 549 203 552 207
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1573 203 1576 207
rect 2584 203 2586 207
rect 2590 203 2593 207
rect 2597 203 2600 207
rect 3608 203 3610 207
rect 3614 203 3617 207
rect 3621 203 3624 207
rect 4632 203 4634 207
rect 4638 203 4641 207
rect 4645 203 4648 207
rect 781 188 782 192
rect 1834 188 1835 192
rect 2102 188 2118 191
rect 3226 188 3227 192
rect 4213 188 4214 192
rect 2701 178 2702 182
rect 1171 168 1174 172
rect 1683 168 1686 172
rect 2330 168 2331 172
rect 2813 168 2814 172
rect 3493 168 3494 172
rect 4254 168 4265 171
rect 202 148 209 151
rect 282 148 297 151
rect 454 151 457 161
rect 454 148 473 151
rect 706 148 713 151
rect 718 148 742 151
rect 766 151 769 161
rect 750 148 769 151
rect 782 148 798 151
rect 802 148 809 151
rect 846 148 854 151
rect 1074 148 1081 151
rect 1086 148 1094 151
rect 1230 151 1233 161
rect 1214 148 1233 151
rect 1246 148 1270 151
rect 1286 151 1289 161
rect 1286 148 1305 151
rect 1350 151 1353 161
rect 1350 148 1369 151
rect 1438 151 1441 161
rect 1722 158 1726 162
rect 1754 158 1758 162
rect 1422 148 1441 151
rect 1826 148 1833 151
rect 1878 151 1881 161
rect 2138 158 2142 162
rect 2158 152 2161 161
rect 1878 148 1897 151
rect 2270 148 2278 151
rect 2302 148 2310 151
rect 62 132 65 142
rect 726 138 734 141
rect 1066 138 1073 141
rect 1598 138 1606 141
rect 1814 138 1825 141
rect 2006 138 2018 141
rect 2222 138 2225 148
rect 2590 148 2598 151
rect 2658 148 2665 151
rect 2670 148 2678 151
rect 2702 148 2710 151
rect 2758 151 2761 161
rect 2906 158 2910 162
rect 2758 148 2777 151
rect 2878 148 2894 151
rect 2898 148 2905 151
rect 2970 148 2985 151
rect 3086 148 3094 151
rect 3390 151 3393 161
rect 3462 158 3481 161
rect 3390 148 3409 151
rect 3646 151 3649 161
rect 3846 158 3858 161
rect 3854 156 3858 158
rect 3594 148 3625 151
rect 3630 148 3649 151
rect 3730 148 3737 151
rect 3838 148 3846 151
rect 4086 151 4089 161
rect 4086 148 4105 151
rect 4198 151 4201 161
rect 4254 152 4257 161
rect 4746 158 4750 162
rect 4182 148 4201 151
rect 4450 148 4465 151
rect 4602 148 4609 151
rect 4670 148 4678 151
rect 4758 151 4761 161
rect 4758 148 4777 151
rect 4802 148 4809 151
rect 4878 151 4881 161
rect 4890 158 4894 162
rect 4862 148 4881 151
rect 5058 148 5065 151
rect 2534 138 2562 141
rect 2890 138 2897 141
rect 3358 138 3369 141
rect 3502 138 3513 141
rect 3602 138 3617 141
rect 3942 138 3950 141
rect 4158 138 4166 141
rect 254 128 273 131
rect 3342 131 3346 133
rect 3342 128 3353 131
rect 4638 131 4642 133
rect 4614 128 4642 131
rect 1048 103 1050 107
rect 1054 103 1057 107
rect 1061 103 1064 107
rect 2072 103 2074 107
rect 2078 103 2081 107
rect 2085 103 2088 107
rect 3096 103 3098 107
rect 3102 103 3105 107
rect 3109 103 3112 107
rect 4112 103 4114 107
rect 4118 103 4121 107
rect 4125 103 4128 107
rect 1062 88 1070 91
rect 1334 78 1353 81
rect 1558 78 1593 81
rect 2766 78 2785 81
rect 70 68 78 71
rect 502 68 505 78
rect 1074 68 1097 71
rect 2022 68 2033 71
rect 2634 68 2649 71
rect 350 58 358 61
rect 590 58 598 61
rect 774 58 793 61
rect 926 58 934 61
rect 1558 58 1566 61
rect 2022 62 2025 68
rect 2662 58 2686 61
rect 3054 62 3057 71
rect 3222 71 3225 81
rect 4278 78 4294 81
rect 4278 74 4282 78
rect 3222 68 3241 71
rect 3342 68 3354 71
rect 3782 68 3790 71
rect 2926 58 2942 61
rect 3222 58 3230 61
rect 3990 62 3993 71
rect 3506 58 3521 61
rect 3678 58 3697 61
rect 3894 58 3902 61
rect 4018 58 4030 61
rect 4222 62 4225 71
rect 5110 68 5118 71
rect 774 48 777 58
rect 954 48 958 52
rect 1798 48 1801 58
rect 3034 48 3038 52
rect 3678 48 3681 58
rect 4066 48 4070 52
rect 4078 48 4094 51
rect 4242 48 4246 52
rect 4370 48 4374 52
rect 4402 48 4406 52
rect 2690 38 2691 42
rect 4254 38 4265 41
rect 2078 18 2094 21
rect 536 3 538 7
rect 542 3 545 7
rect 549 3 552 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1573 3 1576 7
rect 2584 3 2586 7
rect 2590 3 2593 7
rect 2597 3 2600 7
rect 3608 3 3610 7
rect 3614 3 3617 7
rect 3621 3 3624 7
rect 4632 3 4634 7
rect 4638 3 4641 7
rect 4645 3 4648 7
<< m2contact >>
rect 1050 4903 1054 4907
rect 1057 4903 1061 4907
rect 2074 4903 2078 4907
rect 2081 4903 2085 4907
rect 3098 4903 3102 4907
rect 3105 4903 3109 4907
rect 4114 4903 4118 4907
rect 4121 4903 4125 4907
rect 974 4888 978 4892
rect 2302 4888 2306 4892
rect 2414 4888 2418 4892
rect 3614 4888 3618 4892
rect 3982 4888 3986 4892
rect 4998 4888 5002 4892
rect 830 4878 834 4882
rect 846 4878 850 4882
rect 878 4878 882 4882
rect 1254 4878 1258 4882
rect 78 4868 82 4872
rect 230 4868 234 4872
rect 270 4868 274 4872
rect 286 4868 290 4872
rect 374 4868 378 4872
rect 454 4868 458 4872
rect 582 4868 586 4872
rect 598 4868 602 4872
rect 142 4858 146 4862
rect 182 4858 186 4862
rect 214 4859 218 4863
rect 246 4858 250 4862
rect 262 4858 266 4862
rect 318 4858 322 4862
rect 478 4858 482 4862
rect 574 4858 578 4862
rect 614 4859 618 4863
rect 718 4868 722 4872
rect 862 4868 866 4872
rect 878 4868 882 4872
rect 894 4868 898 4872
rect 982 4868 986 4872
rect 1070 4868 1074 4872
rect 1150 4868 1154 4872
rect 1246 4868 1250 4872
rect 1270 4878 1274 4882
rect 1830 4878 1834 4882
rect 2270 4878 2274 4882
rect 3830 4878 3834 4882
rect 3862 4878 3866 4882
rect 4078 4878 4082 4882
rect 4222 4878 4226 4882
rect 1502 4868 1506 4872
rect 1518 4868 1522 4872
rect 1558 4868 1562 4872
rect 1662 4868 1666 4872
rect 1678 4868 1682 4872
rect 1774 4868 1778 4872
rect 638 4858 642 4862
rect 686 4858 690 4862
rect 694 4858 698 4862
rect 710 4858 714 4862
rect 766 4858 770 4862
rect 790 4858 794 4862
rect 830 4858 834 4862
rect 854 4858 858 4862
rect 910 4859 914 4863
rect 1046 4858 1050 4862
rect 1190 4858 1194 4862
rect 1238 4858 1242 4862
rect 1286 4858 1290 4862
rect 1294 4858 1298 4862
rect 1350 4859 1354 4863
rect 1374 4858 1378 4862
rect 1486 4859 1490 4863
rect 1526 4858 1530 4862
rect 1542 4858 1546 4862
rect 1598 4858 1602 4862
rect 1622 4858 1626 4862
rect 1670 4858 1674 4862
rect 1758 4859 1762 4863
rect 1814 4868 1818 4872
rect 1886 4868 1890 4872
rect 1974 4868 1978 4872
rect 2078 4868 2082 4872
rect 2134 4868 2138 4872
rect 2150 4868 2154 4872
rect 2262 4868 2266 4872
rect 2294 4868 2298 4872
rect 2382 4868 2386 4872
rect 2422 4868 2426 4872
rect 2462 4868 2466 4872
rect 2598 4868 2602 4872
rect 2694 4868 2698 4872
rect 2726 4868 2730 4872
rect 2814 4868 2818 4872
rect 2894 4868 2898 4872
rect 2982 4868 2986 4872
rect 3070 4868 3074 4872
rect 3126 4868 3130 4872
rect 3214 4868 3218 4872
rect 3254 4868 3258 4872
rect 3342 4868 3346 4872
rect 3382 4868 3386 4872
rect 3398 4868 3402 4872
rect 3870 4868 3874 4872
rect 3910 4868 3914 4872
rect 4062 4868 4066 4872
rect 5166 4878 5170 4882
rect 4238 4868 4242 4872
rect 4246 4868 4250 4872
rect 4358 4868 4362 4872
rect 4502 4868 4506 4872
rect 4702 4868 4706 4872
rect 4918 4868 4922 4872
rect 5030 4868 5034 4872
rect 1790 4858 1794 4862
rect 1814 4858 1818 4862
rect 1998 4858 2002 4862
rect 2086 4858 2090 4862
rect 2094 4858 2098 4862
rect 2126 4858 2130 4862
rect 2174 4858 2178 4862
rect 2254 4858 2258 4862
rect 2294 4858 2298 4862
rect 2366 4859 2370 4863
rect 2398 4858 2402 4862
rect 2422 4858 2426 4862
rect 2446 4858 2450 4862
rect 2478 4859 2482 4863
rect 2510 4858 2514 4862
rect 2550 4858 2554 4862
rect 2694 4858 2698 4862
rect 2702 4858 2706 4862
rect 2726 4858 2730 4862
rect 2790 4858 2794 4862
rect 2830 4858 2834 4862
rect 2966 4858 2970 4862
rect 3006 4858 3010 4862
rect 3070 4858 3074 4862
rect 3094 4858 3098 4862
rect 3150 4858 3154 4862
rect 3222 4858 3226 4862
rect 3278 4858 3282 4862
rect 3350 4858 3354 4862
rect 3366 4858 3370 4862
rect 3374 4858 3378 4862
rect 3406 4858 3410 4862
rect 3486 4858 3490 4862
rect 3558 4858 3562 4862
rect 3582 4858 3586 4862
rect 3670 4858 3674 4862
rect 3694 4858 3698 4862
rect 3766 4858 3770 4862
rect 3782 4858 3786 4862
rect 3846 4858 3850 4862
rect 3878 4858 3882 4862
rect 3918 4858 3922 4862
rect 4046 4859 4050 4863
rect 4142 4858 4146 4862
rect 4166 4858 4170 4862
rect 4206 4858 4210 4862
rect 4254 4858 4258 4862
rect 4286 4859 4290 4863
rect 4318 4858 4322 4862
rect 4574 4858 4578 4862
rect 4598 4858 4602 4862
rect 4686 4859 4690 4863
rect 4750 4858 4754 4862
rect 4774 4858 4778 4862
rect 4846 4858 4850 4862
rect 4870 4858 4874 4862
rect 4934 4859 4938 4863
rect 5022 4858 5026 4862
rect 5070 4858 5074 4862
rect 5102 4859 5106 4863
rect 5134 4858 5138 4862
rect 246 4848 250 4852
rect 558 4848 562 4852
rect 574 4848 578 4852
rect 710 4848 714 4852
rect 1542 4848 1546 4852
rect 1686 4848 1690 4852
rect 1790 4848 1794 4852
rect 2270 4848 2274 4852
rect 2446 4848 2450 4852
rect 2686 4848 2690 4852
rect 2702 4848 2706 4852
rect 3094 4848 3098 4852
rect 3238 4848 3242 4852
rect 3366 4848 3370 4852
rect 5006 4848 5010 4852
rect 958 4838 962 4842
rect 1214 4838 1218 4842
rect 1230 4838 1234 4842
rect 1710 4838 1714 4842
rect 2054 4838 2058 4842
rect 2110 4838 2114 4842
rect 2254 4838 2258 4842
rect 2670 4838 2674 4842
rect 3046 4838 3050 4842
rect 3190 4838 3194 4842
rect 3222 4838 3226 4842
rect 3318 4838 3322 4842
rect 5150 4838 5154 4842
rect 2734 4828 2738 4832
rect 14 4818 18 4822
rect 150 4818 154 4822
rect 366 4818 370 4822
rect 430 4818 434 4822
rect 534 4818 538 4822
rect 678 4818 682 4822
rect 1126 4818 1130 4822
rect 1310 4818 1314 4822
rect 1414 4818 1418 4822
rect 1422 4818 1426 4822
rect 1654 4818 1658 4822
rect 1694 4818 1698 4822
rect 1950 4818 1954 4822
rect 2230 4818 2234 4822
rect 2542 4818 2546 4822
rect 2566 4818 2570 4822
rect 2654 4818 2658 4822
rect 2838 4818 2842 4822
rect 3062 4818 3066 4822
rect 3206 4818 3210 4822
rect 3334 4818 3338 4822
rect 3430 4818 3434 4822
rect 3726 4818 3730 4822
rect 3822 4818 3826 4822
rect 3974 4818 3978 4822
rect 4094 4818 4098 4822
rect 4198 4818 4202 4822
rect 4350 4818 4354 4822
rect 4414 4818 4418 4822
rect 4438 4818 4442 4822
rect 4558 4818 4562 4822
rect 4622 4818 4626 4822
rect 4806 4818 4810 4822
rect 4902 4818 4906 4822
rect 5022 4818 5026 4822
rect 5038 4818 5042 4822
rect 5158 4818 5162 4822
rect 538 4803 542 4807
rect 545 4803 549 4807
rect 1562 4803 1566 4807
rect 1569 4803 1573 4807
rect 2586 4803 2590 4807
rect 2593 4803 2597 4807
rect 3610 4803 3614 4807
rect 3617 4803 3621 4807
rect 4634 4803 4638 4807
rect 4641 4803 4645 4807
rect 190 4788 194 4792
rect 318 4788 322 4792
rect 478 4788 482 4792
rect 558 4788 562 4792
rect 718 4788 722 4792
rect 1334 4788 1338 4792
rect 1686 4788 1690 4792
rect 1734 4788 1738 4792
rect 2502 4788 2506 4792
rect 3398 4788 3402 4792
rect 3462 4788 3466 4792
rect 4678 4788 4682 4792
rect 670 4778 674 4782
rect 4102 4778 4106 4782
rect 4198 4778 4202 4782
rect 94 4768 98 4772
rect 134 4768 138 4772
rect 206 4768 210 4772
rect 342 4768 346 4772
rect 502 4768 506 4772
rect 574 4768 578 4772
rect 726 4768 730 4772
rect 822 4768 826 4772
rect 918 4768 922 4772
rect 1014 4768 1018 4772
rect 1550 4768 1554 4772
rect 1606 4768 1610 4772
rect 1670 4768 1674 4772
rect 1750 4768 1754 4772
rect 2150 4768 2154 4772
rect 2198 4768 2202 4772
rect 2326 4768 2330 4772
rect 2358 4768 2362 4772
rect 2486 4768 2490 4772
rect 2518 4768 2522 4772
rect 2718 4768 2722 4772
rect 2758 4768 2762 4772
rect 3430 4768 3434 4772
rect 3806 4768 3810 4772
rect 3894 4768 3898 4772
rect 3910 4768 3914 4772
rect 4622 4768 4626 4772
rect 4694 4768 4698 4772
rect 38 4748 42 4752
rect 110 4748 114 4752
rect 118 4748 122 4752
rect 150 4748 154 4752
rect 190 4748 194 4752
rect 246 4748 250 4752
rect 318 4748 322 4752
rect 358 4748 362 4752
rect 398 4747 402 4751
rect 422 4748 426 4752
rect 478 4748 482 4752
rect 686 4758 690 4762
rect 702 4758 706 4762
rect 710 4758 714 4762
rect 726 4758 730 4762
rect 734 4758 738 4762
rect 790 4758 794 4762
rect 806 4758 810 4762
rect 1190 4758 1194 4762
rect 1574 4758 1578 4762
rect 1622 4758 1626 4762
rect 1638 4758 1642 4762
rect 1702 4758 1706 4762
rect 2182 4758 2186 4762
rect 2206 4758 2210 4762
rect 2222 4758 2226 4762
rect 558 4748 562 4752
rect 614 4748 618 4752
rect 638 4748 642 4752
rect 686 4748 690 4752
rect 750 4748 754 4752
rect 774 4748 778 4752
rect 790 4748 794 4752
rect 806 4748 810 4752
rect 854 4747 858 4751
rect 878 4748 882 4752
rect 966 4748 970 4752
rect 1070 4748 1074 4752
rect 1150 4748 1154 4752
rect 1182 4748 1186 4752
rect 1246 4748 1250 4752
rect 1310 4748 1314 4752
rect 1358 4748 1362 4752
rect 1398 4748 1402 4752
rect 1494 4748 1498 4752
rect 1518 4748 1522 4752
rect 1566 4748 1570 4752
rect 1590 4748 1594 4752
rect 1622 4748 1626 4752
rect 1638 4748 1642 4752
rect 1670 4748 1674 4752
rect 1702 4748 1706 4752
rect 1734 4748 1738 4752
rect 1790 4748 1794 4752
rect 1806 4748 1810 4752
rect 1854 4748 1858 4752
rect 1886 4748 1890 4752
rect 1942 4748 1946 4752
rect 1958 4748 1962 4752
rect 2006 4748 2010 4752
rect 2038 4748 2042 4752
rect 2054 4748 2058 4752
rect 2102 4747 2106 4751
rect 2182 4748 2186 4752
rect 2222 4748 2226 4752
rect 2278 4748 2282 4752
rect 2342 4748 2346 4752
rect 2374 4748 2378 4752
rect 2382 4748 2386 4752
rect 2430 4748 2434 4752
rect 2454 4748 2458 4752
rect 2502 4748 2506 4752
rect 2542 4748 2546 4752
rect 2558 4748 2562 4752
rect 2582 4748 2586 4752
rect 2622 4747 2626 4751
rect 2654 4748 2658 4752
rect 2702 4748 2706 4752
rect 2742 4758 2746 4762
rect 3382 4758 3386 4762
rect 3414 4758 3418 4762
rect 3446 4758 3450 4762
rect 3582 4758 3586 4762
rect 2742 4748 2746 4752
rect 2814 4748 2818 4752
rect 2902 4748 2906 4752
rect 2998 4748 3002 4752
rect 3110 4748 3114 4752
rect 3142 4747 3146 4751
rect 3174 4748 3178 4752
rect 3222 4748 3226 4752
rect 3230 4748 3234 4752
rect 3262 4748 3266 4752
rect 3318 4748 3322 4752
rect 3342 4748 3346 4752
rect 3398 4748 3402 4752
rect 3430 4748 3434 4752
rect 3462 4748 3466 4752
rect 3510 4748 3514 4752
rect 3582 4748 3586 4752
rect 3622 4758 3626 4762
rect 3854 4758 3858 4762
rect 3638 4748 3642 4752
rect 3710 4748 3714 4752
rect 3766 4748 3770 4752
rect 3798 4748 3802 4752
rect 3838 4748 3842 4752
rect 4086 4758 4090 4762
rect 4158 4758 4162 4762
rect 3870 4748 3874 4752
rect 3878 4748 3882 4752
rect 3950 4748 3954 4752
rect 4038 4748 4042 4752
rect 4102 4748 4106 4752
rect 4142 4748 4146 4752
rect 4542 4758 4546 4762
rect 4662 4758 4666 4762
rect 4990 4758 4994 4762
rect 4182 4748 4186 4752
rect 4246 4748 4250 4752
rect 4318 4748 4322 4752
rect 4390 4747 4394 4751
rect 4470 4748 4474 4752
rect 4526 4748 4530 4752
rect 4574 4747 4578 4751
rect 4678 4748 4682 4752
rect 4750 4748 4754 4752
rect 4766 4748 4770 4752
rect 4830 4748 4834 4752
rect 4846 4748 4850 4752
rect 4862 4748 4866 4752
rect 4902 4748 4906 4752
rect 4926 4748 4930 4752
rect 4974 4748 4978 4752
rect 4990 4748 4994 4752
rect 5030 4748 5034 4752
rect 5046 4748 5050 4752
rect 5126 4748 5130 4752
rect 5142 4748 5146 4752
rect 14 4738 18 4742
rect 102 4738 106 4742
rect 158 4738 162 4742
rect 182 4738 186 4742
rect 222 4738 226 4742
rect 310 4738 314 4742
rect 366 4738 370 4742
rect 470 4738 474 4742
rect 526 4738 530 4742
rect 550 4738 554 4742
rect 678 4738 682 4742
rect 726 4738 730 4742
rect 758 4738 762 4742
rect 766 4738 770 4742
rect 798 4738 802 4742
rect 958 4738 962 4742
rect 1046 4738 1050 4742
rect 1182 4738 1186 4742
rect 1206 4738 1210 4742
rect 1222 4738 1226 4742
rect 1350 4738 1354 4742
rect 1374 4738 1378 4742
rect 1598 4738 1602 4742
rect 1630 4738 1634 4742
rect 1662 4738 1666 4742
rect 1694 4738 1698 4742
rect 1718 4738 1722 4742
rect 1726 4738 1730 4742
rect 1862 4738 1866 4742
rect 1918 4738 1922 4742
rect 2022 4738 2026 4742
rect 2046 4738 2050 4742
rect 2086 4738 2090 4742
rect 2174 4738 2178 4742
rect 2230 4738 2234 4742
rect 2246 4738 2250 4742
rect 2334 4738 2338 4742
rect 2390 4738 2394 4742
rect 2494 4738 2498 4742
rect 2526 4738 2530 4742
rect 2566 4738 2570 4742
rect 2694 4738 2698 4742
rect 2750 4738 2754 4742
rect 2838 4738 2842 4742
rect 2878 4738 2882 4742
rect 2974 4738 2978 4742
rect 3158 4738 3162 4742
rect 3190 4738 3194 4742
rect 3214 4738 3218 4742
rect 3238 4738 3242 4742
rect 3254 4738 3258 4742
rect 3366 4738 3370 4742
rect 3406 4738 3410 4742
rect 3438 4738 3442 4742
rect 3470 4738 3474 4742
rect 3486 4738 3490 4742
rect 3574 4738 3578 4742
rect 3646 4738 3650 4742
rect 3734 4738 3738 4742
rect 3774 4738 3778 4742
rect 3790 4738 3794 4742
rect 3822 4738 3826 4742
rect 3830 4738 3834 4742
rect 3886 4738 3890 4742
rect 3974 4738 3978 4742
rect 4070 4738 4074 4742
rect 4110 4738 4114 4742
rect 4134 4738 4138 4742
rect 4166 4738 4170 4742
rect 4190 4738 4194 4742
rect 4278 4738 4282 4742
rect 4358 4738 4362 4742
rect 4406 4738 4410 4742
rect 4446 4738 4450 4742
rect 4518 4738 4522 4742
rect 4542 4738 4546 4742
rect 4558 4738 4562 4742
rect 4686 4738 4690 4742
rect 4710 4738 4714 4742
rect 4854 4738 4858 4742
rect 4950 4738 4954 4742
rect 4966 4738 4970 4742
rect 5150 4738 5154 4742
rect 166 4728 170 4732
rect 1134 4728 1138 4732
rect 1270 4728 1274 4732
rect 1326 4728 1330 4732
rect 1870 4728 1874 4732
rect 1902 4728 1906 4732
rect 2030 4728 2034 4732
rect 2854 4728 2858 4732
rect 3198 4728 3202 4732
rect 3302 4728 3306 4732
rect 3750 4728 3754 4732
rect 4814 4728 4818 4732
rect 174 4718 178 4722
rect 302 4718 306 4722
rect 462 4718 466 4722
rect 918 4718 922 4722
rect 1126 4718 1130 4722
rect 1166 4718 1170 4722
rect 1198 4718 1202 4722
rect 1302 4718 1306 4722
rect 1454 4718 1458 4722
rect 1566 4718 1570 4722
rect 1710 4718 1714 4722
rect 1846 4718 1850 4722
rect 1998 4718 2002 4722
rect 2014 4718 2018 4722
rect 2166 4718 2170 4722
rect 2686 4718 2690 4722
rect 2862 4718 2866 4722
rect 2958 4718 2962 4722
rect 3054 4718 3058 4722
rect 3078 4718 3082 4722
rect 3182 4718 3186 4722
rect 3206 4718 3210 4722
rect 3566 4718 3570 4722
rect 3654 4718 3658 4722
rect 3814 4718 3818 4722
rect 3990 4718 3994 4722
rect 4302 4718 4306 4722
rect 4326 4718 4330 4722
rect 4510 4718 4514 4722
rect 4638 4718 4642 4722
rect 4694 4718 4698 4722
rect 4718 4718 4722 4722
rect 4870 4718 4874 4722
rect 4998 4718 5002 4722
rect 5094 4718 5098 4722
rect 1050 4703 1054 4707
rect 1057 4703 1061 4707
rect 2074 4703 2078 4707
rect 2081 4703 2085 4707
rect 3098 4703 3102 4707
rect 3105 4703 3109 4707
rect 4114 4703 4118 4707
rect 4121 4703 4125 4707
rect 94 4688 98 4692
rect 342 4688 346 4692
rect 398 4688 402 4692
rect 1158 4688 1162 4692
rect 1262 4688 1266 4692
rect 1334 4688 1338 4692
rect 1430 4688 1434 4692
rect 1606 4688 1610 4692
rect 2054 4688 2058 4692
rect 2102 4688 2106 4692
rect 2350 4688 2354 4692
rect 3118 4688 3122 4692
rect 3182 4688 3186 4692
rect 3294 4688 3298 4692
rect 3534 4688 3538 4692
rect 4038 4688 4042 4692
rect 4086 4688 4090 4692
rect 4166 4688 4170 4692
rect 4390 4688 4394 4692
rect 4470 4688 4474 4692
rect 4606 4688 4610 4692
rect 4662 4688 4666 4692
rect 4766 4688 4770 4692
rect 5014 4688 5018 4692
rect 14 4668 18 4672
rect 110 4668 114 4672
rect 118 4668 122 4672
rect 134 4678 138 4682
rect 430 4678 434 4682
rect 470 4678 474 4682
rect 686 4678 690 4682
rect 782 4678 786 4682
rect 798 4678 802 4682
rect 886 4678 890 4682
rect 166 4668 170 4672
rect 214 4668 218 4672
rect 254 4668 258 4672
rect 310 4668 314 4672
rect 318 4668 322 4672
rect 374 4668 378 4672
rect 390 4668 394 4672
rect 438 4668 442 4672
rect 486 4668 490 4672
rect 518 4668 522 4672
rect 534 4668 538 4672
rect 566 4668 570 4672
rect 654 4668 658 4672
rect 742 4668 746 4672
rect 814 4668 818 4672
rect 838 4668 842 4672
rect 846 4668 850 4672
rect 942 4668 946 4672
rect 1022 4668 1026 4672
rect 1070 4668 1074 4672
rect 1086 4668 1090 4672
rect 1150 4668 1154 4672
rect 1174 4678 1178 4682
rect 1230 4678 1234 4682
rect 1238 4678 1242 4682
rect 1254 4668 1258 4672
rect 1278 4678 1282 4682
rect 1638 4678 1642 4682
rect 1654 4678 1658 4682
rect 2022 4678 2026 4682
rect 2238 4678 2242 4682
rect 2270 4678 2274 4682
rect 2286 4678 2290 4682
rect 2710 4678 2714 4682
rect 2766 4678 2770 4682
rect 3150 4678 3154 4682
rect 3230 4678 3234 4682
rect 3430 4678 3434 4682
rect 3550 4678 3554 4682
rect 3574 4678 3578 4682
rect 3806 4678 3810 4682
rect 3878 4678 3882 4682
rect 4078 4678 4082 4682
rect 4422 4678 4426 4682
rect 4510 4678 4514 4682
rect 4726 4678 4730 4682
rect 4854 4678 4858 4682
rect 5150 4678 5154 4682
rect 1302 4668 1306 4672
rect 1454 4668 1458 4672
rect 1470 4668 1474 4672
rect 1558 4668 1562 4672
rect 1702 4668 1706 4672
rect 1766 4668 1770 4672
rect 1822 4668 1826 4672
rect 1910 4668 1914 4672
rect 1950 4668 1954 4672
rect 38 4658 42 4662
rect 102 4658 106 4662
rect 150 4658 154 4662
rect 190 4658 194 4662
rect 262 4658 266 4662
rect 302 4658 306 4662
rect 326 4658 330 4662
rect 366 4658 370 4662
rect 382 4658 386 4662
rect 414 4658 418 4662
rect 462 4658 466 4662
rect 494 4658 498 4662
rect 590 4658 594 4662
rect 654 4658 658 4662
rect 678 4658 682 4662
rect 702 4658 706 4662
rect 710 4658 714 4662
rect 734 4658 738 4662
rect 758 4658 762 4662
rect 766 4658 770 4662
rect 822 4658 826 4662
rect 854 4658 858 4662
rect 902 4658 906 4662
rect 934 4659 938 4663
rect 1078 4658 1082 4662
rect 1142 4658 1146 4662
rect 1190 4658 1194 4662
rect 1198 4658 1202 4662
rect 1214 4658 1218 4662
rect 1246 4658 1250 4662
rect 1302 4658 1306 4662
rect 1310 4658 1314 4662
rect 1374 4658 1378 4662
rect 1390 4658 1394 4662
rect 1446 4658 1450 4662
rect 1494 4658 1498 4662
rect 1582 4658 1586 4662
rect 1598 4658 1602 4662
rect 1622 4658 1626 4662
rect 1702 4658 1706 4662
rect 1774 4658 1778 4662
rect 1790 4658 1794 4662
rect 1814 4658 1818 4662
rect 1894 4659 1898 4663
rect 1982 4668 1986 4672
rect 1998 4668 2002 4672
rect 2062 4668 2066 4672
rect 2134 4668 2138 4672
rect 2230 4668 2234 4672
rect 2270 4668 2274 4672
rect 2326 4668 2330 4672
rect 2366 4668 2370 4672
rect 2422 4668 2426 4672
rect 2510 4668 2514 4672
rect 2526 4668 2530 4672
rect 2566 4668 2570 4672
rect 2582 4668 2586 4672
rect 2726 4668 2730 4672
rect 2782 4668 2786 4672
rect 2878 4668 2882 4672
rect 3014 4668 3018 4672
rect 3062 4668 3066 4672
rect 3094 4668 3098 4672
rect 3142 4668 3146 4672
rect 3190 4668 3194 4672
rect 3366 4668 3370 4672
rect 3382 4668 3386 4672
rect 3398 4668 3402 4672
rect 3422 4668 3426 4672
rect 3486 4668 3490 4672
rect 3614 4668 3618 4672
rect 3694 4668 3698 4672
rect 3734 4668 3738 4672
rect 3934 4668 3938 4672
rect 3942 4668 3946 4672
rect 3966 4668 3970 4672
rect 4006 4668 4010 4672
rect 4062 4668 4066 4672
rect 4110 4668 4114 4672
rect 4158 4668 4162 4672
rect 4190 4668 4194 4672
rect 4278 4668 4282 4672
rect 4318 4668 4322 4672
rect 1942 4658 1946 4662
rect 1958 4658 1962 4662
rect 1974 4658 1978 4662
rect 2014 4658 2018 4662
rect 2038 4658 2042 4662
rect 2070 4658 2074 4662
rect 2118 4658 2122 4662
rect 2158 4658 2162 4662
rect 2254 4658 2258 4662
rect 2302 4658 2306 4662
rect 2334 4658 2338 4662
rect 2374 4658 2378 4662
rect 2406 4658 2410 4662
rect 2414 4658 2418 4662
rect 2486 4658 2490 4662
rect 2534 4658 2538 4662
rect 2574 4658 2578 4662
rect 2630 4659 2634 4663
rect 2654 4658 2658 4662
rect 2718 4658 2722 4662
rect 2750 4658 2754 4662
rect 2798 4659 2802 4663
rect 2902 4658 2906 4662
rect 2990 4658 2994 4662
rect 3014 4658 3018 4662
rect 3086 4658 3090 4662
rect 3134 4658 3138 4662
rect 3166 4658 3170 4662
rect 3198 4658 3202 4662
rect 3230 4659 3234 4663
rect 3262 4658 3266 4662
rect 3374 4658 3378 4662
rect 3406 4658 3410 4662
rect 3470 4659 3474 4663
rect 3558 4658 3562 4662
rect 3606 4658 3610 4662
rect 3646 4658 3650 4662
rect 3678 4658 3682 4662
rect 3686 4658 3690 4662
rect 3726 4659 3730 4663
rect 3750 4658 3754 4662
rect 3878 4659 3882 4663
rect 3926 4658 3930 4662
rect 3974 4658 3978 4662
rect 3998 4658 4002 4662
rect 4014 4658 4018 4662
rect 4054 4658 4058 4662
rect 4102 4658 4106 4662
rect 4150 4658 4154 4662
rect 4182 4658 4186 4662
rect 4262 4659 4266 4663
rect 4350 4668 4354 4672
rect 4382 4668 4386 4672
rect 4414 4668 4418 4672
rect 4438 4668 4442 4672
rect 4494 4668 4498 4672
rect 4518 4668 4522 4672
rect 4534 4668 4538 4672
rect 4574 4668 4578 4672
rect 4582 4668 4586 4672
rect 4622 4668 4626 4672
rect 4638 4668 4642 4672
rect 4686 4668 4690 4672
rect 4774 4668 4778 4672
rect 4822 4668 4826 4672
rect 4830 4668 4834 4672
rect 4886 4668 4890 4672
rect 4950 4668 4954 4672
rect 4990 4668 4994 4672
rect 5022 4668 5026 4672
rect 5054 4668 5058 4672
rect 4310 4658 4314 4662
rect 4326 4658 4330 4662
rect 4342 4658 4346 4662
rect 4374 4658 4378 4662
rect 4406 4658 4410 4662
rect 4446 4658 4450 4662
rect 4486 4658 4490 4662
rect 4526 4658 4530 4662
rect 4566 4658 4570 4662
rect 4590 4658 4594 4662
rect 4638 4658 4642 4662
rect 4678 4658 4682 4662
rect 4710 4658 4714 4662
rect 4750 4658 4754 4662
rect 4814 4658 4818 4662
rect 4838 4658 4842 4662
rect 4878 4658 4882 4662
rect 4942 4658 4946 4662
rect 4990 4658 4994 4662
rect 5030 4658 5034 4662
rect 5054 4658 5058 4662
rect 5062 4658 5066 4662
rect 5078 4658 5082 4662
rect 5134 4658 5138 4662
rect 286 4648 290 4652
rect 350 4648 354 4652
rect 518 4648 522 4652
rect 678 4648 682 4652
rect 774 4648 778 4652
rect 838 4648 842 4652
rect 854 4648 858 4652
rect 1006 4648 1010 4652
rect 1014 4648 1018 4652
rect 1198 4648 1202 4652
rect 1326 4648 1330 4652
rect 1430 4648 1434 4652
rect 1598 4648 1602 4652
rect 1606 4648 1610 4652
rect 1790 4648 1794 4652
rect 1814 4648 1818 4652
rect 1942 4648 1946 4652
rect 1958 4648 1962 4652
rect 2238 4648 2242 4652
rect 2550 4648 2554 4652
rect 2742 4648 2746 4652
rect 3006 4648 3010 4652
rect 3046 4648 3050 4652
rect 3086 4648 3090 4652
rect 3118 4648 3122 4652
rect 3278 4648 3282 4652
rect 3590 4648 3594 4652
rect 3662 4648 3666 4652
rect 3910 4648 3914 4652
rect 3942 4648 3946 4652
rect 4030 4648 4034 4652
rect 4086 4648 4090 4652
rect 4134 4648 4138 4652
rect 4166 4648 4170 4652
rect 4294 4648 4298 4652
rect 4326 4648 4330 4652
rect 4358 4648 4362 4652
rect 4390 4648 4394 4652
rect 4462 4648 4466 4652
rect 4550 4648 4554 4652
rect 4606 4648 4610 4652
rect 4614 4648 4618 4652
rect 4654 4648 4658 4652
rect 4694 4648 4698 4652
rect 4790 4648 4794 4652
rect 4798 4648 4802 4652
rect 4862 4648 4866 4652
rect 5014 4648 5018 4652
rect 5046 4648 5050 4652
rect 5078 4648 5082 4652
rect 246 4638 250 4642
rect 262 4638 266 4642
rect 870 4638 874 4642
rect 998 4638 1002 4642
rect 1134 4638 1138 4642
rect 1798 4638 1802 4642
rect 1830 4638 1834 4642
rect 1926 4638 1930 4642
rect 2390 4638 2394 4642
rect 2430 4638 2434 4642
rect 2694 4638 2698 4642
rect 2846 4638 2850 4642
rect 2862 4638 2866 4642
rect 2990 4638 2994 4642
rect 3062 4638 3066 4642
rect 3518 4638 3522 4642
rect 3926 4638 3930 4642
rect 4150 4638 4154 4642
rect 4310 4638 4314 4642
rect 4374 4638 4378 4642
rect 4422 4638 4426 4642
rect 4894 4638 4898 4642
rect 5086 4628 5090 4632
rect 478 4618 482 4622
rect 646 4618 650 4622
rect 694 4618 698 4622
rect 726 4618 730 4622
rect 790 4618 794 4622
rect 806 4618 810 4622
rect 1310 4618 1314 4622
rect 1550 4618 1554 4622
rect 1646 4618 1650 4622
rect 1662 4618 1666 4622
rect 1758 4618 1762 4622
rect 2102 4618 2106 4622
rect 2230 4618 2234 4622
rect 2278 4618 2282 4622
rect 2294 4618 2298 4622
rect 2702 4618 2706 4622
rect 2974 4618 2978 4622
rect 3022 4618 3026 4622
rect 3310 4618 3314 4622
rect 3438 4618 3442 4622
rect 3534 4618 3538 4622
rect 3542 4618 3546 4622
rect 3606 4618 3610 4622
rect 3790 4618 3794 4622
rect 3798 4618 3802 4622
rect 3814 4618 3818 4622
rect 3982 4618 3986 4622
rect 4070 4618 4074 4622
rect 4198 4618 4202 4622
rect 4502 4618 4506 4622
rect 4710 4618 4714 4622
rect 4814 4618 4818 4622
rect 538 4603 542 4607
rect 545 4603 549 4607
rect 1562 4603 1566 4607
rect 1569 4603 1573 4607
rect 2586 4603 2590 4607
rect 2593 4603 2597 4607
rect 3610 4603 3614 4607
rect 3617 4603 3621 4607
rect 4634 4603 4638 4607
rect 4641 4603 4645 4607
rect 262 4588 266 4592
rect 670 4588 674 4592
rect 1446 4588 1450 4592
rect 1606 4588 1610 4592
rect 2982 4588 2986 4592
rect 3030 4588 3034 4592
rect 5078 4588 5082 4592
rect 646 4578 650 4582
rect 278 4568 282 4572
rect 654 4568 658 4572
rect 766 4568 770 4572
rect 830 4568 834 4572
rect 942 4568 946 4572
rect 958 4568 962 4572
rect 1422 4568 1426 4572
rect 1590 4568 1594 4572
rect 1966 4568 1970 4572
rect 2086 4568 2090 4572
rect 2238 4568 2242 4572
rect 3054 4568 3058 4572
rect 3750 4568 3754 4572
rect 4078 4568 4082 4572
rect 4134 4568 4138 4572
rect 4246 4568 4250 4572
rect 4286 4568 4290 4572
rect 4390 4568 4394 4572
rect 4398 4568 4402 4572
rect 4414 4568 4418 4572
rect 4470 4568 4474 4572
rect 4558 4568 4562 4572
rect 4582 4568 4586 4572
rect 4734 4568 4738 4572
rect 4742 4568 4746 4572
rect 4934 4568 4938 4572
rect 6 4548 10 4552
rect 54 4548 58 4552
rect 94 4548 98 4552
rect 190 4548 194 4552
rect 278 4548 282 4552
rect 302 4558 306 4562
rect 350 4558 354 4562
rect 334 4548 338 4552
rect 718 4558 722 4562
rect 366 4548 370 4552
rect 374 4548 378 4552
rect 414 4547 418 4551
rect 486 4548 490 4552
rect 518 4548 522 4552
rect 590 4548 594 4552
rect 670 4548 674 4552
rect 686 4548 690 4552
rect 750 4548 754 4552
rect 790 4548 794 4552
rect 814 4548 818 4552
rect 966 4558 970 4562
rect 1198 4558 1202 4562
rect 1214 4558 1218 4562
rect 1246 4558 1250 4562
rect 1926 4558 1930 4562
rect 1942 4558 1946 4562
rect 1950 4558 1954 4562
rect 1990 4558 1994 4562
rect 2166 4558 2170 4562
rect 2190 4558 2194 4562
rect 2222 4558 2226 4562
rect 2462 4558 2466 4562
rect 854 4548 858 4552
rect 894 4547 898 4551
rect 1030 4548 1034 4552
rect 1134 4548 1138 4552
rect 1158 4548 1162 4552
rect 1230 4548 1234 4552
rect 1294 4548 1298 4552
rect 1350 4548 1354 4552
rect 1382 4548 1386 4552
rect 1446 4548 1450 4552
rect 1494 4548 1498 4552
rect 1606 4548 1610 4552
rect 1622 4548 1626 4552
rect 1670 4548 1674 4552
rect 1710 4548 1714 4552
rect 1798 4548 1802 4552
rect 1886 4547 1890 4551
rect 1926 4548 1930 4552
rect 2030 4548 2034 4552
rect 2134 4548 2138 4552
rect 2158 4548 2162 4552
rect 2206 4548 2210 4552
rect 2278 4548 2282 4552
rect 2390 4548 2394 4552
rect 2422 4547 2426 4551
rect 2454 4548 2458 4552
rect 2462 4548 2466 4552
rect 2486 4558 2490 4562
rect 2526 4558 2530 4562
rect 2566 4558 2570 4562
rect 2702 4558 2706 4562
rect 2718 4558 2722 4562
rect 2950 4558 2954 4562
rect 2990 4558 2994 4562
rect 3014 4558 3018 4562
rect 2526 4548 2530 4552
rect 46 4538 50 4542
rect 70 4538 74 4542
rect 166 4538 170 4542
rect 318 4538 322 4542
rect 326 4538 330 4542
rect 382 4538 386 4542
rect 398 4538 402 4542
rect 494 4538 498 4542
rect 566 4538 570 4542
rect 614 4538 618 4542
rect 678 4538 682 4542
rect 702 4538 706 4542
rect 734 4538 738 4542
rect 742 4538 746 4542
rect 774 4538 778 4542
rect 798 4538 802 4542
rect 806 4538 810 4542
rect 846 4538 850 4542
rect 862 4538 866 4542
rect 878 4538 882 4542
rect 982 4538 986 4542
rect 1070 4538 1074 4542
rect 1214 4538 1218 4542
rect 1222 4538 1226 4542
rect 1286 4538 1290 4542
rect 1358 4538 1362 4542
rect 1374 4538 1378 4542
rect 1406 4538 1410 4542
rect 1454 4538 1458 4542
rect 1470 4538 1474 4542
rect 1614 4538 1618 4542
rect 1630 4538 1634 4542
rect 1638 4538 1642 4542
rect 1686 4538 1690 4542
rect 1774 4538 1778 4542
rect 1790 4538 1794 4542
rect 1798 4538 1802 4542
rect 1902 4538 1906 4542
rect 1918 4538 1922 4542
rect 1966 4538 1970 4542
rect 1974 4538 1978 4542
rect 2102 4538 2106 4542
rect 2126 4538 2130 4542
rect 2182 4538 2186 4542
rect 2222 4538 2226 4542
rect 2238 4538 2242 4542
rect 2270 4538 2274 4542
rect 2342 4538 2346 4542
rect 2350 4538 2354 4542
rect 2606 4547 2610 4551
rect 2686 4548 2690 4552
rect 2702 4548 2706 4552
rect 2710 4548 2714 4552
rect 2798 4548 2802 4552
rect 2862 4547 2866 4551
rect 3030 4548 3034 4552
rect 3086 4558 3090 4562
rect 3278 4558 3282 4562
rect 3302 4558 3306 4562
rect 3350 4558 3354 4562
rect 3502 4558 3506 4562
rect 3510 4558 3514 4562
rect 3550 4558 3554 4562
rect 3646 4558 3650 4562
rect 3910 4558 3914 4562
rect 3942 4558 3946 4562
rect 3078 4548 3082 4552
rect 3142 4548 3146 4552
rect 3158 4548 3162 4552
rect 3174 4548 3178 4552
rect 3238 4548 3242 4552
rect 3318 4548 3322 4552
rect 3358 4548 3362 4552
rect 3406 4547 3410 4551
rect 3486 4548 3490 4552
rect 3566 4548 3570 4552
rect 3598 4547 3602 4551
rect 3638 4548 3642 4552
rect 3662 4548 3666 4552
rect 3710 4548 3714 4552
rect 3806 4548 3810 4552
rect 3830 4548 3834 4552
rect 3886 4548 3890 4552
rect 3902 4548 3906 4552
rect 3926 4548 3930 4552
rect 4014 4558 4018 4562
rect 4086 4558 4090 4562
rect 3966 4548 3970 4552
rect 3982 4548 3986 4552
rect 4006 4548 4010 4552
rect 4038 4548 4042 4552
rect 4086 4548 4090 4552
rect 4102 4548 4106 4552
rect 4190 4548 4194 4552
rect 4446 4558 4450 4562
rect 4478 4558 4482 4562
rect 4518 4558 4522 4562
rect 4534 4558 4538 4562
rect 4838 4558 4842 4562
rect 4894 4558 4898 4562
rect 4270 4548 4274 4552
rect 4302 4548 4306 4552
rect 4430 4548 4434 4552
rect 4494 4548 4498 4552
rect 4534 4548 4538 4552
rect 4566 4548 4570 4552
rect 4662 4548 4666 4552
rect 4686 4547 4690 4551
rect 4806 4547 4810 4551
rect 4838 4548 4842 4552
rect 4862 4548 4866 4552
rect 4878 4548 4882 4552
rect 5054 4558 5058 4562
rect 4910 4548 4914 4552
rect 4918 4548 4922 4552
rect 4990 4548 4994 4552
rect 5038 4548 5042 4552
rect 5166 4558 5170 4562
rect 5078 4548 5082 4552
rect 2502 4538 2506 4542
rect 2510 4538 2514 4542
rect 2534 4538 2538 4542
rect 2574 4538 2578 4542
rect 2590 4538 2594 4542
rect 2614 4538 2618 4542
rect 2678 4538 2682 4542
rect 2710 4538 2714 4542
rect 2846 4538 2850 4542
rect 2966 4538 2970 4542
rect 2974 4538 2978 4542
rect 2998 4538 3002 4542
rect 3022 4538 3026 4542
rect 3078 4538 3082 4542
rect 3102 4538 3106 4542
rect 3166 4538 3170 4542
rect 3262 4538 3266 4542
rect 3294 4538 3298 4542
rect 3318 4538 3322 4542
rect 3334 4538 3338 4542
rect 3390 4538 3394 4542
rect 3478 4538 3482 4542
rect 3494 4538 3498 4542
rect 3526 4538 3530 4542
rect 3670 4538 3674 4542
rect 3686 4538 3690 4542
rect 3918 4538 3922 4542
rect 3974 4538 3978 4542
rect 3982 4538 3986 4542
rect 4062 4538 4066 4542
rect 4110 4538 4114 4542
rect 4214 4538 4218 4542
rect 4230 4538 4234 4542
rect 4278 4538 4282 4542
rect 4302 4538 4306 4542
rect 4374 4538 4378 4542
rect 4398 4538 4402 4542
rect 4422 4538 4426 4542
rect 4454 4538 4458 4542
rect 4502 4538 4506 4542
rect 4510 4538 4514 4542
rect 4542 4538 4546 4542
rect 4566 4538 4570 4542
rect 4718 4538 4722 4542
rect 4822 4538 4826 4542
rect 4862 4538 4866 4542
rect 4870 4538 4874 4542
rect 4926 4538 4930 4542
rect 22 4528 26 4532
rect 550 4528 554 4532
rect 1246 4528 1250 4532
rect 1398 4528 1402 4532
rect 1582 4528 1586 4532
rect 1654 4528 1658 4532
rect 1774 4528 1778 4532
rect 1814 4528 1818 4532
rect 2022 4528 2026 4532
rect 2110 4528 2114 4532
rect 2142 4528 2146 4532
rect 2158 4528 2162 4532
rect 2806 4528 2810 4532
rect 3126 4528 3130 4532
rect 3374 4528 3378 4532
rect 5030 4538 5034 4542
rect 5086 4538 5090 4542
rect 5094 4538 5098 4542
rect 5158 4538 5162 4542
rect 5182 4538 5186 4542
rect 4014 4528 4018 4532
rect 4390 4528 4394 4532
rect 4614 4528 4618 4532
rect 4734 4528 4738 4532
rect 4966 4528 4970 4532
rect 4998 4528 5002 4532
rect 38 4518 42 4522
rect 150 4518 154 4522
rect 478 4518 482 4522
rect 502 4518 506 4522
rect 726 4518 730 4522
rect 974 4518 978 4522
rect 990 4518 994 4522
rect 1190 4518 1194 4522
rect 1342 4518 1346 4522
rect 1414 4518 1418 4522
rect 1550 4518 1554 4522
rect 1558 4518 1562 4522
rect 1766 4518 1770 4522
rect 1822 4518 1826 4522
rect 1990 4518 1994 4522
rect 2174 4518 2178 4522
rect 2190 4518 2194 4522
rect 2334 4518 2338 4522
rect 2358 4518 2362 4522
rect 2518 4518 2522 4522
rect 2670 4518 2674 4522
rect 2742 4518 2746 4522
rect 2942 4518 2946 4522
rect 2958 4518 2962 4522
rect 3006 4518 3010 4522
rect 3086 4518 3090 4522
rect 3182 4518 3186 4522
rect 3286 4518 3290 4522
rect 3302 4518 3306 4522
rect 3470 4518 3474 4522
rect 3510 4518 3514 4522
rect 3534 4518 3538 4522
rect 3766 4518 3770 4522
rect 3878 4518 3882 4522
rect 3950 4518 3954 4522
rect 4054 4518 4058 4522
rect 4254 4518 4258 4522
rect 4286 4518 4290 4522
rect 4446 4518 4450 4522
rect 4470 4518 4474 4522
rect 4478 4518 4482 4522
rect 4590 4518 4594 4522
rect 4606 4518 4610 4522
rect 5174 4518 5178 4522
rect 1050 4503 1054 4507
rect 1057 4503 1061 4507
rect 2074 4503 2078 4507
rect 2081 4503 2085 4507
rect 3098 4503 3102 4507
rect 3105 4503 3109 4507
rect 4114 4503 4118 4507
rect 4121 4503 4125 4507
rect 94 4488 98 4492
rect 118 4488 122 4492
rect 286 4488 290 4492
rect 550 4488 554 4492
rect 750 4488 754 4492
rect 1134 4488 1138 4492
rect 1182 4488 1186 4492
rect 1606 4488 1610 4492
rect 2006 4488 2010 4492
rect 2222 4488 2226 4492
rect 2430 4488 2434 4492
rect 2566 4488 2570 4492
rect 2678 4488 2682 4492
rect 2798 4488 2802 4492
rect 2830 4488 2834 4492
rect 3502 4488 3506 4492
rect 3726 4488 3730 4492
rect 3758 4488 3762 4492
rect 3910 4488 3914 4492
rect 4062 4488 4066 4492
rect 4390 4488 4394 4492
rect 4654 4488 4658 4492
rect 4710 4488 4714 4492
rect 4798 4488 4802 4492
rect 4862 4488 4866 4492
rect 5174 4488 5178 4492
rect 150 4478 154 4482
rect 214 4478 218 4482
rect 382 4478 386 4482
rect 766 4478 770 4482
rect 1350 4478 1354 4482
rect 1750 4478 1754 4482
rect 1766 4478 1770 4482
rect 1806 4478 1810 4482
rect 2390 4478 2394 4482
rect 2534 4478 2538 4482
rect 2614 4478 2618 4482
rect 3158 4478 3162 4482
rect 3398 4478 3402 4482
rect 3606 4478 3610 4482
rect 3766 4478 3770 4482
rect 3942 4478 3946 4482
rect 4014 4478 4018 4482
rect 4326 4478 4330 4482
rect 4630 4478 4634 4482
rect 4782 4478 4786 4482
rect 14 4468 18 4472
rect 110 4468 114 4472
rect 166 4468 170 4472
rect 254 4468 258 4472
rect 334 4468 338 4472
rect 406 4468 410 4472
rect 422 4468 426 4472
rect 454 4468 458 4472
rect 494 4468 498 4472
rect 574 4468 578 4472
rect 614 4468 618 4472
rect 702 4468 706 4472
rect 734 4468 738 4472
rect 782 4468 786 4472
rect 870 4468 874 4472
rect 926 4468 930 4472
rect 982 4468 986 4472
rect 1014 4468 1018 4472
rect 1094 4468 1098 4472
rect 1102 4468 1106 4472
rect 1158 4468 1162 4472
rect 1166 4468 1170 4472
rect 1190 4468 1194 4472
rect 1238 4468 1242 4472
rect 1422 4468 1426 4472
rect 1502 4468 1506 4472
rect 1510 4468 1514 4472
rect 1598 4468 1602 4472
rect 1622 4468 1626 4472
rect 1646 4468 1650 4472
rect 1686 4468 1690 4472
rect 1798 4468 1802 4472
rect 1838 4468 1842 4472
rect 1918 4468 1922 4472
rect 1934 4468 1938 4472
rect 1950 4468 1954 4472
rect 1958 4468 1962 4472
rect 1982 4468 1986 4472
rect 2038 4468 2042 4472
rect 2238 4468 2242 4472
rect 2294 4468 2298 4472
rect 2342 4468 2346 4472
rect 2374 4468 2378 4472
rect 2422 4468 2426 4472
rect 2454 4468 2458 4472
rect 38 4458 42 4462
rect 102 4458 106 4462
rect 134 4458 138 4462
rect 190 4458 194 4462
rect 262 4458 266 4462
rect 350 4459 354 4463
rect 398 4458 402 4462
rect 430 4458 434 4462
rect 502 4458 506 4462
rect 518 4458 522 4462
rect 582 4458 586 4462
rect 590 4458 594 4462
rect 630 4459 634 4463
rect 710 4458 714 4462
rect 806 4458 810 4462
rect 878 4458 882 4462
rect 918 4458 922 4462
rect 934 4458 938 4462
rect 942 4458 946 4462
rect 966 4458 970 4462
rect 982 4458 986 4462
rect 1014 4458 1018 4462
rect 1038 4458 1042 4462
rect 1110 4458 1114 4462
rect 1166 4458 1170 4462
rect 1222 4458 1226 4462
rect 1230 4458 1234 4462
rect 1270 4459 1274 4463
rect 1294 4458 1298 4462
rect 1430 4458 1434 4462
rect 1438 4458 1442 4462
rect 1494 4458 1498 4462
rect 1622 4458 1626 4462
rect 1678 4459 1682 4463
rect 1766 4458 1770 4462
rect 1798 4458 1802 4462
rect 1846 4458 1850 4462
rect 1854 4458 1858 4462
rect 1910 4458 1914 4462
rect 1942 4458 1946 4462
rect 1966 4458 1970 4462
rect 1990 4458 1994 4462
rect 1998 4458 2002 4462
rect 2022 4458 2026 4462
rect 2030 4458 2034 4462
rect 2150 4459 2154 4463
rect 2518 4468 2522 4472
rect 2526 4468 2530 4472
rect 2542 4468 2546 4472
rect 2686 4468 2690 4472
rect 2734 4468 2738 4472
rect 2742 4468 2746 4472
rect 2790 4468 2794 4472
rect 2822 4468 2826 4472
rect 2894 4468 2898 4472
rect 2942 4468 2946 4472
rect 2974 4468 2978 4472
rect 3198 4468 3202 4472
rect 3254 4468 3258 4472
rect 3382 4468 3386 4472
rect 3414 4468 3418 4472
rect 3486 4468 3490 4472
rect 3534 4468 3538 4472
rect 3542 4468 3546 4472
rect 3598 4468 3602 4472
rect 3670 4468 3674 4472
rect 3734 4468 3738 4472
rect 3806 4468 3810 4472
rect 3870 4468 3874 4472
rect 3902 4468 3906 4472
rect 3926 4468 3930 4472
rect 4118 4468 4122 4472
rect 4126 4468 4130 4472
rect 4142 4468 4146 4472
rect 4214 4468 4218 4472
rect 4294 4468 4298 4472
rect 4398 4468 4402 4472
rect 4454 4468 4458 4472
rect 4462 4468 4466 4472
rect 4486 4468 4490 4472
rect 4518 4468 4522 4472
rect 4670 4468 4674 4472
rect 4702 4468 4706 4472
rect 4734 4468 4738 4472
rect 4822 4468 4826 4472
rect 4870 4468 4874 4472
rect 4934 4468 4938 4472
rect 4998 4468 5002 4472
rect 5022 4468 5026 4472
rect 5062 4468 5066 4472
rect 5078 4468 5082 4472
rect 5094 4468 5098 4472
rect 2182 4458 2186 4462
rect 2246 4458 2250 4462
rect 2254 4458 2258 4462
rect 2278 4458 2282 4462
rect 2302 4458 2306 4462
rect 2366 4458 2370 4462
rect 2414 4458 2418 4462
rect 2446 4458 2450 4462
rect 2478 4458 2482 4462
rect 2486 4458 2490 4462
rect 2494 4458 2498 4462
rect 2550 4458 2554 4462
rect 2614 4459 2618 4463
rect 2694 4458 2698 4462
rect 2774 4458 2778 4462
rect 2790 4458 2794 4462
rect 2814 4458 2818 4462
rect 2902 4458 2906 4462
rect 2950 4458 2954 4462
rect 2982 4458 2986 4462
rect 3038 4458 3042 4462
rect 3062 4458 3066 4462
rect 3134 4458 3138 4462
rect 3190 4458 3194 4462
rect 3238 4458 3242 4462
rect 3262 4458 3266 4462
rect 3278 4458 3282 4462
rect 3334 4458 3338 4462
rect 3358 4458 3362 4462
rect 3502 4458 3506 4462
rect 3534 4458 3538 4462
rect 3550 4458 3554 4462
rect 3598 4458 3602 4462
rect 3662 4459 3666 4463
rect 3742 4458 3746 4462
rect 3782 4458 3786 4462
rect 3798 4458 3802 4462
rect 3854 4458 3858 4462
rect 3862 4458 3866 4462
rect 3886 4458 3890 4462
rect 3902 4458 3906 4462
rect 3998 4458 4002 4462
rect 4046 4458 4050 4462
rect 4054 4458 4058 4462
rect 4078 4458 4082 4462
rect 4094 4458 4098 4462
rect 4150 4458 4154 4462
rect 4158 4458 4162 4462
rect 4206 4458 4210 4462
rect 4270 4458 4274 4462
rect 4294 4458 4298 4462
rect 4334 4458 4338 4462
rect 4406 4458 4410 4462
rect 4446 4458 4450 4462
rect 4470 4458 4474 4462
rect 4510 4458 4514 4462
rect 4566 4458 4570 4462
rect 4582 4458 4586 4462
rect 4694 4458 4698 4462
rect 4726 4458 4730 4462
rect 4758 4458 4762 4462
rect 4814 4458 4818 4462
rect 4846 4458 4850 4462
rect 4886 4458 4890 4462
rect 4934 4458 4938 4462
rect 4990 4458 4994 4462
rect 5054 4458 5058 4462
rect 5110 4459 5114 4463
rect 262 4448 266 4452
rect 278 4448 282 4452
rect 438 4448 442 4452
rect 446 4448 450 4452
rect 598 4448 602 4452
rect 726 4448 730 4452
rect 1006 4448 1010 4452
rect 1126 4448 1130 4452
rect 1182 4448 1186 4452
rect 1206 4448 1210 4452
rect 1478 4448 1482 4452
rect 1614 4448 1618 4452
rect 1646 4448 1650 4452
rect 1774 4448 1778 4452
rect 1822 4448 1826 4452
rect 1838 4448 1842 4452
rect 1894 4448 1898 4452
rect 2222 4448 2226 4452
rect 2326 4448 2330 4452
rect 2350 4448 2354 4452
rect 2390 4448 2394 4452
rect 2414 4448 2418 4452
rect 2430 4448 2434 4452
rect 2462 4448 2466 4452
rect 2718 4448 2722 4452
rect 2758 4448 2762 4452
rect 2798 4448 2802 4452
rect 2966 4448 2970 4452
rect 2998 4448 3002 4452
rect 3118 4448 3122 4452
rect 3214 4448 3218 4452
rect 3238 4448 3242 4452
rect 3278 4448 3282 4452
rect 3510 4448 3514 4452
rect 3566 4448 3570 4452
rect 3758 4448 3762 4452
rect 3782 4448 3786 4452
rect 3838 4448 3842 4452
rect 3878 4448 3882 4452
rect 3910 4448 3914 4452
rect 4166 4448 4170 4452
rect 4430 4448 4434 4452
rect 4494 4448 4498 4452
rect 4654 4448 4658 4452
rect 4678 4448 4682 4452
rect 4694 4448 4698 4452
rect 4710 4448 4714 4452
rect 4742 4448 4746 4452
rect 4838 4448 4842 4452
rect 4902 4448 4906 4452
rect 4926 4448 4930 4452
rect 5038 4448 5042 4452
rect 5054 4448 5058 4452
rect 678 4438 682 4442
rect 750 4438 754 4442
rect 862 4438 866 4442
rect 902 4438 906 4442
rect 1726 4438 1730 4442
rect 1926 4438 1930 4442
rect 2478 4438 2482 4442
rect 2574 4438 2578 4442
rect 3590 4438 3594 4442
rect 3942 4438 3946 4442
rect 3966 4438 3970 4442
rect 4374 4438 4378 4442
rect 4406 4438 4410 4442
rect 4822 4438 4826 4442
rect 878 4428 882 4432
rect 2302 4428 2306 4432
rect 2950 4428 2954 4432
rect 94 4418 98 4422
rect 246 4418 250 4422
rect 566 4418 570 4422
rect 694 4418 698 4422
rect 710 4418 714 4422
rect 958 4418 962 4422
rect 1086 4418 1090 4422
rect 1366 4418 1370 4422
rect 1454 4418 1458 4422
rect 1566 4418 1570 4422
rect 1742 4418 1746 4422
rect 1790 4418 1794 4422
rect 1814 4418 1818 4422
rect 1862 4418 1866 4422
rect 2094 4418 2098 4422
rect 2214 4418 2218 4422
rect 2270 4418 2274 4422
rect 2366 4418 2370 4422
rect 2382 4418 2386 4422
rect 2694 4418 2698 4422
rect 2982 4418 2986 4422
rect 3006 4418 3010 4422
rect 3134 4418 3138 4422
rect 3174 4418 3178 4422
rect 3262 4418 3266 4422
rect 3406 4418 3410 4422
rect 3470 4418 3474 4422
rect 3526 4418 3530 4422
rect 3630 4418 3634 4422
rect 3774 4418 3778 4422
rect 4262 4418 4266 4422
rect 4526 4418 4530 4422
rect 4622 4418 4626 4422
rect 4758 4418 4762 4422
rect 4862 4418 4866 4422
rect 4942 4418 4946 4422
rect 538 4403 542 4407
rect 545 4403 549 4407
rect 1562 4403 1566 4407
rect 1569 4403 1573 4407
rect 2586 4403 2590 4407
rect 2593 4403 2597 4407
rect 3610 4403 3614 4407
rect 3617 4403 3621 4407
rect 4634 4403 4638 4407
rect 4641 4403 4645 4407
rect 254 4388 258 4392
rect 1030 4388 1034 4392
rect 1334 4388 1338 4392
rect 1694 4388 1698 4392
rect 2062 4388 2066 4392
rect 2462 4388 2466 4392
rect 2782 4388 2786 4392
rect 2822 4388 2826 4392
rect 3678 4388 3682 4392
rect 4102 4388 4106 4392
rect 4278 4388 4282 4392
rect 4542 4388 4546 4392
rect 5014 4388 5018 4392
rect 742 4378 746 4382
rect 622 4368 626 4372
rect 766 4368 770 4372
rect 798 4368 802 4372
rect 990 4368 994 4372
rect 1470 4368 1474 4372
rect 1710 4368 1714 4372
rect 1806 4368 1810 4372
rect 1846 4368 1850 4372
rect 2006 4368 2010 4372
rect 2110 4368 2114 4372
rect 2398 4368 2402 4372
rect 190 4358 194 4362
rect 6 4348 10 4352
rect 38 4348 42 4352
rect 54 4348 58 4352
rect 86 4347 90 4351
rect 158 4348 162 4352
rect 230 4348 234 4352
rect 270 4348 274 4352
rect 294 4358 298 4362
rect 318 4358 322 4362
rect 574 4358 578 4362
rect 382 4348 386 4352
rect 398 4348 402 4352
rect 470 4348 474 4352
rect 494 4348 498 4352
rect 574 4348 578 4352
rect 598 4358 602 4362
rect 750 4358 754 4362
rect 614 4348 618 4352
rect 638 4348 642 4352
rect 686 4348 690 4352
rect 774 4348 778 4352
rect 838 4358 842 4362
rect 3446 4368 3450 4372
rect 3622 4368 3626 4372
rect 3646 4368 3650 4372
rect 3790 4368 3794 4372
rect 4046 4368 4050 4372
rect 4166 4368 4170 4372
rect 4342 4368 4346 4372
rect 5182 4368 5186 4372
rect 1006 4358 1010 4362
rect 1014 4358 1018 4362
rect 1182 4358 1186 4362
rect 1230 4358 1234 4362
rect 1486 4358 1490 4362
rect 822 4348 826 4352
rect 886 4347 890 4351
rect 966 4348 970 4352
rect 982 4348 986 4352
rect 1030 4348 1034 4352
rect 1094 4348 1098 4352
rect 1166 4348 1170 4352
rect 1174 4348 1178 4352
rect 1214 4348 1218 4352
rect 1262 4347 1266 4351
rect 1294 4348 1298 4352
rect 1334 4348 1338 4352
rect 1390 4348 1394 4352
rect 1470 4348 1474 4352
rect 1486 4348 1490 4352
rect 1502 4348 1506 4352
rect 46 4338 50 4342
rect 70 4338 74 4342
rect 166 4338 170 4342
rect 206 4338 210 4342
rect 262 4338 266 4342
rect 310 4338 314 4342
rect 334 4338 338 4342
rect 446 4338 450 4342
rect 542 4338 546 4342
rect 614 4338 618 4342
rect 646 4338 650 4342
rect 678 4338 682 4342
rect 766 4338 770 4342
rect 774 4338 778 4342
rect 806 4338 810 4342
rect 830 4338 834 4342
rect 854 4338 858 4342
rect 894 4338 898 4342
rect 958 4338 962 4342
rect 990 4338 994 4342
rect 1038 4338 1042 4342
rect 1070 4338 1074 4342
rect 1094 4338 1098 4342
rect 1158 4338 1162 4342
rect 1206 4338 1210 4342
rect 1230 4338 1234 4342
rect 1246 4338 1250 4342
rect 1366 4338 1370 4342
rect 1478 4338 1482 4342
rect 1598 4347 1602 4351
rect 1646 4348 1650 4352
rect 1686 4348 1690 4352
rect 1694 4348 1698 4352
rect 1750 4348 1754 4352
rect 1822 4348 1826 4352
rect 1830 4348 1834 4352
rect 1910 4358 1914 4362
rect 2078 4358 2082 4362
rect 2134 4358 2138 4362
rect 2190 4358 2194 4362
rect 2470 4358 2474 4362
rect 2478 4358 2482 4362
rect 2534 4358 2538 4362
rect 2582 4358 2586 4362
rect 2718 4358 2722 4362
rect 2790 4358 2794 4362
rect 2878 4358 2882 4362
rect 2894 4358 2898 4362
rect 3134 4358 3138 4362
rect 3150 4358 3154 4362
rect 3190 4358 3194 4362
rect 3350 4358 3354 4362
rect 3430 4358 3434 4362
rect 3462 4358 3466 4362
rect 1870 4348 1874 4352
rect 1902 4348 1906 4352
rect 1966 4348 1970 4352
rect 2062 4348 2066 4352
rect 2086 4348 2090 4352
rect 2110 4348 2114 4352
rect 2150 4348 2154 4352
rect 2278 4347 2282 4351
rect 2334 4347 2338 4351
rect 2406 4348 2410 4352
rect 2414 4348 2418 4352
rect 2438 4348 2442 4352
rect 2478 4348 2482 4352
rect 2494 4348 2498 4352
rect 2510 4348 2514 4352
rect 2542 4348 2546 4352
rect 2630 4347 2634 4351
rect 2662 4348 2666 4352
rect 2734 4348 2738 4352
rect 2758 4348 2762 4352
rect 2774 4348 2778 4352
rect 2798 4348 2802 4352
rect 2846 4348 2850 4352
rect 2966 4347 2970 4351
rect 3046 4348 3050 4352
rect 3150 4348 3154 4352
rect 3174 4348 3178 4352
rect 3270 4348 3274 4352
rect 3398 4347 3402 4351
rect 3446 4348 3450 4352
rect 3462 4348 3466 4352
rect 3478 4348 3482 4352
rect 3526 4348 3530 4352
rect 3542 4348 3546 4352
rect 1518 4338 1522 4342
rect 1582 4338 1586 4342
rect 1630 4338 1634 4342
rect 1654 4338 1658 4342
rect 1670 4338 1674 4342
rect 1678 4338 1682 4342
rect 1726 4338 1730 4342
rect 1766 4338 1770 4342
rect 1814 4338 1818 4342
rect 1870 4338 1874 4342
rect 1926 4338 1930 4342
rect 2046 4338 2050 4342
rect 2054 4338 2058 4342
rect 2094 4338 2098 4342
rect 2134 4338 2138 4342
rect 2142 4338 2146 4342
rect 2158 4338 2162 4342
rect 2174 4338 2178 4342
rect 2262 4338 2266 4342
rect 2454 4338 2458 4342
rect 2502 4338 2506 4342
rect 2518 4338 2522 4342
rect 2566 4338 2570 4342
rect 2590 4338 2594 4342
rect 2702 4338 2706 4342
rect 2718 4338 2722 4342
rect 2774 4338 2778 4342
rect 2838 4338 2842 4342
rect 2854 4338 2858 4342
rect 2878 4338 2882 4342
rect 3038 4338 3042 4342
rect 3078 4338 3082 4342
rect 3126 4338 3130 4342
rect 3166 4338 3170 4342
rect 3198 4338 3202 4342
rect 3246 4338 3250 4342
rect 3294 4338 3298 4342
rect 3310 4338 3314 4342
rect 22 4328 26 4332
rect 182 4328 186 4332
rect 246 4328 250 4332
rect 1190 4328 1194 4332
rect 1350 4328 1354 4332
rect 1382 4328 1386 4332
rect 1886 4328 1890 4332
rect 1958 4328 1962 4332
rect 2558 4328 2562 4332
rect 2814 4328 2818 4332
rect 3414 4338 3418 4342
rect 3454 4338 3458 4342
rect 3742 4347 3746 4351
rect 3830 4348 3834 4352
rect 3854 4348 3858 4352
rect 3894 4348 3898 4352
rect 3926 4358 3930 4362
rect 4030 4358 4034 4362
rect 4086 4358 4090 4362
rect 4134 4358 4138 4362
rect 4294 4358 4298 4362
rect 4350 4358 4354 4362
rect 4390 4358 4394 4362
rect 4494 4358 4498 4362
rect 4574 4358 4578 4362
rect 3942 4348 3946 4352
rect 3974 4348 3978 4352
rect 4054 4348 4058 4352
rect 4102 4348 4106 4352
rect 4134 4348 4138 4352
rect 4158 4348 4162 4352
rect 4222 4348 4226 4352
rect 4262 4348 4266 4352
rect 4310 4348 4314 4352
rect 4366 4348 4370 4352
rect 4430 4348 4434 4352
rect 4454 4348 4458 4352
rect 4510 4348 4514 4352
rect 4726 4358 4730 4362
rect 4742 4358 4746 4362
rect 4758 4358 4762 4362
rect 4790 4358 4794 4362
rect 4822 4358 4826 4362
rect 4878 4358 4882 4362
rect 4598 4348 4602 4352
rect 4662 4348 4666 4352
rect 4694 4347 4698 4351
rect 4742 4348 4746 4352
rect 4758 4348 4762 4352
rect 4774 4348 4778 4352
rect 4798 4348 4802 4352
rect 4806 4348 4810 4352
rect 4838 4348 4842 4352
rect 4854 4348 4858 4352
rect 4862 4348 4866 4352
rect 4902 4358 4906 4362
rect 5054 4358 5058 4362
rect 4902 4348 4906 4352
rect 4974 4348 4978 4352
rect 5038 4348 5042 4352
rect 5070 4348 5074 4352
rect 5078 4348 5082 4352
rect 3486 4338 3490 4342
rect 3502 4338 3506 4342
rect 3590 4338 3594 4342
rect 3630 4338 3634 4342
rect 3654 4338 3658 4342
rect 3718 4338 3722 4342
rect 3758 4338 3762 4342
rect 3774 4338 3778 4342
rect 3894 4338 3898 4342
rect 3910 4338 3914 4342
rect 3950 4338 3954 4342
rect 3998 4338 4002 4342
rect 4006 4338 4010 4342
rect 4030 4338 4034 4342
rect 4078 4338 4082 4342
rect 4118 4338 4122 4342
rect 4158 4338 4162 4342
rect 4246 4338 4250 4342
rect 4286 4338 4290 4342
rect 4318 4338 4322 4342
rect 4326 4338 4330 4342
rect 4358 4338 4362 4342
rect 4478 4338 4482 4342
rect 4518 4338 4522 4342
rect 4558 4338 4562 4342
rect 4622 4338 4626 4342
rect 4750 4338 4754 4342
rect 5118 4347 5122 4351
rect 4782 4338 4786 4342
rect 4814 4338 4818 4342
rect 4846 4338 4850 4342
rect 4854 4338 4858 4342
rect 4910 4338 4914 4342
rect 4950 4338 4954 4342
rect 4998 4338 5002 4342
rect 5030 4338 5034 4342
rect 5086 4338 5090 4342
rect 5102 4338 5106 4342
rect 3366 4328 3370 4332
rect 3966 4328 3970 4332
rect 4534 4328 4538 4332
rect 4550 4328 4554 4332
rect 5022 4328 5026 4332
rect 150 4318 154 4322
rect 174 4318 178 4322
rect 214 4318 218 4322
rect 286 4318 290 4322
rect 326 4318 330 4322
rect 430 4318 434 4322
rect 846 4318 850 4322
rect 950 4318 954 4322
rect 1006 4318 1010 4322
rect 1150 4318 1154 4322
rect 1198 4318 1202 4322
rect 1326 4318 1330 4322
rect 1446 4318 1450 4322
rect 1534 4318 1538 4322
rect 1806 4318 1810 4322
rect 1918 4318 1922 4322
rect 2022 4318 2026 4322
rect 2038 4318 2042 4322
rect 2190 4318 2194 4322
rect 2198 4318 2202 4322
rect 2430 4318 2434 4322
rect 2574 4318 2578 4322
rect 2694 4318 2698 4322
rect 2710 4318 2714 4322
rect 2870 4318 2874 4322
rect 2894 4318 2898 4322
rect 2902 4318 2906 4322
rect 3118 4318 3122 4322
rect 3190 4318 3194 4322
rect 3326 4318 3330 4322
rect 3582 4318 3586 4322
rect 3598 4318 3602 4322
rect 3638 4318 3642 4322
rect 3662 4318 3666 4322
rect 3790 4318 3794 4322
rect 3886 4318 3890 4322
rect 3958 4318 3962 4322
rect 4014 4318 4018 4322
rect 4038 4318 4042 4322
rect 4334 4318 4338 4322
rect 4494 4318 4498 4322
rect 4526 4318 4530 4322
rect 4582 4318 4586 4322
rect 4630 4318 4634 4322
rect 4822 4318 4826 4322
rect 4918 4318 4922 4322
rect 1050 4303 1054 4307
rect 1057 4303 1061 4307
rect 2074 4303 2078 4307
rect 2081 4303 2085 4307
rect 3098 4303 3102 4307
rect 3105 4303 3109 4307
rect 4114 4303 4118 4307
rect 4121 4303 4125 4307
rect 70 4288 74 4292
rect 238 4288 242 4292
rect 382 4288 386 4292
rect 598 4288 602 4292
rect 886 4288 890 4292
rect 1206 4288 1210 4292
rect 1230 4288 1234 4292
rect 1286 4288 1290 4292
rect 1438 4288 1442 4292
rect 1942 4288 1946 4292
rect 1998 4288 2002 4292
rect 2166 4288 2170 4292
rect 2302 4288 2306 4292
rect 2334 4288 2338 4292
rect 2654 4288 2658 4292
rect 3046 4288 3050 4292
rect 3094 4288 3098 4292
rect 3934 4288 3938 4292
rect 3974 4288 3978 4292
rect 4198 4288 4202 4292
rect 4214 4288 4218 4292
rect 4702 4288 4706 4292
rect 22 4278 26 4282
rect 414 4278 418 4282
rect 694 4278 698 4282
rect 750 4278 754 4282
rect 918 4278 922 4282
rect 974 4278 978 4282
rect 1094 4278 1098 4282
rect 1222 4278 1226 4282
rect 1342 4278 1346 4282
rect 1446 4278 1450 4282
rect 1766 4278 1770 4282
rect 1798 4278 1802 4282
rect 46 4268 50 4272
rect 126 4268 130 4272
rect 142 4268 146 4272
rect 262 4268 266 4272
rect 358 4268 362 4272
rect 374 4268 378 4272
rect 454 4268 458 4272
rect 542 4268 546 4272
rect 590 4268 594 4272
rect 662 4268 666 4272
rect 726 4268 730 4272
rect 734 4268 738 4272
rect 782 4268 786 4272
rect 798 4268 802 4272
rect 814 4268 818 4272
rect 878 4268 882 4272
rect 990 4268 994 4272
rect 1046 4268 1050 4272
rect 1166 4268 1170 4272
rect 1190 4268 1194 4272
rect 1254 4268 1258 4272
rect 1262 4268 1266 4272
rect 1302 4268 1306 4272
rect 1382 4268 1386 4272
rect 1574 4268 1578 4272
rect 1638 4268 1642 4272
rect 1694 4268 1698 4272
rect 1830 4268 1834 4272
rect 1846 4268 1850 4272
rect 1990 4268 1994 4272
rect 2014 4278 2018 4282
rect 2214 4278 2218 4282
rect 2438 4278 2442 4282
rect 2590 4278 2594 4282
rect 2686 4278 2690 4282
rect 2750 4278 2754 4282
rect 2934 4278 2938 4282
rect 3078 4278 3082 4282
rect 3318 4278 3322 4282
rect 3510 4278 3514 4282
rect 3718 4278 3722 4282
rect 3990 4278 3994 4282
rect 4286 4278 4290 4282
rect 4302 4278 4306 4282
rect 2062 4268 2066 4272
rect 2150 4268 2154 4272
rect 2198 4268 2202 4272
rect 2222 4268 2226 4272
rect 2270 4268 2274 4272
rect 2278 4268 2282 4272
rect 2310 4268 2314 4272
rect 2662 4268 2666 4272
rect 2710 4268 2714 4272
rect 2966 4268 2970 4272
rect 3038 4268 3042 4272
rect 3086 4268 3090 4272
rect 3150 4268 3154 4272
rect 3246 4268 3250 4272
rect 3302 4268 3306 4272
rect 3342 4268 3346 4272
rect 3374 4268 3378 4272
rect 3414 4268 3418 4272
rect 3478 4268 3482 4272
rect 6 4258 10 4262
rect 54 4258 58 4262
rect 174 4258 178 4262
rect 246 4258 250 4262
rect 286 4258 290 4262
rect 366 4258 370 4262
rect 398 4258 402 4262
rect 422 4258 426 4262
rect 430 4258 434 4262
rect 438 4258 442 4262
rect 550 4258 554 4262
rect 654 4258 658 4262
rect 710 4258 714 4262
rect 742 4258 746 4262
rect 806 4258 810 4262
rect 822 4258 826 4262
rect 830 4258 834 4262
rect 854 4258 858 4262
rect 870 4258 874 4262
rect 902 4258 906 4262
rect 926 4258 930 4262
rect 934 4258 938 4262
rect 958 4258 962 4262
rect 998 4258 1002 4262
rect 1054 4258 1058 4262
rect 1094 4259 1098 4263
rect 1166 4258 1170 4262
rect 1206 4258 1210 4262
rect 1246 4258 1250 4262
rect 1294 4258 1298 4262
rect 1326 4258 1330 4262
rect 1382 4258 1386 4262
rect 1494 4258 1498 4262
rect 1518 4258 1522 4262
rect 1582 4258 1586 4262
rect 1590 4258 1594 4262
rect 1646 4258 1650 4262
rect 1686 4258 1690 4262
rect 1758 4258 1762 4262
rect 1878 4258 1882 4262
rect 1958 4258 1962 4262
rect 1974 4258 1978 4262
rect 1982 4258 1986 4262
rect 2038 4258 2042 4262
rect 2086 4258 2090 4262
rect 2190 4258 2194 4262
rect 2238 4258 2242 4262
rect 2270 4258 2274 4262
rect 2286 4258 2290 4262
rect 2318 4258 2322 4262
rect 2342 4258 2346 4262
rect 2350 4258 2354 4262
rect 2374 4258 2378 4262
rect 2390 4258 2394 4262
rect 2398 4258 2402 4262
rect 2422 4258 2426 4262
rect 2518 4259 2522 4263
rect 2598 4258 2602 4262
rect 2702 4258 2706 4262
rect 2734 4258 2738 4262
rect 2782 4259 2786 4263
rect 2814 4258 2818 4262
rect 2854 4258 2858 4262
rect 2862 4258 2866 4262
rect 2886 4258 2890 4262
rect 2894 4258 2898 4262
rect 2918 4258 2922 4262
rect 2958 4258 2962 4262
rect 2990 4258 2994 4262
rect 3014 4258 3018 4262
rect 3022 4258 3026 4262
rect 3030 4258 3034 4262
rect 3062 4258 3066 4262
rect 3142 4258 3146 4262
rect 3158 4258 3162 4262
rect 3166 4258 3170 4262
rect 3190 4258 3194 4262
rect 3238 4258 3242 4262
rect 3334 4258 3338 4262
rect 3350 4258 3354 4262
rect 3366 4258 3370 4262
rect 3406 4259 3410 4263
rect 3606 4268 3610 4272
rect 3622 4268 3626 4272
rect 3702 4268 3706 4272
rect 3750 4268 3754 4272
rect 3774 4268 3778 4272
rect 3782 4268 3786 4272
rect 3486 4258 3490 4262
rect 3510 4258 3514 4262
rect 3534 4258 3538 4262
rect 3558 4258 3562 4262
rect 3566 4258 3570 4262
rect 3574 4258 3578 4262
rect 3590 4258 3594 4262
rect 3630 4258 3634 4262
rect 3638 4258 3642 4262
rect 3718 4259 3722 4263
rect 3838 4268 3842 4272
rect 3870 4268 3874 4272
rect 3878 4268 3882 4272
rect 3910 4268 3914 4272
rect 3918 4268 3922 4272
rect 3942 4268 3946 4272
rect 3958 4268 3962 4272
rect 4030 4268 4034 4272
rect 4062 4268 4066 4272
rect 4182 4268 4186 4272
rect 4222 4268 4226 4272
rect 4254 4268 4258 4272
rect 4262 4268 4266 4272
rect 4670 4278 4674 4282
rect 4830 4278 4834 4282
rect 4326 4268 4330 4272
rect 4374 4268 4378 4272
rect 4454 4268 4458 4272
rect 4486 4268 4490 4272
rect 4566 4268 4570 4272
rect 4678 4268 4682 4272
rect 4782 4268 4786 4272
rect 4798 4268 4802 4272
rect 4854 4268 4858 4272
rect 4942 4268 4946 4272
rect 4958 4268 4962 4272
rect 5014 4268 5018 4272
rect 5102 4268 5106 4272
rect 5118 4268 5122 4272
rect 3766 4258 3770 4262
rect 3790 4258 3794 4262
rect 3814 4258 3818 4262
rect 3830 4258 3834 4262
rect 3846 4258 3850 4262
rect 4022 4258 4026 4262
rect 4062 4258 4066 4262
rect 4070 4258 4074 4262
rect 4078 4258 4082 4262
rect 4102 4258 4106 4262
rect 4134 4258 4138 4262
rect 4142 4258 4146 4262
rect 4166 4258 4170 4262
rect 4230 4258 4234 4262
rect 4246 4258 4250 4262
rect 4286 4258 4290 4262
rect 4318 4258 4322 4262
rect 4334 4258 4338 4262
rect 4366 4259 4370 4263
rect 4478 4258 4482 4262
rect 4494 4258 4498 4262
rect 4510 4258 4514 4262
rect 4566 4258 4570 4262
rect 4630 4258 4634 4262
rect 4694 4258 4698 4262
rect 4766 4259 4770 4263
rect 4806 4258 4810 4262
rect 4846 4258 4850 4262
rect 4918 4258 4922 4262
rect 4966 4258 4970 4262
rect 5006 4258 5010 4262
rect 5070 4258 5074 4262
rect 446 4248 450 4252
rect 574 4248 578 4252
rect 766 4248 770 4252
rect 1038 4248 1042 4252
rect 1182 4248 1186 4252
rect 1286 4248 1290 4252
rect 1318 4248 1322 4252
rect 1606 4248 1610 4252
rect 1686 4248 1690 4252
rect 1814 4248 1818 4252
rect 1974 4248 1978 4252
rect 2166 4248 2170 4252
rect 2174 4248 2178 4252
rect 2238 4248 2242 4252
rect 2246 4248 2250 4252
rect 2302 4248 2306 4252
rect 2334 4248 2338 4252
rect 2678 4248 2682 4252
rect 2726 4248 2730 4252
rect 2918 4248 2922 4252
rect 2974 4248 2978 4252
rect 3102 4248 3106 4252
rect 3118 4248 3122 4252
rect 3142 4248 3146 4252
rect 3318 4248 3322 4252
rect 3350 4248 3354 4252
rect 3502 4248 3506 4252
rect 3574 4248 3578 4252
rect 3646 4248 3650 4252
rect 3750 4248 3754 4252
rect 3806 4248 3810 4252
rect 3814 4248 3818 4252
rect 3902 4248 3906 4252
rect 3934 4248 3938 4252
rect 3958 4248 3962 4252
rect 3982 4248 3986 4252
rect 4006 4248 4010 4252
rect 4038 4248 4042 4252
rect 4198 4248 4202 4252
rect 4206 4248 4210 4252
rect 4230 4248 4234 4252
rect 4278 4248 4282 4252
rect 4510 4248 4514 4252
rect 4614 4248 4618 4252
rect 4678 4248 4682 4252
rect 4822 4248 4826 4252
rect 4982 4248 4986 4252
rect 1014 4238 1018 4242
rect 1158 4238 1162 4242
rect 1222 4238 1226 4242
rect 1422 4238 1426 4242
rect 1550 4238 1554 4242
rect 1662 4238 1666 4242
rect 3878 4238 3882 4242
rect 4438 4238 4442 4242
rect 4878 4238 4882 4242
rect 5006 4238 5010 4242
rect 5022 4238 5026 4242
rect 1702 4228 1706 4232
rect 2846 4228 2850 4232
rect 30 4218 34 4222
rect 222 4218 226 4222
rect 510 4218 514 4222
rect 550 4218 554 4222
rect 758 4218 762 4222
rect 846 4218 850 4222
rect 950 4218 954 4222
rect 982 4218 986 4222
rect 1454 4218 1458 4222
rect 1806 4218 1810 4222
rect 1822 4218 1826 4222
rect 2142 4218 2146 4222
rect 2158 4218 2162 4222
rect 2190 4218 2194 4222
rect 2206 4218 2210 4222
rect 2262 4218 2266 4222
rect 2358 4218 2362 4222
rect 2414 4218 2418 4222
rect 2446 4218 2450 4222
rect 2454 4218 2458 4222
rect 2670 4218 2674 4222
rect 2694 4218 2698 4222
rect 2870 4218 2874 4222
rect 2998 4218 3002 4222
rect 3174 4218 3178 4222
rect 3470 4218 3474 4222
rect 3518 4218 3522 4222
rect 3550 4218 3554 4222
rect 3654 4218 3658 4222
rect 3790 4218 3794 4222
rect 3950 4218 3954 4222
rect 3998 4218 4002 4222
rect 4022 4218 4026 4222
rect 4054 4218 4058 4222
rect 4094 4218 4098 4222
rect 4150 4218 4154 4222
rect 4430 4218 4434 4222
rect 4518 4218 4522 4222
rect 4630 4218 4634 4222
rect 4862 4218 4866 4222
rect 5174 4218 5178 4222
rect 538 4203 542 4207
rect 545 4203 549 4207
rect 1562 4203 1566 4207
rect 1569 4203 1573 4207
rect 2586 4203 2590 4207
rect 2593 4203 2597 4207
rect 3610 4203 3614 4207
rect 3617 4203 3621 4207
rect 4634 4203 4638 4207
rect 4641 4203 4645 4207
rect 94 4188 98 4192
rect 782 4188 786 4192
rect 934 4188 938 4192
rect 1166 4188 1170 4192
rect 1358 4188 1362 4192
rect 1374 4188 1378 4192
rect 2342 4188 2346 4192
rect 2726 4188 2730 4192
rect 2782 4188 2786 4192
rect 2838 4188 2842 4192
rect 3054 4188 3058 4192
rect 3478 4188 3482 4192
rect 3526 4188 3530 4192
rect 3854 4188 3858 4192
rect 4494 4188 4498 4192
rect 1326 4178 1330 4182
rect 2310 4178 2314 4182
rect 4718 4178 4722 4182
rect 734 4168 738 4172
rect 1222 4168 1226 4172
rect 1878 4168 1882 4172
rect 1918 4168 1922 4172
rect 1966 4168 1970 4172
rect 2006 4168 2010 4172
rect 2022 4168 2026 4172
rect 2358 4168 2362 4172
rect 3286 4168 3290 4172
rect 3430 4168 3434 4172
rect 3558 4168 3562 4172
rect 3638 4168 3642 4172
rect 3782 4168 3786 4172
rect 3966 4168 3970 4172
rect 3998 4168 4002 4172
rect 4086 4168 4090 4172
rect 4206 4168 4210 4172
rect 4462 4168 4466 4172
rect 4574 4168 4578 4172
rect 5054 4168 5058 4172
rect 5182 4168 5186 4172
rect 30 4147 34 4151
rect 62 4148 66 4152
rect 134 4148 138 4152
rect 214 4148 218 4152
rect 222 4148 226 4152
rect 246 4158 250 4162
rect 270 4158 274 4162
rect 302 4148 306 4152
rect 326 4158 330 4162
rect 350 4158 354 4162
rect 382 4158 386 4162
rect 422 4158 426 4162
rect 518 4158 522 4162
rect 742 4158 746 4162
rect 366 4148 370 4152
rect 422 4148 426 4152
rect 438 4148 442 4152
rect 470 4148 474 4152
rect 478 4148 482 4152
rect 494 4148 498 4152
rect 566 4148 570 4152
rect 590 4148 594 4152
rect 670 4148 674 4152
rect 750 4148 754 4152
rect 758 4148 762 4152
rect 782 4148 786 4152
rect 806 4158 810 4162
rect 894 4158 898 4162
rect 958 4158 962 4162
rect 1006 4158 1010 4162
rect 1182 4158 1186 4162
rect 1198 4158 1202 4162
rect 1206 4158 1210 4162
rect 1278 4158 1282 4162
rect 830 4148 834 4152
rect 838 4148 842 4152
rect 878 4148 882 4152
rect 910 4148 914 4152
rect 950 4148 954 4152
rect 990 4148 994 4152
rect 1014 4148 1018 4152
rect 1022 4148 1026 4152
rect 1046 4148 1050 4152
rect 1110 4148 1114 4152
rect 1182 4148 1186 4152
rect 1222 4148 1226 4152
rect 1246 4148 1250 4152
rect 1406 4158 1410 4162
rect 1526 4158 1530 4162
rect 1534 4158 1538 4162
rect 1302 4148 1306 4152
rect 1342 4148 1346 4152
rect 1358 4148 1362 4152
rect 1382 4148 1386 4152
rect 1446 4148 1450 4152
rect 1558 4148 1562 4152
rect 1582 4148 1586 4152
rect 1606 4148 1610 4152
rect 1630 4158 1634 4162
rect 1710 4158 1714 4162
rect 1726 4158 1730 4162
rect 1734 4158 1738 4162
rect 1662 4148 1666 4152
rect 1686 4148 1690 4152
rect 1694 4148 1698 4152
rect 1710 4148 1714 4152
rect 1822 4147 1826 4151
rect 1870 4148 1874 4152
rect 1910 4148 1914 4152
rect 1934 4148 1938 4152
rect 1950 4148 1954 4152
rect 1990 4158 1994 4162
rect 2110 4158 2114 4162
rect 2278 4158 2282 4162
rect 2294 4158 2298 4162
rect 2326 4158 2330 4162
rect 2366 4158 2370 4162
rect 2630 4158 2634 4162
rect 2686 4158 2690 4162
rect 1990 4148 1994 4152
rect 2062 4148 2066 4152
rect 2166 4148 2170 4152
rect 2230 4148 2234 4152
rect 2278 4148 2282 4152
rect 2310 4148 2314 4152
rect 2342 4148 2346 4152
rect 2398 4148 2402 4152
rect 2422 4148 2426 4152
rect 2430 4148 2434 4152
rect 2454 4148 2458 4152
rect 2470 4148 2474 4152
rect 2486 4148 2490 4152
rect 2534 4148 2538 4152
rect 2614 4148 2618 4152
rect 2670 4148 2674 4152
rect 2678 4148 2682 4152
rect 2702 4148 2706 4152
rect 2726 4148 2730 4152
rect 2750 4158 2754 4162
rect 2806 4158 2810 4162
rect 2862 4158 2866 4162
rect 2934 4158 2938 4162
rect 3414 4158 3418 4162
rect 3446 4158 3450 4162
rect 3566 4158 3570 4162
rect 3742 4158 3746 4162
rect 3758 4158 3762 4162
rect 3950 4158 3954 4162
rect 4190 4158 4194 4162
rect 4222 4158 4226 4162
rect 4422 4158 4426 4162
rect 2798 4148 2802 4152
rect 2854 4148 2858 4152
rect 2862 4148 2866 4152
rect 2878 4148 2882 4152
rect 2918 4148 2922 4152
rect 2998 4148 3002 4152
rect 3038 4148 3042 4152
rect 3070 4148 3074 4152
rect 3134 4148 3138 4152
rect 142 4138 146 4142
rect 230 4138 234 4142
rect 262 4138 266 4142
rect 286 4138 290 4142
rect 294 4138 298 4142
rect 318 4138 322 4142
rect 342 4138 346 4142
rect 358 4138 362 4142
rect 374 4138 378 4142
rect 398 4138 402 4142
rect 430 4138 434 4142
rect 486 4138 490 4142
rect 526 4138 530 4142
rect 662 4138 666 4142
rect 766 4138 770 4142
rect 822 4138 826 4142
rect 894 4138 898 4142
rect 918 4138 922 4142
rect 974 4138 978 4142
rect 982 4138 986 4142
rect 1086 4138 1090 4142
rect 1174 4138 1178 4142
rect 1222 4138 1226 4142
rect 1254 4138 1258 4142
rect 1262 4138 1266 4142
rect 1310 4138 1314 4142
rect 1390 4138 1394 4142
rect 1422 4138 1426 4142
rect 1510 4138 1514 4142
rect 1526 4138 1530 4142
rect 1630 4138 1634 4142
rect 1646 4138 1650 4142
rect 1702 4138 1706 4142
rect 1750 4138 1754 4142
rect 1838 4138 1842 4142
rect 1894 4138 1898 4142
rect 1942 4138 1946 4142
rect 1998 4138 2002 4142
rect 2102 4138 2106 4142
rect 2118 4138 2122 4142
rect 2134 4138 2138 4142
rect 2254 4138 2258 4142
rect 2270 4138 2274 4142
rect 2302 4138 2306 4142
rect 2334 4138 2338 4142
rect 2366 4138 2370 4142
rect 2382 4138 2386 4142
rect 2478 4138 2482 4142
rect 2574 4138 2578 4142
rect 2606 4138 2610 4142
rect 2710 4138 2714 4142
rect 2766 4138 2770 4142
rect 2822 4138 2826 4142
rect 3206 4147 3210 4151
rect 3246 4148 3250 4152
rect 3326 4148 3330 4152
rect 3398 4148 3402 4152
rect 3406 4148 3410 4152
rect 3430 4148 3434 4152
rect 3454 4148 3458 4152
rect 3502 4148 3506 4152
rect 3510 4148 3514 4152
rect 3590 4148 3594 4152
rect 3694 4148 3698 4152
rect 3742 4148 3746 4152
rect 3782 4148 3786 4152
rect 3830 4148 3834 4152
rect 3846 4148 3850 4152
rect 3894 4148 3898 4152
rect 2926 4138 2930 4142
rect 2982 4138 2986 4142
rect 3022 4138 3026 4142
rect 3062 4138 3066 4142
rect 3078 4138 3082 4142
rect 3222 4138 3226 4142
rect 3238 4138 3242 4142
rect 3270 4138 3274 4142
rect 3302 4138 3306 4142
rect 3390 4138 3394 4142
rect 3422 4138 3426 4142
rect 3494 4138 3498 4142
rect 3542 4138 3546 4142
rect 3582 4138 3586 4142
rect 3702 4138 3706 4142
rect 3734 4138 3738 4142
rect 3766 4138 3770 4142
rect 3918 4147 3922 4151
rect 3974 4148 3978 4152
rect 4126 4148 4130 4152
rect 4158 4147 4162 4151
rect 4206 4148 4210 4152
rect 4222 4148 4226 4152
rect 4238 4148 4242 4152
rect 4302 4148 4306 4152
rect 4350 4148 4354 4152
rect 4382 4148 4386 4152
rect 4510 4158 4514 4162
rect 4542 4158 4546 4162
rect 4566 4158 4570 4162
rect 4686 4158 4690 4162
rect 4910 4158 4914 4162
rect 4446 4148 4450 4152
rect 4478 4148 4482 4152
rect 4526 4148 4530 4152
rect 4630 4148 4634 4152
rect 4686 4148 4690 4152
rect 4702 4148 4706 4152
rect 4774 4148 4778 4152
rect 4814 4148 4818 4152
rect 4894 4148 4898 4152
rect 4934 4158 4938 4162
rect 5070 4158 5074 4162
rect 5078 4158 5082 4162
rect 4934 4148 4938 4152
rect 5006 4148 5010 4152
rect 5054 4148 5058 4152
rect 5118 4147 5122 4151
rect 3814 4138 3818 4142
rect 3822 4138 3826 4142
rect 3974 4138 3978 4142
rect 3982 4138 3986 4142
rect 4006 4138 4010 4142
rect 4078 4138 4082 4142
rect 4214 4138 4218 4142
rect 4246 4138 4250 4142
rect 4294 4138 4298 4142
rect 4334 4138 4338 4142
rect 4358 4138 4362 4142
rect 4374 4138 4378 4142
rect 4406 4138 4410 4142
rect 4454 4138 4458 4142
rect 4478 4138 4482 4142
rect 4486 4138 4490 4142
rect 4518 4138 4522 4142
rect 4542 4138 4546 4142
rect 4550 4138 4554 4142
rect 4654 4138 4658 4142
rect 4710 4138 4714 4142
rect 4798 4138 4802 4142
rect 4878 4138 4882 4142
rect 4886 4138 4890 4142
rect 4942 4138 4946 4142
rect 5030 4138 5034 4142
rect 5046 4138 5050 4142
rect 5102 4138 5106 4142
rect 878 4128 882 4132
rect 1318 4128 1322 4132
rect 1342 4128 1346 4132
rect 1366 4128 1370 4132
rect 1566 4128 1570 4132
rect 1854 4128 1858 4132
rect 2142 4128 2146 4132
rect 2438 4128 2442 4132
rect 2686 4128 2690 4132
rect 2902 4128 2906 4132
rect 3118 4128 3122 4132
rect 3470 4128 3474 4132
rect 3606 4128 3610 4132
rect 4398 4128 4402 4132
rect 5086 4128 5090 4132
rect 278 4118 282 4122
rect 462 4118 466 4122
rect 534 4118 538 4122
rect 846 4118 850 4122
rect 886 4118 890 4122
rect 958 4118 962 4122
rect 1006 4118 1010 4122
rect 1038 4118 1042 4122
rect 1166 4118 1170 4122
rect 1214 4118 1218 4122
rect 1286 4118 1290 4122
rect 1406 4118 1410 4122
rect 1502 4118 1506 4122
rect 1526 4118 1530 4122
rect 1670 4118 1674 4122
rect 1742 4118 1746 4122
rect 1758 4118 1762 4122
rect 2150 4118 2154 4122
rect 2414 4118 2418 4122
rect 2494 4118 2498 4122
rect 2654 4118 2658 4122
rect 2806 4118 2810 4122
rect 2942 4118 2946 4122
rect 3054 4118 3058 4122
rect 3086 4118 3090 4122
rect 3142 4118 3146 4122
rect 3262 4118 3266 4122
rect 3382 4118 3386 4122
rect 3558 4118 3562 4122
rect 3574 4118 3578 4122
rect 3774 4118 3778 4122
rect 3990 4118 3994 4122
rect 4254 4118 4258 4122
rect 4430 4118 4434 4122
rect 4462 4118 4466 4122
rect 4566 4118 4570 4122
rect 4950 4118 4954 4122
rect 1050 4103 1054 4107
rect 1057 4103 1061 4107
rect 2074 4103 2078 4107
rect 2081 4103 2085 4107
rect 3098 4103 3102 4107
rect 3105 4103 3109 4107
rect 4114 4103 4118 4107
rect 4121 4103 4125 4107
rect 94 4088 98 4092
rect 454 4088 458 4092
rect 502 4088 506 4092
rect 518 4088 522 4092
rect 622 4088 626 4092
rect 694 4088 698 4092
rect 742 4088 746 4092
rect 854 4088 858 4092
rect 1390 4088 1394 4092
rect 1534 4088 1538 4092
rect 1918 4088 1922 4092
rect 1974 4088 1978 4092
rect 2142 4088 2146 4092
rect 2182 4088 2186 4092
rect 2302 4088 2306 4092
rect 2542 4088 2546 4092
rect 2934 4088 2938 4092
rect 2974 4088 2978 4092
rect 3206 4088 3210 4092
rect 3318 4088 3322 4092
rect 3358 4088 3362 4092
rect 3398 4088 3402 4092
rect 3430 4088 3434 4092
rect 3454 4088 3458 4092
rect 3662 4088 3666 4092
rect 3694 4088 3698 4092
rect 3862 4088 3866 4092
rect 4070 4088 4074 4092
rect 4206 4088 4210 4092
rect 4334 4088 4338 4092
rect 4446 4088 4450 4092
rect 4646 4088 4650 4092
rect 4742 4088 4746 4092
rect 5078 4088 5082 4092
rect 150 4078 154 4082
rect 510 4078 514 4082
rect 630 4078 634 4082
rect 862 4078 866 4082
rect 1222 4078 1226 4082
rect 1382 4078 1386 4082
rect 1438 4078 1442 4082
rect 2150 4078 2154 4082
rect 2526 4078 2530 4082
rect 2582 4078 2586 4082
rect 2902 4078 2906 4082
rect 3046 4078 3050 4082
rect 110 4068 114 4072
rect 126 4068 130 4072
rect 166 4068 170 4072
rect 318 4068 322 4072
rect 446 4068 450 4072
rect 470 4068 474 4072
rect 494 4068 498 4072
rect 534 4068 538 4072
rect 590 4068 594 4072
rect 678 4068 682 4072
rect 734 4068 738 4072
rect 758 4068 762 4072
rect 774 4068 778 4072
rect 886 4068 890 4072
rect 894 4068 898 4072
rect 910 4068 914 4072
rect 1054 4068 1058 4072
rect 1086 4068 1090 4072
rect 1150 4068 1154 4072
rect 1190 4068 1194 4072
rect 1310 4068 1314 4072
rect 1374 4068 1378 4072
rect 1406 4068 1410 4072
rect 1494 4068 1498 4072
rect 1550 4068 1554 4072
rect 1630 4068 1634 4072
rect 1766 4068 1770 4072
rect 1790 4068 1794 4072
rect 1814 4068 1818 4072
rect 1822 4068 1826 4072
rect 1854 4068 1858 4072
rect 1934 4068 1938 4072
rect 1982 4068 1986 4072
rect 1990 4068 1994 4072
rect 2102 4068 2106 4072
rect 2118 4068 2122 4072
rect 2158 4068 2162 4072
rect 2206 4068 2210 4072
rect 2214 4068 2218 4072
rect 2246 4068 2250 4072
rect 2270 4068 2274 4072
rect 2318 4068 2322 4072
rect 2326 4068 2330 4072
rect 2350 4068 2354 4072
rect 2518 4068 2522 4072
rect 2566 4068 2570 4072
rect 2614 4068 2618 4072
rect 2638 4068 2642 4072
rect 2646 4068 2650 4072
rect 2758 4068 2762 4072
rect 2774 4068 2778 4072
rect 2830 4068 2834 4072
rect 2950 4068 2954 4072
rect 2958 4068 2962 4072
rect 3198 4078 3202 4082
rect 3246 4078 3250 4082
rect 3278 4078 3282 4082
rect 3390 4078 3394 4082
rect 3446 4078 3450 4082
rect 3886 4078 3890 4082
rect 4014 4078 4018 4082
rect 4238 4078 4242 4082
rect 4246 4078 4250 4082
rect 4318 4078 4322 4082
rect 4486 4078 4490 4082
rect 4598 4078 4602 4082
rect 4750 4078 4754 4082
rect 3062 4068 3066 4072
rect 3070 4068 3074 4072
rect 3182 4068 3186 4072
rect 3310 4068 3314 4072
rect 3334 4068 3338 4072
rect 3382 4068 3386 4072
rect 3462 4068 3466 4072
rect 3494 4068 3498 4072
rect 3526 4068 3530 4072
rect 3534 4068 3538 4072
rect 3566 4068 3570 4072
rect 3638 4068 3642 4072
rect 3734 4068 3738 4072
rect 3766 4068 3770 4072
rect 3798 4068 3802 4072
rect 3854 4068 3858 4072
rect 3974 4068 3978 4072
rect 4006 4068 4010 4072
rect 4054 4068 4058 4072
rect 4062 4068 4066 4072
rect 4182 4068 4186 4072
rect 4230 4068 4234 4072
rect 4254 4068 4258 4072
rect 4310 4068 4314 4072
rect 4414 4068 4418 4072
rect 4430 4068 4434 4072
rect 4478 4068 4482 4072
rect 4582 4068 4586 4072
rect 4654 4068 4658 4072
rect 4734 4068 4738 4072
rect 4758 4068 4762 4072
rect 4798 4068 4802 4072
rect 4886 4068 4890 4072
rect 4982 4068 4986 4072
rect 4998 4068 5002 4072
rect 5062 4068 5066 4072
rect 5086 4068 5090 4072
rect 5174 4068 5178 4072
rect 38 4058 42 4062
rect 62 4058 66 4062
rect 102 4058 106 4062
rect 134 4058 138 4062
rect 190 4058 194 4062
rect 270 4058 274 4062
rect 326 4058 330 4062
rect 334 4058 338 4062
rect 358 4058 362 4062
rect 374 4058 378 4062
rect 382 4058 386 4062
rect 438 4058 442 4062
rect 582 4058 586 4062
rect 590 4058 594 4062
rect 638 4058 642 4062
rect 646 4058 650 4062
rect 670 4058 674 4062
rect 710 4058 714 4062
rect 798 4058 802 4062
rect 886 4058 890 4062
rect 918 4058 922 4062
rect 926 4058 930 4062
rect 950 4058 954 4062
rect 966 4058 970 4062
rect 998 4058 1002 4062
rect 1006 4058 1010 4062
rect 1062 4058 1066 4062
rect 1126 4058 1130 4062
rect 1142 4058 1146 4062
rect 1150 4058 1154 4062
rect 1190 4058 1194 4062
rect 1254 4058 1258 4062
rect 1262 4058 1266 4062
rect 1294 4059 1298 4063
rect 1398 4058 1402 4062
rect 1414 4058 1418 4062
rect 1454 4058 1458 4062
rect 1462 4058 1466 4062
rect 1486 4058 1490 4062
rect 1502 4058 1506 4062
rect 1518 4058 1522 4062
rect 1566 4058 1570 4062
rect 1606 4058 1610 4062
rect 1614 4058 1618 4062
rect 1654 4058 1658 4062
rect 1726 4058 1730 4062
rect 1750 4058 1754 4062
rect 1758 4058 1762 4062
rect 1774 4058 1778 4062
rect 1830 4058 1834 4062
rect 1886 4058 1890 4062
rect 1894 4058 1898 4062
rect 1902 4058 1906 4062
rect 1942 4058 1946 4062
rect 1958 4058 1962 4062
rect 1998 4058 2002 4062
rect 2014 4058 2018 4062
rect 2078 4058 2082 4062
rect 2134 4058 2138 4062
rect 2166 4058 2170 4062
rect 2222 4058 2226 4062
rect 2294 4058 2298 4062
rect 2334 4058 2338 4062
rect 2358 4058 2362 4062
rect 2366 4058 2370 4062
rect 2390 4058 2394 4062
rect 2414 4058 2418 4062
rect 2438 4058 2442 4062
rect 2446 4058 2450 4062
rect 2558 4058 2562 4062
rect 2606 4058 2610 4062
rect 2646 4058 2650 4062
rect 2742 4059 2746 4063
rect 2774 4058 2778 4062
rect 2822 4058 2826 4062
rect 2894 4058 2898 4062
rect 2990 4058 2994 4062
rect 3014 4058 3018 4062
rect 3022 4058 3026 4062
rect 3030 4058 3034 4062
rect 3078 4058 3082 4062
rect 3158 4058 3162 4062
rect 3270 4058 3274 4062
rect 3342 4058 3346 4062
rect 3406 4058 3410 4062
rect 3414 4058 3418 4062
rect 3470 4058 3474 4062
rect 3518 4058 3522 4062
rect 3574 4058 3578 4062
rect 3630 4058 3634 4062
rect 3646 4058 3650 4062
rect 3670 4058 3674 4062
rect 3710 4058 3714 4062
rect 3758 4058 3762 4062
rect 3790 4058 3794 4062
rect 3806 4058 3810 4062
rect 3814 4058 3818 4062
rect 3838 4058 3842 4062
rect 3886 4058 3890 4062
rect 3910 4058 3914 4062
rect 3934 4058 3938 4062
rect 3942 4058 3946 4062
rect 3950 4058 3954 4062
rect 3998 4058 4002 4062
rect 4038 4058 4042 4062
rect 4046 4058 4050 4062
rect 4086 4058 4090 4062
rect 4094 4058 4098 4062
rect 4118 4058 4122 4062
rect 4126 4058 4130 4062
rect 4166 4058 4170 4062
rect 4190 4058 4194 4062
rect 4262 4058 4266 4062
rect 4302 4058 4306 4062
rect 4390 4058 4394 4062
rect 4446 4058 4450 4062
rect 4470 4058 4474 4062
rect 4558 4058 4562 4062
rect 4614 4058 4618 4062
rect 4662 4058 4666 4062
rect 4766 4058 4770 4062
rect 4782 4058 4786 4062
rect 4862 4058 4866 4062
rect 4958 4058 4962 4062
rect 5158 4059 5162 4063
rect 278 4048 282 4052
rect 302 4048 306 4052
rect 422 4048 426 4052
rect 454 4048 458 4052
rect 478 4048 482 4052
rect 518 4048 522 4052
rect 534 4048 538 4052
rect 574 4048 578 4052
rect 614 4048 618 4052
rect 718 4048 722 4052
rect 742 4048 746 4052
rect 862 4048 866 4052
rect 1126 4048 1130 4052
rect 1214 4048 1218 4052
rect 1238 4048 1242 4052
rect 1430 4048 1434 4052
rect 1526 4048 1530 4052
rect 1534 4048 1538 4052
rect 1798 4048 1802 4052
rect 1846 4048 1850 4052
rect 1966 4048 1970 4052
rect 2014 4048 2018 4052
rect 2190 4048 2194 4052
rect 2262 4048 2266 4052
rect 2302 4048 2306 4052
rect 2350 4048 2354 4052
rect 2542 4048 2546 4052
rect 2622 4048 2626 4052
rect 2670 4048 2674 4052
rect 2822 4048 2826 4052
rect 2934 4048 2938 4052
rect 2974 4048 2978 4052
rect 3326 4048 3330 4052
rect 3366 4048 3370 4052
rect 3478 4048 3482 4052
rect 3558 4048 3562 4052
rect 3590 4048 3594 4052
rect 3742 4048 3746 4052
rect 3774 4048 3778 4052
rect 3982 4048 3986 4052
rect 4030 4048 4034 4052
rect 4078 4048 4082 4052
rect 4150 4048 4154 4052
rect 4214 4048 4218 4052
rect 4278 4048 4282 4052
rect 4302 4048 4306 4052
rect 4446 4048 4450 4052
rect 4454 4048 4458 4052
rect 4782 4048 4786 4052
rect 5070 4048 5074 4052
rect 230 4038 234 4042
rect 494 4038 498 4042
rect 1254 4038 1258 4042
rect 1958 4038 1962 4042
rect 2582 4038 2586 4042
rect 2798 4038 2802 4042
rect 2838 4038 2842 4042
rect 3094 4038 3098 4042
rect 3790 4038 3794 4042
rect 1478 4028 1482 4032
rect 3518 4028 3522 4032
rect 3758 4028 3762 4032
rect 4502 4028 4506 4032
rect 262 4018 266 4022
rect 350 4018 354 4022
rect 398 4018 402 4022
rect 598 4018 602 4022
rect 726 4018 730 4022
rect 942 4018 946 4022
rect 990 4018 994 4022
rect 1118 4018 1122 4022
rect 1174 4018 1178 4022
rect 1198 4018 1202 4022
rect 1230 4018 1234 4022
rect 1414 4018 1418 4022
rect 1446 4018 1450 4022
rect 1598 4018 1602 4022
rect 1710 4018 1714 4022
rect 1742 4018 1746 4022
rect 2022 4018 2026 4022
rect 2222 4018 2226 4022
rect 2374 4018 2378 4022
rect 2422 4018 2426 4022
rect 2462 4018 2466 4022
rect 2534 4018 2538 4022
rect 2630 4018 2634 4022
rect 2654 4018 2658 4022
rect 2678 4018 2682 4022
rect 2998 4018 3002 4022
rect 3214 4018 3218 4022
rect 3542 4018 3546 4022
rect 3630 4018 3634 4022
rect 3894 4018 3898 4022
rect 3926 4018 3930 4022
rect 3998 4018 4002 4022
rect 4022 4018 4026 4022
rect 4102 4018 4106 4022
rect 4326 4018 4330 4022
rect 4494 4018 4498 4022
rect 4678 4018 4682 4022
rect 4902 4018 4906 4022
rect 5006 4018 5010 4022
rect 5094 4018 5098 4022
rect 538 4003 542 4007
rect 545 4003 549 4007
rect 1562 4003 1566 4007
rect 1569 4003 1573 4007
rect 2586 4003 2590 4007
rect 2593 4003 2597 4007
rect 3610 4003 3614 4007
rect 3617 4003 3621 4007
rect 4634 4003 4638 4007
rect 4641 4003 4645 4007
rect 342 3988 346 3992
rect 606 3988 610 3992
rect 622 3988 626 3992
rect 1022 3988 1026 3992
rect 1142 3988 1146 3992
rect 1254 3988 1258 3992
rect 1278 3988 1282 3992
rect 1310 3988 1314 3992
rect 1654 3988 1658 3992
rect 1870 3988 1874 3992
rect 2326 3988 2330 3992
rect 2534 3988 2538 3992
rect 2758 3988 2762 3992
rect 2982 3988 2986 3992
rect 3726 3988 3730 3992
rect 4182 3988 4186 3992
rect 4270 3988 4274 3992
rect 4398 3988 4402 3992
rect 4750 3988 4754 3992
rect 4774 3988 4778 3992
rect 4926 3988 4930 3992
rect 5110 3988 5114 3992
rect 1534 3978 1538 3982
rect 3854 3978 3858 3982
rect 94 3968 98 3972
rect 838 3968 842 3972
rect 878 3968 882 3972
rect 982 3968 986 3972
rect 1094 3968 1098 3972
rect 1174 3968 1178 3972
rect 1606 3968 1610 3972
rect 1686 3968 1690 3972
rect 1710 3968 1714 3972
rect 1894 3968 1898 3972
rect 2022 3968 2026 3972
rect 2086 3968 2090 3972
rect 2358 3968 2362 3972
rect 2726 3968 2730 3972
rect 2782 3968 2786 3972
rect 2830 3968 2834 3972
rect 2870 3968 2874 3972
rect 3062 3968 3066 3972
rect 3374 3968 3378 3972
rect 4574 3968 4578 3972
rect 4670 3968 4674 3972
rect 4734 3968 4738 3972
rect 4878 3968 4882 3972
rect 4966 3968 4970 3972
rect 310 3958 314 3962
rect 358 3958 362 3962
rect 374 3958 378 3962
rect 382 3958 386 3962
rect 406 3958 410 3962
rect 38 3948 42 3952
rect 62 3948 66 3952
rect 102 3948 106 3952
rect 134 3948 138 3952
rect 158 3948 162 3952
rect 190 3948 194 3952
rect 246 3948 250 3952
rect 358 3948 362 3952
rect 438 3948 442 3952
rect 462 3958 466 3962
rect 614 3958 618 3962
rect 718 3958 722 3962
rect 542 3948 546 3952
rect 678 3948 682 3952
rect 734 3948 738 3952
rect 782 3948 786 3952
rect 854 3948 858 3952
rect 862 3948 866 3952
rect 1126 3958 1130 3962
rect 1158 3958 1162 3962
rect 1182 3958 1186 3962
rect 1214 3958 1218 3962
rect 1246 3958 1250 3962
rect 1542 3958 1546 3962
rect 894 3948 898 3952
rect 950 3948 954 3952
rect 1014 3948 1018 3952
rect 1038 3948 1042 3952
rect 1062 3948 1066 3952
rect 1070 3948 1074 3952
rect 1118 3948 1122 3952
rect 1142 3948 1146 3952
rect 1198 3948 1202 3952
rect 1230 3948 1234 3952
rect 1326 3948 1330 3952
rect 1366 3948 1370 3952
rect 1390 3948 1394 3952
rect 1486 3948 1490 3952
rect 1590 3948 1594 3952
rect 1670 3958 1674 3962
rect 1782 3958 1786 3962
rect 1654 3948 1658 3952
rect 1686 3948 1690 3952
rect 1726 3948 1730 3952
rect 1838 3958 1842 3962
rect 1862 3958 1866 3962
rect 1990 3958 1994 3962
rect 2278 3958 2282 3962
rect 1806 3948 1810 3952
rect 1862 3948 1866 3952
rect 1958 3947 1962 3951
rect 1998 3948 2002 3952
rect 2006 3948 2010 3952
rect 2022 3948 2026 3952
rect 2038 3948 2042 3952
rect 2134 3947 2138 3951
rect 2198 3948 2202 3952
rect 2222 3948 2226 3952
rect 2662 3958 2666 3962
rect 2702 3958 2706 3962
rect 2742 3958 2746 3962
rect 2798 3958 2802 3962
rect 2838 3958 2842 3962
rect 2886 3958 2890 3962
rect 2990 3958 2994 3962
rect 3070 3958 3074 3962
rect 3270 3958 3274 3962
rect 3406 3958 3410 3962
rect 2302 3948 2306 3952
rect 2342 3948 2346 3952
rect 2366 3948 2370 3952
rect 2374 3948 2378 3952
rect 2382 3948 2386 3952
rect 2390 3948 2394 3952
rect 2414 3948 2418 3952
rect 2462 3948 2466 3952
rect 2494 3947 2498 3951
rect 2542 3948 2546 3952
rect 2598 3948 2602 3952
rect 2630 3947 2634 3951
rect 2678 3948 2682 3952
rect 2726 3948 2730 3952
rect 2758 3948 2762 3952
rect 2782 3948 2786 3952
rect 2814 3948 2818 3952
rect 2854 3948 2858 3952
rect 2870 3948 2874 3952
rect 2918 3947 2922 3951
rect 3038 3948 3042 3952
rect 3062 3948 3066 3952
rect 3086 3948 3090 3952
rect 3166 3948 3170 3952
rect 3190 3948 3194 3952
rect 3254 3948 3258 3952
rect 3310 3948 3314 3952
rect 3342 3947 3346 3951
rect 3390 3948 3394 3952
rect 3430 3958 3434 3962
rect 3574 3958 3578 3962
rect 3486 3948 3490 3952
rect 3510 3948 3514 3952
rect 3574 3948 3578 3952
rect 3598 3958 3602 3962
rect 3846 3958 3850 3962
rect 4102 3958 4106 3962
rect 4118 3958 4122 3962
rect 4166 3958 4170 3962
rect 4174 3958 4178 3962
rect 4198 3958 4202 3962
rect 4214 3958 4218 3962
rect 4246 3958 4250 3962
rect 4302 3958 4306 3962
rect 4430 3958 4434 3962
rect 4526 3958 4530 3962
rect 3662 3947 3666 3951
rect 3790 3948 3794 3952
rect 3918 3947 3922 3951
rect 3966 3948 3970 3952
rect 3998 3948 4002 3952
rect 4054 3948 4058 3952
rect 4150 3948 4154 3952
rect 4230 3948 4234 3952
rect 4254 3948 4258 3952
rect 4262 3948 4266 3952
rect 4318 3948 4322 3952
rect 4350 3948 4354 3952
rect 4382 3948 4386 3952
rect 4390 3948 4394 3952
rect 4446 3948 4450 3952
rect 4470 3948 4474 3952
rect 4478 3948 4482 3952
rect 4486 3948 4490 3952
rect 4518 3948 4522 3952
rect 4550 3948 4554 3952
rect 4590 3958 4594 3962
rect 4686 3958 4690 3962
rect 4710 3958 4714 3962
rect 4614 3948 4618 3952
rect 4782 3958 4786 3962
rect 4910 3958 4914 3962
rect 4942 3958 4946 3962
rect 4734 3948 4738 3952
rect 4822 3948 4826 3952
rect 4894 3948 4898 3952
rect 4918 3948 4922 3952
rect 4926 3948 4930 3952
rect 5014 3947 5018 3951
rect 5054 3948 5058 3952
rect 5062 3948 5066 3952
rect 5078 3958 5082 3962
rect 5150 3958 5154 3962
rect 5094 3948 5098 3952
rect 5134 3948 5138 3952
rect 5174 3948 5178 3952
rect 110 3938 114 3942
rect 126 3938 130 3942
rect 166 3938 170 3942
rect 222 3938 226 3942
rect 326 3938 330 3942
rect 398 3938 402 3942
rect 406 3938 410 3942
rect 422 3938 426 3942
rect 430 3938 434 3942
rect 454 3938 458 3942
rect 478 3938 482 3942
rect 566 3938 570 3942
rect 598 3938 602 3942
rect 670 3938 674 3942
rect 742 3938 746 3942
rect 774 3938 778 3942
rect 846 3938 850 3942
rect 902 3938 906 3942
rect 918 3938 922 3942
rect 1078 3938 1082 3942
rect 1102 3938 1106 3942
rect 1110 3938 1114 3942
rect 1158 3938 1162 3942
rect 1174 3938 1178 3942
rect 1190 3938 1194 3942
rect 1206 3938 1210 3942
rect 1238 3938 1242 3942
rect 1262 3938 1266 3942
rect 1302 3938 1306 3942
rect 1430 3938 1434 3942
rect 1486 3938 1490 3942
rect 1558 3938 1562 3942
rect 1582 3938 1586 3942
rect 1614 3938 1618 3942
rect 1638 3938 1642 3942
rect 1646 3938 1650 3942
rect 1678 3938 1682 3942
rect 1726 3938 1730 3942
rect 1758 3938 1762 3942
rect 1766 3938 1770 3942
rect 1814 3938 1818 3942
rect 1822 3938 1826 3942
rect 1838 3938 1842 3942
rect 1974 3938 1978 3942
rect 2014 3938 2018 3942
rect 2046 3938 2050 3942
rect 2262 3938 2266 3942
rect 2278 3938 2282 3942
rect 2510 3938 2514 3942
rect 2670 3938 2674 3942
rect 2734 3938 2738 3942
rect 2766 3938 2770 3942
rect 2774 3938 2778 3942
rect 2806 3938 2810 3942
rect 2830 3938 2834 3942
rect 2854 3938 2858 3942
rect 2862 3938 2866 3942
rect 2902 3938 2906 3942
rect 3014 3938 3018 3942
rect 3046 3938 3050 3942
rect 3094 3938 3098 3942
rect 3254 3938 3258 3942
rect 3390 3938 3394 3942
rect 3398 3938 3402 3942
rect 3446 3938 3450 3942
rect 3614 3938 3618 3942
rect 3670 3938 3674 3942
rect 3782 3938 3786 3942
rect 3814 3938 3818 3942
rect 3830 3938 3834 3942
rect 3934 3938 3938 3942
rect 3990 3938 3994 3942
rect 4086 3938 4090 3942
rect 4102 3938 4106 3942
rect 4134 3938 4138 3942
rect 4190 3938 4194 3942
rect 4198 3938 4202 3942
rect 4214 3938 4218 3942
rect 4246 3938 4250 3942
rect 4326 3938 4330 3942
rect 4374 3938 4378 3942
rect 4414 3938 4418 3942
rect 4534 3938 4538 3942
rect 4558 3938 4562 3942
rect 4590 3938 4594 3942
rect 4622 3938 4626 3942
rect 4646 3938 4650 3942
rect 4670 3938 4674 3942
rect 4694 3938 4698 3942
rect 4766 3938 4770 3942
rect 4814 3938 4818 3942
rect 4886 3938 4890 3942
rect 4918 3938 4922 3942
rect 5030 3938 5034 3942
rect 5046 3938 5050 3942
rect 5102 3938 5106 3942
rect 5126 3938 5130 3942
rect 5158 3938 5162 3942
rect 5190 3938 5194 3942
rect 150 3928 154 3932
rect 206 3928 210 3932
rect 334 3928 338 3932
rect 1094 3928 1098 3932
rect 1870 3928 1874 3932
rect 1886 3928 1890 3932
rect 2318 3928 2322 3932
rect 2526 3928 2530 3932
rect 2702 3928 2706 3932
rect 3230 3928 3234 3932
rect 3950 3928 3954 3932
rect 4334 3928 4338 3932
rect 4406 3928 4410 3932
rect 4534 3928 4538 3932
rect 4758 3928 4762 3932
rect 5118 3928 5122 3932
rect 174 3918 178 3922
rect 302 3918 306 3922
rect 318 3918 322 3922
rect 390 3918 394 3922
rect 486 3918 490 3922
rect 718 3918 722 3922
rect 998 3918 1002 3922
rect 1214 3918 1218 3922
rect 1542 3918 1546 3922
rect 1710 3918 1714 3922
rect 1790 3918 1794 3922
rect 1830 3918 1834 3922
rect 1854 3918 1858 3922
rect 2070 3918 2074 3922
rect 2254 3918 2258 3922
rect 2398 3918 2402 3922
rect 2430 3918 2434 3922
rect 2566 3918 2570 3922
rect 2838 3918 2842 3922
rect 2998 3918 3002 3922
rect 3022 3918 3026 3922
rect 3054 3918 3058 3922
rect 3238 3918 3242 3922
rect 3374 3918 3378 3922
rect 3558 3918 3562 3922
rect 3734 3918 3738 3922
rect 3846 3918 3850 3922
rect 3982 3918 3986 3922
rect 4006 3918 4010 3922
rect 4166 3918 4170 3922
rect 4366 3918 4370 3922
rect 4430 3918 4434 3922
rect 4454 3918 4458 3922
rect 4502 3918 4506 3922
rect 4598 3918 4602 3922
rect 4654 3918 4658 3922
rect 4678 3918 4682 3922
rect 4950 3918 4954 3922
rect 1050 3903 1054 3907
rect 1057 3903 1061 3907
rect 2074 3903 2078 3907
rect 2081 3903 2085 3907
rect 3098 3903 3102 3907
rect 3105 3903 3109 3907
rect 4114 3903 4118 3907
rect 4121 3903 4125 3907
rect 94 3888 98 3892
rect 102 3888 106 3892
rect 430 3888 434 3892
rect 662 3888 666 3892
rect 1110 3888 1114 3892
rect 1198 3888 1202 3892
rect 1318 3888 1322 3892
rect 1366 3888 1370 3892
rect 1398 3888 1402 3892
rect 1822 3888 1826 3892
rect 1926 3888 1930 3892
rect 2142 3888 2146 3892
rect 2302 3888 2306 3892
rect 2502 3888 2506 3892
rect 2982 3888 2986 3892
rect 3078 3888 3082 3892
rect 3694 3888 3698 3892
rect 3798 3888 3802 3892
rect 3878 3888 3882 3892
rect 4134 3888 4138 3892
rect 4182 3888 4186 3892
rect 4262 3888 4266 3892
rect 4550 3888 4554 3892
rect 198 3878 202 3882
rect 438 3878 442 3882
rect 926 3878 930 3882
rect 942 3878 946 3882
rect 982 3878 986 3882
rect 1118 3878 1122 3882
rect 1126 3878 1130 3882
rect 1142 3878 1146 3882
rect 1294 3878 1298 3882
rect 1310 3878 1314 3882
rect 1454 3878 1458 3882
rect 1462 3878 1466 3882
rect 1638 3878 1642 3882
rect 1734 3878 1738 3882
rect 1870 3878 1874 3882
rect 2022 3878 2026 3882
rect 2110 3878 2114 3882
rect 2374 3878 2378 3882
rect 2414 3878 2418 3882
rect 2470 3878 2474 3882
rect 2734 3878 2738 3882
rect 2790 3878 2794 3882
rect 2838 3878 2842 3882
rect 3222 3878 3226 3882
rect 3502 3878 3506 3882
rect 182 3868 186 3872
rect 262 3868 266 3872
rect 278 3868 282 3872
rect 326 3868 330 3872
rect 366 3868 370 3872
rect 486 3868 490 3872
rect 566 3868 570 3872
rect 590 3868 594 3872
rect 838 3868 842 3872
rect 958 3868 962 3872
rect 1006 3868 1010 3872
rect 1022 3868 1026 3872
rect 1166 3868 1170 3872
rect 1182 3868 1186 3872
rect 1246 3868 1250 3872
rect 1278 3868 1282 3872
rect 1358 3868 1362 3872
rect 1390 3868 1394 3872
rect 1430 3868 1434 3872
rect 1446 3868 1450 3872
rect 1470 3868 1474 3872
rect 1486 3868 1490 3872
rect 1614 3868 1618 3872
rect 1790 3868 1794 3872
rect 1846 3868 1850 3872
rect 1870 3868 1874 3872
rect 1974 3868 1978 3872
rect 2054 3868 2058 3872
rect 2102 3868 2106 3872
rect 2150 3868 2154 3872
rect 2166 3868 2170 3872
rect 2222 3868 2226 3872
rect 2310 3868 2314 3872
rect 2326 3868 2330 3872
rect 2342 3868 2346 3872
rect 2510 3868 2514 3872
rect 2518 3868 2522 3872
rect 2758 3868 2762 3872
rect 2766 3868 2770 3872
rect 2934 3868 2938 3872
rect 2950 3868 2954 3872
rect 2966 3868 2970 3872
rect 3006 3868 3010 3872
rect 3014 3868 3018 3872
rect 3046 3868 3050 3872
rect 3070 3868 3074 3872
rect 3166 3868 3170 3872
rect 3246 3868 3250 3872
rect 3374 3868 3378 3872
rect 3382 3868 3386 3872
rect 3430 3868 3434 3872
rect 3974 3878 3978 3882
rect 4718 3878 4722 3882
rect 4990 3878 4994 3882
rect 3526 3868 3530 3872
rect 3750 3868 3754 3872
rect 3766 3868 3770 3872
rect 3822 3868 3826 3872
rect 3958 3868 3962 3872
rect 3990 3868 3994 3872
rect 4014 3868 4018 3872
rect 4142 3868 4146 3872
rect 4190 3868 4194 3872
rect 4198 3868 4202 3872
rect 4254 3868 4258 3872
rect 4478 3868 4482 3872
rect 4486 3868 4490 3872
rect 4542 3868 4546 3872
rect 4606 3868 4610 3872
rect 4614 3868 4618 3872
rect 4670 3868 4674 3872
rect 4702 3868 4706 3872
rect 4758 3868 4762 3872
rect 4814 3868 4818 3872
rect 4822 3868 4826 3872
rect 4862 3868 4866 3872
rect 4878 3868 4882 3872
rect 4966 3868 4970 3872
rect 5022 3868 5026 3872
rect 5086 3868 5090 3872
rect 38 3858 42 3862
rect 62 3858 66 3862
rect 166 3859 170 3863
rect 222 3858 226 3862
rect 302 3858 306 3862
rect 374 3858 378 3862
rect 414 3858 418 3862
rect 478 3858 482 3862
rect 598 3858 602 3862
rect 702 3858 706 3862
rect 726 3858 730 3862
rect 790 3858 794 3862
rect 814 3858 818 3862
rect 822 3858 826 3862
rect 862 3858 866 3862
rect 998 3858 1002 3862
rect 1030 3858 1034 3862
rect 1054 3858 1058 3862
rect 1062 3858 1066 3862
rect 1086 3858 1090 3862
rect 1102 3858 1106 3862
rect 1142 3858 1146 3862
rect 1166 3858 1170 3862
rect 1174 3858 1178 3862
rect 1262 3859 1266 3863
rect 1326 3858 1330 3862
rect 1350 3858 1354 3862
rect 1382 3858 1386 3862
rect 1422 3858 1426 3862
rect 1478 3858 1482 3862
rect 1502 3858 1506 3862
rect 1510 3858 1514 3862
rect 1534 3858 1538 3862
rect 1558 3858 1562 3862
rect 1598 3858 1602 3862
rect 1606 3858 1610 3862
rect 1622 3858 1626 3862
rect 1646 3858 1650 3862
rect 1654 3858 1658 3862
rect 1710 3858 1714 3862
rect 1742 3858 1746 3862
rect 1750 3858 1754 3862
rect 1774 3858 1778 3862
rect 1798 3858 1802 3862
rect 1846 3858 1850 3862
rect 1854 3858 1858 3862
rect 1878 3858 1882 3862
rect 1886 3858 1890 3862
rect 1910 3858 1914 3862
rect 1990 3859 1994 3863
rect 2046 3858 2050 3862
rect 2126 3858 2130 3862
rect 2158 3858 2162 3862
rect 2174 3858 2178 3862
rect 2198 3858 2202 3862
rect 2206 3858 2210 3862
rect 2246 3858 2250 3862
rect 2318 3858 2322 3862
rect 2342 3858 2346 3862
rect 2398 3858 2402 3862
rect 2422 3858 2426 3862
rect 2430 3858 2434 3862
rect 2462 3858 2466 3862
rect 2486 3858 2490 3862
rect 2518 3858 2522 3862
rect 2534 3858 2538 3862
rect 2558 3858 2562 3862
rect 2566 3858 2570 3862
rect 2598 3858 2602 3862
rect 2622 3858 2626 3862
rect 2630 3858 2634 3862
rect 2638 3858 2642 3862
rect 2646 3858 2650 3862
rect 2670 3858 2674 3862
rect 2694 3858 2698 3862
rect 2718 3858 2722 3862
rect 2726 3858 2730 3862
rect 2750 3858 2754 3862
rect 2814 3858 2818 3862
rect 2918 3859 2922 3863
rect 2958 3858 2962 3862
rect 2998 3858 3002 3862
rect 3014 3858 3018 3862
rect 3142 3858 3146 3862
rect 3158 3858 3162 3862
rect 3222 3858 3226 3862
rect 3254 3858 3258 3862
rect 3262 3858 3266 3862
rect 3286 3858 3290 3862
rect 3334 3858 3338 3862
rect 3342 3858 3346 3862
rect 3366 3858 3370 3862
rect 3414 3858 3418 3862
rect 3422 3858 3426 3862
rect 3438 3858 3442 3862
rect 3446 3858 3450 3862
rect 3470 3858 3474 3862
rect 3486 3858 3490 3862
rect 3510 3858 3514 3862
rect 3534 3858 3538 3862
rect 3566 3859 3570 3863
rect 3598 3858 3602 3862
rect 3638 3858 3642 3862
rect 3686 3858 3690 3862
rect 3710 3858 3714 3862
rect 3718 3858 3722 3862
rect 3726 3858 3730 3862
rect 3758 3858 3762 3862
rect 3774 3858 3778 3862
rect 3814 3858 3818 3862
rect 3838 3858 3842 3862
rect 3862 3858 3866 3862
rect 3870 3858 3874 3862
rect 3942 3859 3946 3863
rect 3990 3858 3994 3862
rect 4022 3858 4026 3862
rect 4062 3858 4066 3862
rect 4086 3858 4090 3862
rect 4150 3858 4154 3862
rect 4206 3858 4210 3862
rect 4246 3858 4250 3862
rect 4294 3858 4298 3862
rect 4318 3858 4322 3862
rect 4366 3858 4370 3862
rect 4390 3858 4394 3862
rect 4398 3858 4402 3862
rect 4414 3858 4418 3862
rect 4438 3858 4442 3862
rect 4446 3858 4450 3862
rect 4454 3858 4458 3862
rect 4470 3858 4474 3862
rect 4494 3858 4498 3862
rect 4526 3858 4530 3862
rect 4534 3858 4538 3862
rect 4630 3859 4634 3863
rect 4694 3858 4698 3862
rect 4726 3858 4730 3862
rect 4766 3858 4770 3862
rect 4806 3858 4810 3862
rect 4830 3858 4834 3862
rect 4870 3858 4874 3862
rect 4926 3858 4930 3862
rect 4934 3858 4938 3862
rect 5014 3858 5018 3862
rect 5078 3858 5082 3862
rect 5126 3858 5130 3862
rect 5150 3858 5154 3862
rect 222 3848 226 3852
rect 246 3848 250 3852
rect 390 3848 394 3852
rect 398 3848 402 3852
rect 974 3848 978 3852
rect 1334 3848 1338 3852
rect 1350 3848 1354 3852
rect 1366 3848 1370 3852
rect 1398 3848 1402 3852
rect 1446 3848 1450 3852
rect 1494 3848 1498 3852
rect 1582 3848 1586 3852
rect 1638 3848 1642 3852
rect 1694 3848 1698 3852
rect 1814 3848 1818 3852
rect 1822 3848 1826 3852
rect 2086 3848 2090 3852
rect 2334 3848 2338 3852
rect 2350 3848 2354 3852
rect 2374 3848 2378 3852
rect 2414 3848 2418 3852
rect 2734 3848 2738 3852
rect 2782 3848 2786 3852
rect 2830 3848 2834 3852
rect 2974 3848 2978 3852
rect 2982 3848 2986 3852
rect 3086 3848 3090 3852
rect 3246 3848 3250 3852
rect 3350 3848 3354 3852
rect 3398 3848 3402 3852
rect 3654 3848 3658 3852
rect 3790 3848 3794 3852
rect 4222 3848 4226 3852
rect 4246 3848 4250 3852
rect 4454 3848 4458 3852
rect 4510 3848 4514 3852
rect 4678 3848 4682 3852
rect 4782 3848 4786 3852
rect 4846 3848 4850 3852
rect 4998 3848 5002 3852
rect 5054 3848 5058 3852
rect 5078 3848 5082 3852
rect 918 3838 922 3842
rect 1190 3838 1194 3842
rect 2766 3838 2770 3842
rect 3070 3838 3074 3842
rect 3198 3838 3202 3842
rect 3230 3838 3234 3842
rect 4166 3838 4170 3842
rect 4886 3838 4890 3842
rect 206 3828 210 3832
rect 2438 3828 2442 3832
rect 4374 3828 4378 3832
rect 5094 3828 5098 3832
rect 358 3818 362 3822
rect 374 3818 378 3822
rect 414 3818 418 3822
rect 550 3818 554 3822
rect 774 3818 778 3822
rect 806 3818 810 3822
rect 934 3818 938 3822
rect 950 3818 954 3822
rect 966 3818 970 3822
rect 1078 3818 1082 3822
rect 1134 3818 1138 3822
rect 1302 3818 1306 3822
rect 1526 3818 1530 3822
rect 1662 3818 1666 3822
rect 1766 3818 1770 3822
rect 1798 3818 1802 3822
rect 1902 3818 1906 3822
rect 2030 3818 2034 3822
rect 2606 3818 2610 3822
rect 2662 3818 2666 3822
rect 2710 3818 2714 3822
rect 2814 3818 2818 3822
rect 3022 3818 3026 3822
rect 3326 3818 3330 3822
rect 3366 3818 3370 3822
rect 3462 3818 3466 3822
rect 3694 3818 3698 3822
rect 3854 3818 3858 3822
rect 4150 3818 4154 3822
rect 4422 3818 4426 3822
rect 4710 3818 4714 3822
rect 4806 3818 4810 3822
rect 4982 3818 4986 3822
rect 5014 3818 5018 3822
rect 538 3803 542 3807
rect 545 3803 549 3807
rect 1562 3803 1566 3807
rect 1569 3803 1573 3807
rect 2586 3803 2590 3807
rect 2593 3803 2597 3807
rect 3610 3803 3614 3807
rect 3617 3803 3621 3807
rect 4634 3803 4638 3807
rect 4641 3803 4645 3807
rect 334 3788 338 3792
rect 590 3788 594 3792
rect 686 3788 690 3792
rect 998 3788 1002 3792
rect 1158 3788 1162 3792
rect 1182 3788 1186 3792
rect 1702 3788 1706 3792
rect 1750 3788 1754 3792
rect 2254 3788 2258 3792
rect 2630 3788 2634 3792
rect 2654 3788 2658 3792
rect 2838 3788 2842 3792
rect 3358 3788 3362 3792
rect 3414 3788 3418 3792
rect 3702 3788 3706 3792
rect 4070 3788 4074 3792
rect 4158 3788 4162 3792
rect 4462 3788 4466 3792
rect 406 3778 410 3782
rect 2270 3778 2274 3782
rect 4998 3778 5002 3782
rect 894 3768 898 3772
rect 1366 3768 1370 3772
rect 1734 3768 1738 3772
rect 1894 3768 1898 3772
rect 2022 3768 2026 3772
rect 2390 3768 2394 3772
rect 2918 3768 2922 3772
rect 2934 3768 2938 3772
rect 3646 3768 3650 3772
rect 3750 3768 3754 3772
rect 3950 3768 3954 3772
rect 4174 3768 4178 3772
rect 4366 3768 4370 3772
rect 4622 3768 4626 3772
rect 4750 3768 4754 3772
rect 5094 3768 5098 3772
rect 342 3758 346 3762
rect 46 3748 50 3752
rect 134 3748 138 3752
rect 238 3747 242 3751
rect 310 3748 314 3752
rect 382 3748 386 3752
rect 406 3748 410 3752
rect 430 3758 434 3762
rect 654 3758 658 3762
rect 502 3748 506 3752
rect 686 3748 690 3752
rect 710 3758 714 3762
rect 742 3748 746 3752
rect 766 3748 770 3752
rect 774 3748 778 3752
rect 782 3748 786 3752
rect 830 3747 834 3751
rect 910 3748 914 3752
rect 918 3748 922 3752
rect 934 3758 938 3762
rect 958 3758 962 3762
rect 1014 3758 1018 3762
rect 974 3748 978 3752
rect 998 3748 1002 3752
rect 1030 3748 1034 3752
rect 1062 3758 1066 3762
rect 1102 3748 1106 3752
rect 1126 3758 1130 3762
rect 1294 3758 1298 3762
rect 1326 3758 1330 3762
rect 1126 3748 1130 3752
rect 1174 3748 1178 3752
rect 1238 3748 1242 3752
rect 1310 3748 1314 3752
rect 1462 3758 1466 3762
rect 1342 3748 1346 3752
rect 1350 3748 1354 3752
rect 1422 3748 1426 3752
rect 1518 3748 1522 3752
rect 1622 3748 1626 3752
rect 1646 3758 1650 3762
rect 1670 3758 1674 3762
rect 1694 3758 1698 3762
rect 1766 3758 1770 3762
rect 1750 3748 1754 3752
rect 1806 3748 1810 3752
rect 1830 3748 1834 3752
rect 1854 3748 1858 3752
rect 1862 3748 1866 3752
rect 1878 3748 1882 3752
rect 2046 3758 2050 3762
rect 2070 3758 2074 3762
rect 2166 3758 2170 3762
rect 2246 3758 2250 3762
rect 1910 3748 1914 3752
rect 1918 3748 1922 3752
rect 86 3738 90 3742
rect 246 3738 250 3742
rect 318 3738 322 3742
rect 358 3738 362 3742
rect 390 3738 394 3742
rect 398 3738 402 3742
rect 446 3738 450 3742
rect 486 3738 490 3742
rect 654 3738 658 3742
rect 670 3738 674 3742
rect 678 3738 682 3742
rect 726 3738 730 3742
rect 814 3738 818 3742
rect 902 3738 906 3742
rect 950 3738 954 3742
rect 982 3738 986 3742
rect 990 3738 994 3742
rect 1022 3738 1026 3742
rect 1038 3738 1042 3742
rect 1958 3747 1962 3751
rect 1990 3748 1994 3752
rect 2126 3748 2130 3752
rect 2206 3748 2210 3752
rect 2238 3748 2242 3752
rect 2350 3747 2354 3751
rect 2382 3748 2386 3752
rect 2414 3758 2418 3762
rect 2438 3758 2442 3762
rect 2590 3758 2594 3762
rect 2454 3748 2458 3752
rect 2518 3748 2522 3752
rect 2654 3748 2658 3752
rect 2678 3758 2682 3762
rect 3326 3758 3330 3762
rect 3374 3758 3378 3762
rect 3542 3758 3546 3762
rect 3574 3758 3578 3762
rect 3670 3758 3674 3762
rect 3686 3758 3690 3762
rect 3710 3758 3714 3762
rect 3718 3758 3722 3762
rect 3894 3758 3898 3762
rect 4102 3758 4106 3762
rect 4150 3758 4154 3762
rect 4302 3758 4306 3762
rect 2694 3748 2698 3752
rect 2710 3748 2714 3752
rect 2742 3748 2746 3752
rect 2750 3748 2754 3752
rect 2854 3748 2858 3752
rect 2862 3748 2866 3752
rect 2894 3748 2898 3752
rect 2910 3748 2914 3752
rect 2974 3748 2978 3752
rect 3134 3748 3138 3752
rect 3198 3748 3202 3752
rect 3230 3748 3234 3752
rect 3278 3747 3282 3751
rect 3382 3748 3386 3752
rect 3390 3748 3394 3752
rect 3406 3748 3410 3752
rect 3494 3747 3498 3751
rect 3558 3748 3562 3752
rect 3566 3748 3570 3752
rect 3614 3748 3618 3752
rect 3726 3748 3730 3752
rect 3734 3748 3738 3752
rect 3782 3748 3786 3752
rect 3814 3747 3818 3751
rect 3902 3748 3906 3752
rect 3982 3747 3986 3751
rect 4014 3748 4018 3752
rect 4054 3748 4058 3752
rect 4078 3748 4082 3752
rect 4126 3748 4130 3752
rect 4150 3748 4154 3752
rect 4206 3748 4210 3752
rect 4254 3748 4258 3752
rect 4262 3748 4266 3752
rect 4286 3748 4290 3752
rect 4318 3748 4322 3752
rect 4342 3748 4346 3752
rect 4702 3758 4706 3762
rect 4990 3758 4994 3762
rect 4398 3748 4402 3752
rect 4422 3748 4426 3752
rect 4430 3748 4434 3752
rect 4454 3748 4458 3752
rect 1094 3738 1098 3742
rect 1142 3738 1146 3742
rect 1246 3738 1250 3742
rect 1262 3738 1266 3742
rect 1278 3738 1282 3742
rect 1302 3738 1306 3742
rect 1358 3738 1362 3742
rect 1414 3738 1418 3742
rect 1478 3738 1482 3742
rect 1494 3738 1498 3742
rect 1630 3738 1634 3742
rect 1670 3738 1674 3742
rect 1686 3738 1690 3742
rect 1710 3738 1714 3742
rect 1766 3738 1770 3742
rect 1782 3738 1786 3742
rect 1822 3738 1826 3742
rect 1870 3738 1874 3742
rect 1926 3738 1930 3742
rect 2030 3738 2034 3742
rect 2054 3738 2058 3742
rect 2118 3738 2122 3742
rect 2214 3738 2218 3742
rect 2230 3738 2234 3742
rect 2262 3738 2266 3742
rect 2318 3738 2322 3742
rect 2366 3738 2370 3742
rect 2382 3738 2386 3742
rect 2430 3738 2434 3742
rect 2446 3738 2450 3742
rect 2462 3738 2466 3742
rect 2502 3738 2506 3742
rect 2550 3738 2554 3742
rect 2566 3738 2570 3742
rect 2590 3738 2594 3742
rect 2606 3738 2610 3742
rect 2646 3738 2650 3742
rect 2702 3738 2706 3742
rect 2758 3738 2762 3742
rect 2822 3738 2826 3742
rect 2902 3738 2906 3742
rect 2998 3738 3002 3742
rect 3014 3738 3018 3742
rect 3086 3738 3090 3742
rect 3110 3738 3114 3742
rect 3158 3738 3162 3742
rect 3206 3738 3210 3742
rect 3262 3738 3266 3742
rect 3310 3738 3314 3742
rect 3366 3738 3370 3742
rect 3398 3738 3402 3742
rect 3510 3738 3514 3742
rect 3526 3738 3530 3742
rect 3550 3738 3554 3742
rect 3630 3738 3634 3742
rect 3662 3738 3666 3742
rect 3670 3738 3674 3742
rect 3686 3738 3690 3742
rect 3742 3738 3746 3742
rect 3862 3738 3866 3742
rect 3878 3738 3882 3742
rect 3934 3738 3938 3742
rect 4086 3738 4090 3742
rect 4126 3738 4130 3742
rect 4526 3747 4530 3751
rect 4558 3748 4562 3752
rect 4566 3748 4570 3752
rect 4590 3748 4594 3752
rect 4598 3748 4602 3752
rect 4646 3748 4650 3752
rect 4694 3748 4698 3752
rect 4702 3748 4706 3752
rect 4718 3748 4722 3752
rect 4734 3748 4738 3752
rect 4750 3748 4754 3752
rect 4814 3748 4818 3752
rect 4902 3748 4906 3752
rect 4926 3748 4930 3752
rect 4966 3748 4970 3752
rect 4990 3748 4994 3752
rect 5030 3748 5034 3752
rect 5038 3748 5042 3752
rect 5126 3748 5130 3752
rect 4222 3738 4226 3742
rect 4294 3738 4298 3742
rect 4326 3738 4330 3742
rect 4334 3738 4338 3742
rect 4358 3738 4362 3742
rect 4382 3738 4386 3742
rect 4390 3738 4394 3742
rect 4438 3738 4442 3742
rect 4542 3738 4546 3742
rect 4606 3738 4610 3742
rect 4686 3738 4690 3742
rect 4726 3738 4730 3742
rect 4734 3738 4738 3742
rect 5158 3747 5162 3751
rect 4782 3738 4786 3742
rect 4966 3738 4970 3742
rect 5078 3738 5082 3742
rect 206 3728 210 3732
rect 334 3728 338 3732
rect 558 3728 562 3732
rect 798 3728 802 3732
rect 1198 3728 1202 3732
rect 1718 3728 1722 3732
rect 1958 3728 1962 3732
rect 2878 3728 2882 3732
rect 3214 3728 3218 3732
rect 3246 3728 3250 3732
rect 3422 3728 3426 3732
rect 3846 3728 3850 3732
rect 4662 3728 4666 3732
rect 4766 3728 4770 3732
rect 6 3718 10 3722
rect 302 3718 306 3722
rect 366 3718 370 3722
rect 542 3718 546 3722
rect 574 3718 578 3722
rect 662 3718 666 3722
rect 758 3718 762 3722
rect 790 3718 794 3722
rect 958 3718 962 3722
rect 1118 3718 1122 3722
rect 1134 3718 1138 3722
rect 1286 3718 1290 3722
rect 1470 3718 1474 3722
rect 1606 3718 1610 3722
rect 1670 3718 1674 3722
rect 1726 3718 1730 3722
rect 1790 3718 1794 3722
rect 1846 3718 1850 3722
rect 2038 3718 2042 3722
rect 2062 3718 2066 3722
rect 2270 3718 2274 3722
rect 2470 3718 2474 3722
rect 2582 3718 2586 3722
rect 2614 3718 2618 3722
rect 2726 3718 2730 3722
rect 3190 3718 3194 3722
rect 3430 3718 3434 3722
rect 3542 3718 3546 3722
rect 3590 3718 3594 3722
rect 3654 3718 3658 3722
rect 3686 3718 3690 3722
rect 3710 3718 3714 3722
rect 3854 3718 3858 3722
rect 3918 3718 3922 3722
rect 3950 3718 3954 3722
rect 4046 3718 4050 3722
rect 4102 3718 4106 3722
rect 4270 3718 4274 3722
rect 4630 3718 4634 3722
rect 4678 3718 4682 3722
rect 4774 3718 4778 3722
rect 4958 3718 4962 3722
rect 1050 3703 1054 3707
rect 1057 3703 1061 3707
rect 2074 3703 2078 3707
rect 2081 3703 2085 3707
rect 3098 3703 3102 3707
rect 3105 3703 3109 3707
rect 4114 3703 4118 3707
rect 4121 3703 4125 3707
rect 38 3688 42 3692
rect 238 3688 242 3692
rect 358 3688 362 3692
rect 502 3688 506 3692
rect 814 3688 818 3692
rect 830 3688 834 3692
rect 862 3688 866 3692
rect 1334 3688 1338 3692
rect 1446 3688 1450 3692
rect 1726 3688 1730 3692
rect 2398 3688 2402 3692
rect 2574 3688 2578 3692
rect 2630 3688 2634 3692
rect 3094 3688 3098 3692
rect 3390 3688 3394 3692
rect 3414 3688 3418 3692
rect 3526 3688 3530 3692
rect 3574 3688 3578 3692
rect 3606 3688 3610 3692
rect 3702 3688 3706 3692
rect 3830 3688 3834 3692
rect 3966 3688 3970 3692
rect 4278 3688 4282 3692
rect 4686 3688 4690 3692
rect 4718 3688 4722 3692
rect 4926 3688 4930 3692
rect 5038 3688 5042 3692
rect 5102 3688 5106 3692
rect 5166 3688 5170 3692
rect 6 3678 10 3682
rect 270 3678 274 3682
rect 350 3678 354 3682
rect 750 3678 754 3682
rect 822 3678 826 3682
rect 966 3678 970 3682
rect 1006 3678 1010 3682
rect 46 3668 50 3672
rect 86 3668 90 3672
rect 158 3668 162 3672
rect 174 3668 178 3672
rect 214 3668 218 3672
rect 230 3668 234 3672
rect 278 3668 282 3672
rect 390 3668 394 3672
rect 478 3668 482 3672
rect 566 3668 570 3672
rect 638 3668 642 3672
rect 686 3668 690 3672
rect 718 3668 722 3672
rect 838 3668 842 3672
rect 854 3668 858 3672
rect 1822 3678 1826 3682
rect 2022 3678 2026 3682
rect 3142 3678 3146 3682
rect 1102 3668 1106 3672
rect 1126 3668 1130 3672
rect 1166 3668 1170 3672
rect 1222 3668 1226 3672
rect 1262 3668 1266 3672
rect 1366 3668 1370 3672
rect 1414 3668 1418 3672
rect 1454 3668 1458 3672
rect 1470 3668 1474 3672
rect 1510 3668 1514 3672
rect 1518 3668 1522 3672
rect 1590 3668 1594 3672
rect 1598 3668 1602 3672
rect 1686 3668 1690 3672
rect 1934 3668 1938 3672
rect 2134 3668 2138 3672
rect 2150 3668 2154 3672
rect 2198 3668 2202 3672
rect 2270 3668 2274 3672
rect 2326 3668 2330 3672
rect 2374 3668 2378 3672
rect 2510 3668 2514 3672
rect 22 3658 26 3662
rect 54 3658 58 3662
rect 94 3658 98 3662
rect 166 3658 170 3662
rect 206 3658 210 3662
rect 222 3658 226 3662
rect 254 3658 258 3662
rect 342 3658 346 3662
rect 366 3658 370 3662
rect 406 3658 410 3662
rect 430 3658 434 3662
rect 438 3658 442 3662
rect 446 3658 450 3662
rect 478 3658 482 3662
rect 486 3658 490 3662
rect 558 3658 562 3662
rect 638 3658 642 3662
rect 646 3658 650 3662
rect 710 3658 714 3662
rect 758 3658 762 3662
rect 846 3658 850 3662
rect 878 3658 882 3662
rect 894 3658 898 3662
rect 910 3658 914 3662
rect 934 3658 938 3662
rect 942 3658 946 3662
rect 950 3658 954 3662
rect 982 3658 986 3662
rect 990 3658 994 3662
rect 1022 3658 1026 3662
rect 1030 3658 1034 3662
rect 1094 3658 1098 3662
rect 1110 3658 1114 3662
rect 1134 3658 1138 3662
rect 1150 3658 1154 3662
rect 1214 3658 1218 3662
rect 1254 3659 1258 3663
rect 1350 3658 1354 3662
rect 1390 3658 1394 3662
rect 1462 3658 1466 3662
rect 1478 3658 1482 3662
rect 1510 3658 1514 3662
rect 1526 3658 1530 3662
rect 1582 3658 1586 3662
rect 1598 3658 1602 3662
rect 1678 3658 1682 3662
rect 1742 3658 1746 3662
rect 1750 3658 1754 3662
rect 1758 3658 1762 3662
rect 1782 3658 1786 3662
rect 1790 3658 1794 3662
rect 1830 3658 1834 3662
rect 1838 3658 1842 3662
rect 1846 3658 1850 3662
rect 1854 3658 1858 3662
rect 1886 3658 1890 3662
rect 1894 3658 1898 3662
rect 1902 3658 1906 3662
rect 1926 3658 1930 3662
rect 1942 3658 1946 3662
rect 1950 3658 1954 3662
rect 1974 3658 1978 3662
rect 1982 3658 1986 3662
rect 2006 3658 2010 3662
rect 2118 3659 2122 3663
rect 2566 3668 2570 3672
rect 2614 3668 2618 3672
rect 2662 3668 2666 3672
rect 2734 3668 2738 3672
rect 2790 3668 2794 3672
rect 2822 3668 2826 3672
rect 2894 3668 2898 3672
rect 2902 3668 2906 3672
rect 2958 3668 2962 3672
rect 2998 3668 3002 3672
rect 3086 3668 3090 3672
rect 3158 3668 3162 3672
rect 3246 3668 3250 3672
rect 3278 3668 3282 3672
rect 3310 3668 3314 3672
rect 3406 3668 3410 3672
rect 3430 3678 3434 3682
rect 3566 3678 3570 3682
rect 3798 3678 3802 3682
rect 3918 3678 3922 3682
rect 4222 3678 4226 3682
rect 4750 3678 4754 3682
rect 4886 3678 4890 3682
rect 3502 3668 3506 3672
rect 3558 3668 3562 3672
rect 3638 3668 3642 3672
rect 3694 3668 3698 3672
rect 3782 3668 3786 3672
rect 3838 3668 3842 3672
rect 3846 3668 3850 3672
rect 3918 3668 3922 3672
rect 3942 3668 3946 3672
rect 3998 3668 4002 3672
rect 4078 3668 4082 3672
rect 4134 3668 4138 3672
rect 4182 3668 4186 3672
rect 4198 3668 4202 3672
rect 4262 3668 4266 3672
rect 4358 3668 4362 3672
rect 4454 3668 4458 3672
rect 4606 3668 4610 3672
rect 4622 3668 4626 3672
rect 4654 3668 4658 3672
rect 4710 3668 4714 3672
rect 4798 3668 4802 3672
rect 4814 3668 4818 3672
rect 4870 3668 4874 3672
rect 4902 3668 4906 3672
rect 4910 3668 4914 3672
rect 5006 3668 5010 3672
rect 5030 3668 5034 3672
rect 5054 3678 5058 3682
rect 5134 3678 5138 3682
rect 5078 3668 5082 3672
rect 5110 3668 5114 3672
rect 5174 3668 5178 3672
rect 2158 3658 2162 3662
rect 2166 3658 2170 3662
rect 2286 3658 2290 3662
rect 2310 3658 2314 3662
rect 2318 3658 2322 3662
rect 2334 3658 2338 3662
rect 2358 3658 2362 3662
rect 2366 3658 2370 3662
rect 2382 3658 2386 3662
rect 2438 3658 2442 3662
rect 2462 3658 2466 3662
rect 2518 3658 2522 3662
rect 2534 3658 2538 3662
rect 2542 3658 2546 3662
rect 2550 3658 2554 3662
rect 2606 3658 2610 3662
rect 2646 3658 2650 3662
rect 2718 3658 2722 3662
rect 2782 3658 2786 3662
rect 2798 3658 2802 3662
rect 2814 3658 2818 3662
rect 2902 3658 2906 3662
rect 2950 3658 2954 3662
rect 2990 3659 2994 3663
rect 3062 3658 3066 3662
rect 3078 3658 3082 3662
rect 3126 3658 3130 3662
rect 3182 3658 3186 3662
rect 3254 3658 3258 3662
rect 3262 3658 3266 3662
rect 3334 3658 3338 3662
rect 3398 3658 3402 3662
rect 3446 3658 3450 3662
rect 3454 3658 3458 3662
rect 3462 3658 3466 3662
rect 3486 3658 3490 3662
rect 3510 3658 3514 3662
rect 3550 3658 3554 3662
rect 3582 3658 3586 3662
rect 3590 3658 3594 3662
rect 3630 3658 3634 3662
rect 3646 3658 3650 3662
rect 3686 3658 3690 3662
rect 3742 3658 3746 3662
rect 3758 3658 3762 3662
rect 3814 3658 3818 3662
rect 3854 3658 3858 3662
rect 3878 3658 3882 3662
rect 3886 3658 3890 3662
rect 3934 3658 3938 3662
rect 3942 3658 3946 3662
rect 3990 3658 3994 3662
rect 4006 3658 4010 3662
rect 4014 3658 4018 3662
rect 4038 3658 4042 3662
rect 4054 3658 4058 3662
rect 4094 3658 4098 3662
rect 4158 3658 4162 3662
rect 4238 3658 4242 3662
rect 4254 3658 4258 3662
rect 4270 3658 4274 3662
rect 4310 3658 4314 3662
rect 4318 3658 4322 3662
rect 4374 3658 4378 3662
rect 4406 3658 4410 3662
rect 4414 3658 4418 3662
rect 4438 3658 4442 3662
rect 4494 3658 4498 3662
rect 4582 3658 4586 3662
rect 4662 3658 4666 3662
rect 4670 3658 4674 3662
rect 4694 3658 4698 3662
rect 4774 3658 4778 3662
rect 4854 3658 4858 3662
rect 4870 3658 4874 3662
rect 4918 3658 4922 3662
rect 4982 3658 4986 3662
rect 5022 3658 5026 3662
rect 5070 3658 5074 3662
rect 5086 3658 5090 3662
rect 5150 3658 5154 3662
rect 5190 3658 5194 3662
rect 374 3648 378 3652
rect 502 3648 506 3652
rect 662 3648 666 3652
rect 670 3648 674 3652
rect 894 3648 898 3652
rect 1078 3648 1082 3652
rect 1190 3648 1194 3652
rect 1478 3648 1482 3652
rect 1558 3648 1562 3652
rect 1614 3648 1618 3652
rect 1990 3648 1994 3652
rect 2182 3648 2186 3652
rect 2398 3648 2402 3652
rect 2518 3648 2522 3652
rect 2582 3648 2586 3652
rect 2686 3648 2690 3652
rect 2766 3648 2770 3652
rect 2782 3648 2786 3652
rect 2798 3648 2802 3652
rect 2926 3648 2930 3652
rect 2950 3648 2954 3652
rect 3038 3648 3042 3652
rect 3294 3648 3298 3652
rect 3534 3648 3538 3652
rect 3662 3648 3666 3652
rect 3974 3648 3978 3652
rect 4054 3648 4058 3652
rect 4214 3648 4218 3652
rect 4470 3648 4474 3652
rect 4494 3648 4498 3652
rect 4686 3648 4690 3652
rect 4814 3648 4818 3652
rect 4830 3648 4834 3652
rect 4838 3648 4842 3652
rect 150 3638 154 3642
rect 190 3638 194 3642
rect 1134 3638 1138 3642
rect 1318 3638 1322 3642
rect 3686 3638 3690 3642
rect 4118 3638 4122 3642
rect 4542 3638 4546 3642
rect 4710 3638 4714 3642
rect 4942 3638 4946 3642
rect 5126 3638 5130 3642
rect 1214 3628 1218 3632
rect 4630 3628 4634 3632
rect 382 3618 386 3622
rect 422 3618 426 3622
rect 454 3618 458 3622
rect 646 3618 650 3622
rect 710 3618 714 3622
rect 918 3618 922 3622
rect 1030 3618 1034 3622
rect 1150 3618 1154 3622
rect 1502 3618 1506 3622
rect 1582 3618 1586 3622
rect 1606 3618 1610 3622
rect 1774 3618 1778 3622
rect 1870 3618 1874 3622
rect 1966 3618 1970 3622
rect 2214 3618 2218 3622
rect 2294 3618 2298 3622
rect 2838 3618 2842 3622
rect 3238 3618 3242 3622
rect 3390 3618 3394 3622
rect 3478 3618 3482 3622
rect 3902 3618 3906 3622
rect 4022 3618 4026 3622
rect 4102 3618 4106 3622
rect 4206 3618 4210 3622
rect 4390 3618 4394 3622
rect 4422 3618 4426 3622
rect 4510 3618 4514 3622
rect 4854 3618 4858 3622
rect 538 3603 542 3607
rect 545 3603 549 3607
rect 1562 3603 1566 3607
rect 1569 3603 1573 3607
rect 2586 3603 2590 3607
rect 2593 3603 2597 3607
rect 3610 3603 3614 3607
rect 3617 3603 3621 3607
rect 4634 3603 4638 3607
rect 4641 3603 4645 3607
rect 470 3588 474 3592
rect 526 3588 530 3592
rect 606 3588 610 3592
rect 630 3588 634 3592
rect 934 3588 938 3592
rect 1246 3588 1250 3592
rect 1270 3588 1274 3592
rect 1326 3588 1330 3592
rect 1662 3588 1666 3592
rect 2454 3588 2458 3592
rect 3310 3588 3314 3592
rect 3350 3588 3354 3592
rect 3430 3588 3434 3592
rect 3734 3588 3738 3592
rect 3958 3588 3962 3592
rect 4398 3588 4402 3592
rect 4726 3588 4730 3592
rect 4774 3588 4778 3592
rect 5134 3588 5138 3592
rect 2710 3578 2714 3582
rect 2822 3578 2826 3582
rect 2982 3578 2986 3582
rect 150 3568 154 3572
rect 246 3568 250 3572
rect 262 3568 266 3572
rect 318 3568 322 3572
rect 510 3568 514 3572
rect 1134 3568 1138 3572
rect 1350 3568 1354 3572
rect 1454 3568 1458 3572
rect 1494 3568 1498 3572
rect 1958 3568 1962 3572
rect 1998 3568 2002 3572
rect 2118 3568 2122 3572
rect 2182 3568 2186 3572
rect 2726 3568 2730 3572
rect 2886 3568 2890 3572
rect 3286 3568 3290 3572
rect 3398 3568 3402 3572
rect 3774 3568 3778 3572
rect 3974 3568 3978 3572
rect 4974 3568 4978 3572
rect 5054 3568 5058 3572
rect 294 3558 298 3562
rect 334 3558 338 3562
rect 350 3558 354 3562
rect 414 3558 418 3562
rect 446 3558 450 3562
rect 582 3558 586 3562
rect 110 3548 114 3552
rect 198 3547 202 3551
rect 278 3548 282 3552
rect 294 3548 298 3552
rect 302 3548 306 3552
rect 318 3548 322 3552
rect 398 3548 402 3552
rect 430 3548 434 3552
rect 454 3548 458 3552
rect 494 3548 498 3552
rect 502 3548 506 3552
rect 542 3548 546 3552
rect 694 3558 698 3562
rect 878 3558 882 3562
rect 606 3548 610 3552
rect 646 3548 650 3552
rect 678 3548 682 3552
rect 734 3548 738 3552
rect 758 3548 762 3552
rect 798 3548 802 3552
rect 830 3548 834 3552
rect 878 3548 882 3552
rect 902 3558 906 3562
rect 926 3558 930 3562
rect 1150 3558 1154 3562
rect 1286 3558 1290 3562
rect 1406 3558 1410 3562
rect 950 3548 954 3552
rect 1022 3548 1026 3552
rect 1078 3548 1082 3552
rect 1134 3548 1138 3552
rect 1182 3547 1186 3551
rect 1254 3548 1258 3552
rect 1310 3548 1314 3552
rect 1374 3548 1378 3552
rect 1438 3548 1442 3552
rect 1622 3558 1626 3562
rect 1702 3558 1706 3562
rect 1814 3558 1818 3562
rect 1478 3548 1482 3552
rect 1550 3548 1554 3552
rect 1622 3548 1626 3552
rect 1638 3548 1642 3552
rect 1678 3548 1682 3552
rect 1774 3547 1778 3551
rect 1814 3548 1818 3552
rect 1838 3558 1842 3562
rect 1854 3548 1858 3552
rect 1902 3548 1906 3552
rect 1926 3548 1930 3552
rect 1974 3548 1978 3552
rect 1982 3548 1986 3552
rect 2134 3558 2138 3562
rect 2150 3558 2154 3562
rect 2390 3558 2394 3562
rect 2014 3548 2018 3552
rect 2054 3548 2058 3552
rect 2134 3548 2138 3552
rect 2150 3548 2154 3552
rect 2166 3548 2170 3552
rect 2238 3548 2242 3552
rect 2310 3548 2314 3552
rect 2694 3558 2698 3562
rect 2854 3558 2858 3562
rect 2870 3558 2874 3562
rect 3006 3558 3010 3562
rect 3054 3558 3058 3562
rect 3270 3558 3274 3562
rect 2414 3548 2418 3552
rect 2454 3548 2458 3552
rect 2566 3547 2570 3551
rect 2614 3548 2618 3552
rect 2662 3548 2666 3552
rect 2678 3548 2682 3552
rect 2710 3548 2714 3552
rect 2758 3547 2762 3551
rect 2790 3548 2794 3552
rect 2838 3548 2842 3552
rect 2854 3548 2858 3552
rect 2870 3548 2874 3552
rect 2918 3547 2922 3551
rect 3006 3548 3010 3552
rect 3022 3548 3026 3552
rect 3038 3548 3042 3552
rect 3062 3548 3066 3552
rect 3070 3548 3074 3552
rect 3094 3548 3098 3552
rect 3134 3548 3138 3552
rect 3150 3548 3154 3552
rect 3190 3548 3194 3552
rect 6 3538 10 3542
rect 86 3538 90 3542
rect 182 3538 186 3542
rect 270 3538 274 3542
rect 326 3538 330 3542
rect 350 3538 354 3542
rect 406 3538 410 3542
rect 422 3538 426 3542
rect 438 3538 442 3542
rect 486 3538 490 3542
rect 566 3538 570 3542
rect 614 3538 618 3542
rect 686 3538 690 3542
rect 806 3538 810 3542
rect 918 3538 922 3542
rect 942 3538 946 3542
rect 1054 3538 1058 3542
rect 1126 3538 1130 3542
rect 1166 3538 1170 3542
rect 1302 3538 1306 3542
rect 1422 3538 1426 3542
rect 1430 3538 1434 3542
rect 1486 3538 1490 3542
rect 1590 3538 1594 3542
rect 1646 3538 1650 3542
rect 1686 3538 1690 3542
rect 1790 3538 1794 3542
rect 1806 3538 1810 3542
rect 1862 3538 1866 3542
rect 1966 3538 1970 3542
rect 2030 3538 2034 3542
rect 2062 3538 2066 3542
rect 2094 3538 2098 3542
rect 2142 3538 2146 3542
rect 2174 3538 2178 3542
rect 2222 3538 2226 3542
rect 2262 3538 2266 3542
rect 2286 3538 2290 3542
rect 2374 3538 2378 3542
rect 2398 3538 2402 3542
rect 2478 3538 2482 3542
rect 2518 3538 2522 3542
rect 2582 3538 2586 3542
rect 2622 3538 2626 3542
rect 2646 3538 2650 3542
rect 2670 3538 2674 3542
rect 2694 3538 2698 3542
rect 2702 3538 2706 3542
rect 2830 3538 2834 3542
rect 2862 3538 2866 3542
rect 2934 3538 2938 3542
rect 3222 3547 3226 3551
rect 3286 3548 3290 3552
rect 3326 3548 3330 3552
rect 3334 3548 3338 3552
rect 3390 3548 3394 3552
rect 3414 3548 3418 3552
rect 3454 3558 3458 3562
rect 3494 3558 3498 3562
rect 3510 3548 3514 3552
rect 3526 3548 3530 3552
rect 3606 3548 3610 3552
rect 3654 3548 3658 3552
rect 3694 3558 3698 3562
rect 3902 3558 3906 3562
rect 3918 3558 3922 3562
rect 3926 3558 3930 3562
rect 4158 3558 4162 3562
rect 3750 3548 3754 3552
rect 3790 3548 3794 3552
rect 3830 3548 3834 3552
rect 3022 3538 3026 3542
rect 3030 3538 3034 3542
rect 3054 3538 3058 3542
rect 3102 3538 3106 3542
rect 3126 3538 3130 3542
rect 3302 3538 3306 3542
rect 3358 3538 3362 3542
rect 3382 3538 3386 3542
rect 3414 3538 3418 3542
rect 3422 3538 3426 3542
rect 3470 3538 3474 3542
rect 3478 3538 3482 3542
rect 3582 3538 3586 3542
rect 3630 3538 3634 3542
rect 3662 3538 3666 3542
rect 3678 3538 3682 3542
rect 3718 3538 3722 3542
rect 3758 3538 3762 3542
rect 3862 3547 3866 3551
rect 3902 3548 3906 3552
rect 3934 3548 3938 3552
rect 3942 3548 3946 3552
rect 4054 3548 4058 3552
rect 4094 3548 4098 3552
rect 4182 3558 4186 3562
rect 4222 3558 4226 3562
rect 4358 3558 4362 3562
rect 4182 3548 4186 3552
rect 4190 3548 4194 3552
rect 4302 3548 4306 3552
rect 4382 3558 4386 3562
rect 4558 3558 4562 3562
rect 4382 3548 4386 3552
rect 4470 3548 4474 3552
rect 4510 3548 4514 3552
rect 4526 3548 4530 3552
rect 4542 3548 4546 3552
rect 4638 3558 4642 3562
rect 4662 3558 4666 3562
rect 4678 3558 4682 3562
rect 4710 3558 4714 3562
rect 4742 3558 4746 3562
rect 4758 3558 4762 3562
rect 4902 3558 4906 3562
rect 4590 3548 4594 3552
rect 4614 3548 4618 3552
rect 4686 3548 4690 3552
rect 4702 3548 4706 3552
rect 4734 3548 4738 3552
rect 4758 3548 4762 3552
rect 4846 3548 4850 3552
rect 4926 3558 4930 3562
rect 5150 3558 5154 3562
rect 4926 3548 4930 3552
rect 5014 3548 5018 3552
rect 5078 3548 5082 3552
rect 5110 3548 5114 3552
rect 3894 3538 3898 3542
rect 3990 3538 3994 3542
rect 4038 3538 4042 3542
rect 4078 3538 4082 3542
rect 4142 3538 4146 3542
rect 4198 3538 4202 3542
rect 4238 3538 4242 3542
rect 4278 3538 4282 3542
rect 4310 3538 4314 3542
rect 4342 3538 4346 3542
rect 4494 3538 4498 3542
rect 4534 3538 4538 3542
rect 4566 3538 4570 3542
rect 4598 3538 4602 3542
rect 4662 3538 4666 3542
rect 4678 3538 4682 3542
rect 4734 3538 4738 3542
rect 4870 3538 4874 3542
rect 4886 3538 4890 3542
rect 4934 3538 4938 3542
rect 5014 3538 5018 3542
rect 5070 3538 5074 3542
rect 5086 3538 5090 3542
rect 5166 3538 5170 3542
rect 358 3528 362 3532
rect 374 3528 378 3532
rect 654 3528 658 3532
rect 814 3528 818 3532
rect 846 3528 850 3532
rect 854 3528 858 3532
rect 990 3528 994 3532
rect 1606 3528 1610 3532
rect 2030 3528 2034 3532
rect 2430 3528 2434 3532
rect 2630 3528 2634 3532
rect 2638 3528 2642 3532
rect 2654 3528 2658 3532
rect 2990 3528 2994 3532
rect 3254 3528 3258 3532
rect 3366 3528 3370 3532
rect 3966 3528 3970 3532
rect 4526 3528 4530 3532
rect 4598 3528 4602 3532
rect 4854 3528 4858 3532
rect 5126 3528 5130 3532
rect 5142 3528 5146 3532
rect 62 3518 66 3522
rect 166 3518 170 3522
rect 366 3518 370 3522
rect 790 3518 794 3522
rect 862 3518 866 3522
rect 966 3518 970 3522
rect 1118 3518 1122 3522
rect 1294 3518 1298 3522
rect 1326 3518 1330 3522
rect 1390 3518 1394 3522
rect 1414 3518 1418 3522
rect 1462 3518 1466 3522
rect 1622 3518 1626 3522
rect 1702 3518 1706 3522
rect 1710 3518 1714 3522
rect 2366 3518 2370 3522
rect 3086 3518 3090 3522
rect 3158 3518 3162 3522
rect 3262 3518 3266 3522
rect 3350 3518 3354 3522
rect 3398 3518 3402 3522
rect 3534 3518 3538 3522
rect 3766 3518 3770 3522
rect 3974 3518 3978 3522
rect 3998 3518 4002 3522
rect 4110 3518 4114 3522
rect 4222 3518 4226 3522
rect 4654 3518 4658 3522
rect 5062 3518 5066 3522
rect 5094 3518 5098 3522
rect 5134 3518 5138 3522
rect 5158 3518 5162 3522
rect 1050 3503 1054 3507
rect 1057 3503 1061 3507
rect 2074 3503 2078 3507
rect 2081 3503 2085 3507
rect 3098 3503 3102 3507
rect 3105 3503 3109 3507
rect 4114 3503 4118 3507
rect 4121 3503 4125 3507
rect 6 3488 10 3492
rect 190 3488 194 3492
rect 238 3488 242 3492
rect 358 3488 362 3492
rect 598 3488 602 3492
rect 694 3488 698 3492
rect 838 3488 842 3492
rect 1246 3488 1250 3492
rect 1270 3488 1274 3492
rect 1350 3488 1354 3492
rect 1398 3488 1402 3492
rect 1478 3488 1482 3492
rect 2030 3488 2034 3492
rect 2342 3488 2346 3492
rect 2558 3488 2562 3492
rect 2598 3488 2602 3492
rect 2894 3488 2898 3492
rect 3134 3488 3138 3492
rect 3366 3488 3370 3492
rect 3574 3488 3578 3492
rect 3686 3488 3690 3492
rect 4462 3488 4466 3492
rect 4566 3488 4570 3492
rect 4678 3488 4682 3492
rect 4694 3488 4698 3492
rect 4734 3488 4738 3492
rect 4798 3488 4802 3492
rect 5150 3488 5154 3492
rect 230 3478 234 3482
rect 462 3478 466 3482
rect 582 3478 586 3482
rect 62 3468 66 3472
rect 86 3468 90 3472
rect 126 3468 130 3472
rect 158 3468 162 3472
rect 166 3468 170 3472
rect 222 3468 226 3472
rect 262 3468 266 3472
rect 278 3468 282 3472
rect 366 3468 370 3472
rect 382 3468 386 3472
rect 414 3468 418 3472
rect 622 3468 626 3472
rect 638 3468 642 3472
rect 646 3468 650 3472
rect 678 3468 682 3472
rect 758 3468 762 3472
rect 782 3468 786 3472
rect 846 3468 850 3472
rect 862 3468 866 3472
rect 870 3468 874 3472
rect 934 3468 938 3472
rect 958 3468 962 3472
rect 990 3468 994 3472
rect 1046 3468 1050 3472
rect 1062 3468 1066 3472
rect 1078 3468 1082 3472
rect 1118 3468 1122 3472
rect 1166 3468 1170 3472
rect 1262 3468 1266 3472
rect 1286 3478 1290 3482
rect 1342 3478 1346 3482
rect 1366 3478 1370 3482
rect 1382 3478 1386 3482
rect 1302 3468 1306 3472
rect 1406 3468 1410 3472
rect 1702 3478 1706 3482
rect 2126 3478 2130 3482
rect 2534 3478 2538 3482
rect 1526 3468 1530 3472
rect 1606 3468 1610 3472
rect 1734 3468 1738 3472
rect 1982 3468 1986 3472
rect 1998 3468 2002 3472
rect 2078 3468 2082 3472
rect 2222 3468 2226 3472
rect 2278 3468 2282 3472
rect 2334 3468 2338 3472
rect 2422 3468 2426 3472
rect 2438 3468 2442 3472
rect 2494 3468 2498 3472
rect 2526 3468 2530 3472
rect 2566 3468 2570 3472
rect 2622 3468 2626 3472
rect 2678 3468 2682 3472
rect 2726 3468 2730 3472
rect 2790 3468 2794 3472
rect 2886 3468 2890 3472
rect 2910 3478 2914 3482
rect 2942 3478 2946 3482
rect 2974 3478 2978 3482
rect 3374 3478 3378 3482
rect 3430 3478 3434 3482
rect 3446 3478 3450 3482
rect 3662 3478 3666 3482
rect 3670 3478 3674 3482
rect 4038 3478 4042 3482
rect 4278 3478 4282 3482
rect 4686 3478 4690 3482
rect 4790 3478 4794 3482
rect 5014 3478 5018 3482
rect 5054 3478 5058 3482
rect 3046 3468 3050 3472
rect 3078 3468 3082 3472
rect 3102 3468 3106 3472
rect 3158 3468 3162 3472
rect 3206 3468 3210 3472
rect 3454 3468 3458 3472
rect 3582 3468 3586 3472
rect 3630 3468 3634 3472
rect 3662 3468 3666 3472
rect 3742 3468 3746 3472
rect 3782 3468 3786 3472
rect 70 3459 74 3463
rect 102 3458 106 3462
rect 118 3458 122 3462
rect 134 3458 138 3462
rect 158 3458 162 3462
rect 174 3458 178 3462
rect 214 3458 218 3462
rect 302 3458 306 3462
rect 326 3458 330 3462
rect 374 3458 378 3462
rect 446 3458 450 3462
rect 470 3458 474 3462
rect 502 3458 506 3462
rect 526 3458 530 3462
rect 542 3458 546 3462
rect 566 3458 570 3462
rect 574 3458 578 3462
rect 598 3458 602 3462
rect 654 3458 658 3462
rect 710 3458 714 3462
rect 734 3458 738 3462
rect 742 3458 746 3462
rect 798 3458 802 3462
rect 990 3458 994 3462
rect 1006 3458 1010 3462
rect 1030 3458 1034 3462
rect 1038 3458 1042 3462
rect 1070 3458 1074 3462
rect 1110 3458 1114 3462
rect 1126 3458 1130 3462
rect 1190 3458 1194 3462
rect 1254 3458 1258 3462
rect 1302 3458 1306 3462
rect 1318 3458 1322 3462
rect 1358 3458 1362 3462
rect 1366 3458 1370 3462
rect 1414 3458 1418 3462
rect 1446 3458 1450 3462
rect 1462 3458 1466 3462
rect 1502 3458 1506 3462
rect 1558 3458 1562 3462
rect 1598 3458 1602 3462
rect 1614 3458 1618 3462
rect 1622 3458 1626 3462
rect 1678 3458 1682 3462
rect 1726 3458 1730 3462
rect 1774 3458 1778 3462
rect 1790 3458 1794 3462
rect 1838 3458 1842 3462
rect 1846 3458 1850 3462
rect 1878 3458 1882 3462
rect 1926 3458 1930 3462
rect 1950 3459 1954 3463
rect 1990 3458 1994 3462
rect 2014 3458 2018 3462
rect 2038 3458 2042 3462
rect 2062 3458 2066 3462
rect 2102 3458 2106 3462
rect 2142 3458 2146 3462
rect 2166 3458 2170 3462
rect 2174 3458 2178 3462
rect 2214 3458 2218 3462
rect 2286 3458 2290 3462
rect 2294 3458 2298 3462
rect 2326 3458 2330 3462
rect 2406 3459 2410 3463
rect 2446 3458 2450 3462
rect 2454 3458 2458 3462
rect 2494 3458 2498 3462
rect 2502 3458 2506 3462
rect 2614 3458 2618 3462
rect 2630 3458 2634 3462
rect 2646 3458 2650 3462
rect 2670 3458 2674 3462
rect 2710 3459 2714 3463
rect 3910 3468 3914 3472
rect 3942 3468 3946 3472
rect 3958 3468 3962 3472
rect 4094 3468 4098 3472
rect 4134 3468 4138 3472
rect 4150 3468 4154 3472
rect 4206 3468 4210 3472
rect 4390 3468 4394 3472
rect 4446 3468 4450 3472
rect 4454 3468 4458 3472
rect 4510 3468 4514 3472
rect 4582 3468 4586 3472
rect 4702 3468 4706 3472
rect 4718 3468 4722 3472
rect 4750 3468 4754 3472
rect 4766 3468 4770 3472
rect 4854 3468 4858 3472
rect 4902 3468 4906 3472
rect 5030 3468 5034 3472
rect 5086 3468 5090 3472
rect 5158 3468 5162 3472
rect 2822 3458 2826 3462
rect 2878 3458 2882 3462
rect 2926 3458 2930 3462
rect 2982 3458 2986 3462
rect 3054 3458 3058 3462
rect 3094 3458 3098 3462
rect 3150 3458 3154 3462
rect 3198 3458 3202 3462
rect 3206 3458 3210 3462
rect 3230 3458 3234 3462
rect 3246 3458 3250 3462
rect 3254 3458 3258 3462
rect 3262 3458 3266 3462
rect 3270 3458 3274 3462
rect 3294 3458 3298 3462
rect 3318 3458 3322 3462
rect 3342 3458 3346 3462
rect 3350 3458 3354 3462
rect 3358 3458 3362 3462
rect 3406 3458 3410 3462
rect 3430 3458 3434 3462
rect 3454 3458 3458 3462
rect 3518 3458 3522 3462
rect 3542 3458 3546 3462
rect 3638 3458 3642 3462
rect 3742 3458 3746 3462
rect 3790 3458 3794 3462
rect 3806 3458 3810 3462
rect 3814 3458 3818 3462
rect 3822 3458 3826 3462
rect 3846 3458 3850 3462
rect 3870 3458 3874 3462
rect 3894 3458 3898 3462
rect 3902 3458 3906 3462
rect 3918 3458 3922 3462
rect 3950 3458 3954 3462
rect 4038 3459 4042 3463
rect 4086 3458 4090 3462
rect 4102 3458 4106 3462
rect 4118 3458 4122 3462
rect 4142 3458 4146 3462
rect 4198 3458 4202 3462
rect 4254 3458 4258 3462
rect 4310 3458 4314 3462
rect 4318 3458 4322 3462
rect 4350 3458 4354 3462
rect 4358 3458 4362 3462
rect 4398 3458 4402 3462
rect 4438 3458 4442 3462
rect 4518 3458 4522 3462
rect 4606 3458 4610 3462
rect 4710 3458 4714 3462
rect 4742 3458 4746 3462
rect 4774 3458 4778 3462
rect 4854 3458 4858 3462
rect 4894 3458 4898 3462
rect 4926 3458 4930 3462
rect 5006 3458 5010 3462
rect 5094 3458 5098 3462
rect 5166 3458 5170 3462
rect 102 3448 106 3452
rect 246 3448 250 3452
rect 262 3448 266 3452
rect 398 3448 402 3452
rect 422 3448 426 3452
rect 438 3448 442 3452
rect 622 3448 626 3452
rect 670 3448 674 3452
rect 694 3448 698 3452
rect 846 3448 850 3452
rect 942 3448 946 3452
rect 1094 3448 1098 3452
rect 1334 3448 1338 3452
rect 1390 3448 1394 3452
rect 1582 3448 1586 3452
rect 1662 3448 1666 3452
rect 1710 3448 1714 3452
rect 1998 3448 2002 3452
rect 2030 3448 2034 3452
rect 2086 3448 2090 3452
rect 2102 3448 2106 3452
rect 2310 3448 2314 3452
rect 2470 3448 2474 3452
rect 2550 3448 2554 3452
rect 2654 3448 2658 3452
rect 3070 3448 3074 3452
rect 3198 3448 3202 3452
rect 3382 3448 3386 3452
rect 3438 3448 3442 3452
rect 3478 3448 3482 3452
rect 3598 3448 3602 3452
rect 3806 3448 3810 3452
rect 3918 3448 3922 3452
rect 3934 3448 3938 3452
rect 3966 3448 3970 3452
rect 4070 3448 4074 3452
rect 4086 3448 4090 3452
rect 4102 3448 4106 3452
rect 4174 3448 4178 3452
rect 4414 3448 4418 3452
rect 4422 3448 4426 3452
rect 4470 3448 4474 3452
rect 4734 3448 4738 3452
rect 4918 3448 4922 3452
rect 5182 3448 5186 3452
rect 150 3438 154 3442
rect 198 3438 202 3442
rect 1230 3438 1234 3442
rect 1430 3438 1434 3442
rect 1886 3438 1890 3442
rect 2054 3438 2058 3442
rect 2254 3438 2258 3442
rect 2270 3438 2274 3442
rect 2630 3438 2634 3442
rect 2670 3438 2674 3442
rect 2774 3438 2778 3442
rect 3038 3438 3042 3442
rect 3174 3438 3178 3442
rect 4198 3438 4202 3442
rect 654 3428 658 3432
rect 3462 3428 3466 3432
rect 494 3418 498 3422
rect 558 3418 562 3422
rect 606 3418 610 3422
rect 630 3418 634 3422
rect 726 3418 730 3422
rect 982 3418 986 3422
rect 1022 3418 1026 3422
rect 1142 3418 1146 3422
rect 1318 3418 1322 3422
rect 1358 3418 1362 3422
rect 1542 3418 1546 3422
rect 1598 3418 1602 3422
rect 1638 3418 1642 3422
rect 1726 3418 1730 3422
rect 1830 3418 1834 3422
rect 1862 3418 1866 3422
rect 2158 3418 2162 3422
rect 2542 3418 2546 3422
rect 2870 3418 2874 3422
rect 2934 3418 2938 3422
rect 3278 3418 3282 3422
rect 3334 3418 3338 3422
rect 3398 3418 3402 3422
rect 3678 3418 3682 3422
rect 3830 3418 3834 3422
rect 3878 3418 3882 3422
rect 3974 3418 3978 3422
rect 4214 3418 4218 3422
rect 4326 3418 4330 3422
rect 4374 3418 4378 3422
rect 4398 3418 4402 3422
rect 4438 3418 4442 3422
rect 4950 3418 4954 3422
rect 5046 3418 5050 3422
rect 5166 3418 5170 3422
rect 538 3403 542 3407
rect 545 3403 549 3407
rect 1562 3403 1566 3407
rect 1569 3403 1573 3407
rect 2586 3403 2590 3407
rect 2593 3403 2597 3407
rect 3610 3403 3614 3407
rect 3617 3403 3621 3407
rect 4634 3403 4638 3407
rect 4641 3403 4645 3407
rect 1694 3388 1698 3392
rect 1934 3388 1938 3392
rect 1974 3388 1978 3392
rect 3422 3388 3426 3392
rect 3990 3388 3994 3392
rect 4102 3388 4106 3392
rect 4142 3388 4146 3392
rect 4446 3388 4450 3392
rect 4694 3388 4698 3392
rect 4726 3388 4730 3392
rect 4806 3388 4810 3392
rect 4990 3388 4994 3392
rect 5158 3388 5162 3392
rect 222 3378 226 3382
rect 750 3378 754 3382
rect 1542 3378 1546 3382
rect 1670 3378 1674 3382
rect 1822 3378 1826 3382
rect 5174 3378 5178 3382
rect 262 3368 266 3372
rect 382 3368 386 3372
rect 502 3368 506 3372
rect 550 3368 554 3372
rect 662 3368 666 3372
rect 710 3368 714 3372
rect 958 3368 962 3372
rect 1078 3368 1082 3372
rect 1158 3368 1162 3372
rect 1318 3368 1322 3372
rect 1574 3368 1578 3372
rect 1782 3368 1786 3372
rect 1838 3368 1842 3372
rect 1998 3368 2002 3372
rect 2038 3368 2042 3372
rect 2198 3368 2202 3372
rect 2302 3368 2306 3372
rect 2430 3368 2434 3372
rect 2814 3368 2818 3372
rect 2942 3368 2946 3372
rect 3086 3368 3090 3372
rect 3310 3368 3314 3372
rect 3326 3368 3330 3372
rect 3518 3368 3522 3372
rect 3710 3368 3714 3372
rect 4006 3368 4010 3372
rect 4062 3368 4066 3372
rect 4358 3368 4362 3372
rect 4934 3368 4938 3372
rect 5006 3368 5010 3372
rect 238 3358 242 3362
rect 94 3348 98 3352
rect 126 3348 130 3352
rect 174 3348 178 3352
rect 238 3348 242 3352
rect 518 3358 522 3362
rect 278 3348 282 3352
rect 318 3347 322 3351
rect 390 3348 394 3352
rect 446 3348 450 3352
rect 518 3348 522 3352
rect 574 3348 578 3352
rect 622 3348 626 3352
rect 694 3348 698 3352
rect 846 3358 850 3362
rect 1110 3358 1114 3362
rect 1142 3358 1146 3362
rect 1214 3358 1218 3362
rect 1310 3358 1314 3362
rect 1414 3358 1418 3362
rect 1430 3358 1434 3362
rect 1526 3358 1530 3362
rect 1710 3358 1714 3362
rect 1750 3358 1754 3362
rect 726 3348 730 3352
rect 734 3348 738 3352
rect 782 3348 786 3352
rect 806 3348 810 3352
rect 902 3348 906 3352
rect 966 3348 970 3352
rect 1022 3348 1026 3352
rect 1110 3348 1114 3352
rect 1126 3348 1130 3352
rect 1134 3348 1138 3352
rect 1166 3348 1170 3352
rect 1174 3348 1178 3352
rect 1214 3348 1218 3352
rect 1230 3348 1234 3352
rect 1254 3348 1258 3352
rect 1294 3348 1298 3352
rect 1350 3348 1354 3352
rect 1358 3348 1362 3352
rect 1454 3348 1458 3352
rect 1494 3348 1498 3352
rect 1510 3348 1514 3352
rect 1526 3348 1530 3352
rect 1534 3348 1538 3352
rect 6 3338 10 3342
rect 118 3338 122 3342
rect 230 3338 234 3342
rect 286 3338 290 3342
rect 326 3338 330 3342
rect 398 3338 402 3342
rect 422 3338 426 3342
rect 510 3338 514 3342
rect 582 3338 586 3342
rect 598 3338 602 3342
rect 686 3338 690 3342
rect 742 3338 746 3342
rect 862 3338 866 3342
rect 878 3338 882 3342
rect 998 3338 1002 3342
rect 1030 3338 1034 3342
rect 1102 3338 1106 3342
rect 1134 3338 1138 3342
rect 1230 3338 1234 3342
rect 1302 3338 1306 3342
rect 1430 3338 1434 3342
rect 1462 3338 1466 3342
rect 1470 3338 1474 3342
rect 1502 3338 1506 3342
rect 1606 3347 1610 3351
rect 1638 3348 1642 3352
rect 1678 3348 1682 3352
rect 1766 3348 1770 3352
rect 1798 3348 1802 3352
rect 1814 3348 1818 3352
rect 1878 3348 1882 3352
rect 1918 3348 1922 3352
rect 1950 3348 1954 3352
rect 1958 3348 1962 3352
rect 1974 3348 1978 3352
rect 2054 3358 2058 3362
rect 2022 3348 2026 3352
rect 2030 3348 2034 3352
rect 2038 3348 2042 3352
rect 1534 3338 1538 3342
rect 1590 3338 1594 3342
rect 1726 3338 1730 3342
rect 1734 3338 1738 3342
rect 1758 3338 1762 3342
rect 1814 3338 1818 3342
rect 1854 3338 1858 3342
rect 1902 3338 1906 3342
rect 1966 3338 1970 3342
rect 2022 3338 2026 3342
rect 2158 3347 2162 3351
rect 2190 3348 2194 3352
rect 2222 3358 2226 3362
rect 2270 3348 2274 3352
rect 2286 3348 2290 3352
rect 2326 3358 2330 3362
rect 2518 3358 2522 3362
rect 2534 3358 2538 3362
rect 2622 3358 2626 3362
rect 2830 3358 2834 3362
rect 2326 3348 2330 3352
rect 2366 3347 2370 3351
rect 2462 3348 2466 3352
rect 2502 3348 2506 3352
rect 2526 3348 2530 3352
rect 2550 3348 2554 3352
rect 2566 3348 2570 3352
rect 2670 3348 2674 3352
rect 2686 3348 2690 3352
rect 2758 3348 2762 3352
rect 2830 3348 2834 3352
rect 2854 3358 2858 3362
rect 2870 3348 2874 3352
rect 2886 3348 2890 3352
rect 2926 3348 2930 3352
rect 3046 3347 3050 3351
rect 3086 3348 3090 3352
rect 3126 3358 3130 3362
rect 3286 3358 3290 3362
rect 3206 3348 3210 3352
rect 3222 3348 3226 3352
rect 3270 3348 3274 3352
rect 3566 3358 3570 3362
rect 3582 3358 3586 3362
rect 3598 3358 3602 3362
rect 3742 3358 3746 3362
rect 3806 3358 3810 3362
rect 3318 3348 3322 3352
rect 3358 3348 3362 3352
rect 3374 3348 3378 3352
rect 3454 3348 3458 3352
rect 3478 3348 3482 3352
rect 3550 3348 3554 3352
rect 3582 3348 3586 3352
rect 3654 3348 3658 3352
rect 3726 3348 3730 3352
rect 3750 3348 3754 3352
rect 3942 3358 3946 3362
rect 4174 3358 4178 3362
rect 3830 3348 3834 3352
rect 3902 3348 3906 3352
rect 3958 3348 3962 3352
rect 3974 3348 3978 3352
rect 4030 3348 4034 3352
rect 4086 3348 4090 3352
rect 4158 3348 4162 3352
rect 4214 3358 4218 3362
rect 4414 3358 4418 3362
rect 4430 3358 4434 3362
rect 4542 3358 4546 3362
rect 4558 3358 4562 3362
rect 4574 3358 4578 3362
rect 4630 3358 4634 3362
rect 4846 3358 4850 3362
rect 4910 3358 4914 3362
rect 4942 3358 4946 3362
rect 4958 3358 4962 3362
rect 4974 3358 4978 3362
rect 5118 3358 5122 3362
rect 5166 3358 5170 3362
rect 4190 3348 4194 3352
rect 4198 3348 4202 3352
rect 4262 3348 4266 3352
rect 4302 3348 4306 3352
rect 4366 3348 4370 3352
rect 4390 3348 4394 3352
rect 4430 3348 4434 3352
rect 4502 3348 4506 3352
rect 4558 3348 4562 3352
rect 4590 3348 4594 3352
rect 4606 3348 4610 3352
rect 4622 3348 4626 3352
rect 4678 3348 4682 3352
rect 4710 3348 4714 3352
rect 4742 3348 4746 3352
rect 4750 3348 4754 3352
rect 4758 3348 4762 3352
rect 4782 3348 4786 3352
rect 4822 3348 4826 3352
rect 4854 3348 4858 3352
rect 4894 3348 4898 3352
rect 4918 3348 4922 3352
rect 4958 3348 4962 3352
rect 4990 3348 4994 3352
rect 5062 3348 5066 3352
rect 5110 3348 5114 3352
rect 5134 3348 5138 3352
rect 2062 3338 2066 3342
rect 2174 3338 2178 3342
rect 2190 3338 2194 3342
rect 2238 3338 2242 3342
rect 2254 3338 2258 3342
rect 2278 3338 2282 3342
rect 2334 3338 2338 3342
rect 2454 3338 2458 3342
rect 2486 3338 2490 3342
rect 2494 3338 2498 3342
rect 2526 3338 2530 3342
rect 2558 3338 2562 3342
rect 2606 3338 2610 3342
rect 2822 3338 2826 3342
rect 2878 3338 2882 3342
rect 2902 3338 2906 3342
rect 2942 3338 2946 3342
rect 2958 3338 2962 3342
rect 2974 3338 2978 3342
rect 3078 3338 3082 3342
rect 3142 3338 3146 3342
rect 3262 3338 3266 3342
rect 3318 3338 3322 3342
rect 3534 3338 3538 3342
rect 3542 3338 3546 3342
rect 3574 3338 3578 3342
rect 3630 3338 3634 3342
rect 3718 3338 3722 3342
rect 3782 3338 3786 3342
rect 3822 3338 3826 3342
rect 3838 3338 3842 3342
rect 3894 3338 3898 3342
rect 3966 3338 3970 3342
rect 4022 3338 4026 3342
rect 4062 3338 4066 3342
rect 4078 3338 4082 3342
rect 4150 3338 4154 3342
rect 4206 3338 4210 3342
rect 4230 3338 4234 3342
rect 4254 3338 4258 3342
rect 4310 3338 4314 3342
rect 4438 3338 4442 3342
rect 4510 3338 4514 3342
rect 4566 3338 4570 3342
rect 4598 3338 4602 3342
rect 4606 3338 4610 3342
rect 4830 3338 4834 3342
rect 4886 3338 4890 3342
rect 4918 3338 4922 3342
rect 4966 3338 4970 3342
rect 4998 3338 5002 3342
rect 5062 3338 5066 3342
rect 5086 3338 5090 3342
rect 5110 3338 5114 3342
rect 5142 3338 5146 3342
rect 5150 3338 5154 3342
rect 78 3328 82 3332
rect 158 3328 162 3332
rect 406 3328 410 3332
rect 982 3328 986 3332
rect 1278 3328 1282 3332
rect 1382 3328 1386 3332
rect 1606 3328 1610 3332
rect 2366 3328 2370 3332
rect 2518 3328 2522 3332
rect 3046 3328 3050 3332
rect 3566 3328 3570 3332
rect 4118 3328 4122 3332
rect 4238 3328 4242 3332
rect 4366 3328 4370 3332
rect 4382 3328 4386 3332
rect 4406 3328 4410 3332
rect 4662 3328 4666 3332
rect 5110 3328 5114 3332
rect 5182 3328 5186 3332
rect 62 3318 66 3322
rect 110 3318 114 3322
rect 678 3318 682 3322
rect 854 3318 858 3322
rect 974 3318 978 3322
rect 1190 3318 1194 3322
rect 1422 3318 1426 3322
rect 1438 3318 1442 3322
rect 1710 3318 1714 3322
rect 1750 3318 1754 3322
rect 2438 3318 2442 3322
rect 2582 3318 2586 3322
rect 2910 3318 2914 3322
rect 2950 3318 2954 3322
rect 3150 3318 3154 3322
rect 3526 3318 3530 3322
rect 3742 3318 3746 3322
rect 3766 3318 3770 3322
rect 3846 3318 3850 3322
rect 3942 3318 3946 3322
rect 3990 3318 3994 3322
rect 4006 3318 4010 3322
rect 4046 3318 4050 3322
rect 4142 3318 4146 3322
rect 4214 3318 4218 3322
rect 4246 3318 4250 3322
rect 4398 3318 4402 3322
rect 4446 3318 4450 3322
rect 4574 3318 4578 3322
rect 4766 3318 4770 3322
rect 4806 3318 4810 3322
rect 4846 3318 4850 3322
rect 4870 3318 4874 3322
rect 4934 3318 4938 3322
rect 1050 3303 1054 3307
rect 1057 3303 1061 3307
rect 2074 3303 2078 3307
rect 2081 3303 2085 3307
rect 3098 3303 3102 3307
rect 3105 3303 3109 3307
rect 4114 3303 4118 3307
rect 4121 3303 4125 3307
rect 214 3288 218 3292
rect 310 3288 314 3292
rect 678 3288 682 3292
rect 926 3288 930 3292
rect 1126 3288 1130 3292
rect 1310 3288 1314 3292
rect 1686 3288 1690 3292
rect 1934 3288 1938 3292
rect 2150 3288 2154 3292
rect 2822 3288 2826 3292
rect 3038 3288 3042 3292
rect 3062 3288 3066 3292
rect 3366 3288 3370 3292
rect 3606 3288 3610 3292
rect 3622 3288 3626 3292
rect 3926 3288 3930 3292
rect 4102 3288 4106 3292
rect 4662 3288 4666 3292
rect 4766 3288 4770 3292
rect 4798 3288 4802 3292
rect 4870 3288 4874 3292
rect 5158 3288 5162 3292
rect 286 3278 290 3282
rect 302 3278 306 3282
rect 414 3278 418 3282
rect 710 3278 714 3282
rect 934 3278 938 3282
rect 950 3278 954 3282
rect 982 3278 986 3282
rect 1198 3278 1202 3282
rect 1206 3278 1210 3282
rect 1710 3278 1714 3282
rect 2358 3278 2362 3282
rect 2654 3278 2658 3282
rect 2750 3278 2754 3282
rect 3030 3278 3034 3282
rect 3046 3278 3050 3282
rect 3150 3278 3154 3282
rect 3214 3278 3218 3282
rect 3406 3278 3410 3282
rect 3662 3278 3666 3282
rect 3718 3278 3722 3282
rect 4214 3278 4218 3282
rect 4230 3278 4234 3282
rect 4286 3278 4290 3282
rect 4454 3278 4458 3282
rect 4574 3278 4578 3282
rect 62 3268 66 3272
rect 118 3268 122 3272
rect 134 3268 138 3272
rect 158 3268 162 3272
rect 222 3268 226 3272
rect 286 3268 290 3272
rect 302 3268 306 3272
rect 318 3268 322 3272
rect 334 3268 338 3272
rect 382 3268 386 3272
rect 494 3268 498 3272
rect 598 3268 602 3272
rect 654 3268 658 3272
rect 670 3268 674 3272
rect 718 3268 722 3272
rect 742 3268 746 3272
rect 782 3268 786 3272
rect 830 3268 834 3272
rect 870 3268 874 3272
rect 910 3268 914 3272
rect 918 3268 922 3272
rect 1030 3268 1034 3272
rect 1150 3268 1154 3272
rect 1318 3268 1322 3272
rect 1334 3268 1338 3272
rect 1382 3268 1386 3272
rect 1470 3268 1474 3272
rect 1542 3268 1546 3272
rect 1606 3268 1610 3272
rect 1670 3268 1674 3272
rect 1758 3268 1762 3272
rect 1806 3268 1810 3272
rect 1854 3268 1858 3272
rect 1918 3268 1922 3272
rect 2006 3268 2010 3272
rect 2054 3268 2058 3272
rect 2070 3268 2074 3272
rect 2126 3268 2130 3272
rect 2182 3268 2186 3272
rect 2230 3268 2234 3272
rect 2294 3268 2298 3272
rect 2310 3268 2314 3272
rect 2350 3268 2354 3272
rect 2550 3268 2554 3272
rect 2574 3268 2578 3272
rect 2630 3268 2634 3272
rect 2646 3268 2650 3272
rect 2798 3268 2802 3272
rect 2846 3268 2850 3272
rect 2974 3268 2978 3272
rect 70 3259 74 3263
rect 158 3258 162 3262
rect 174 3258 178 3262
rect 230 3258 234 3262
rect 246 3258 250 3262
rect 278 3258 282 3262
rect 326 3258 330 3262
rect 342 3258 346 3262
rect 430 3258 434 3262
rect 518 3258 522 3262
rect 606 3258 610 3262
rect 614 3258 618 3262
rect 646 3258 650 3262
rect 662 3258 666 3262
rect 694 3258 698 3262
rect 726 3258 730 3262
rect 774 3259 778 3263
rect 846 3258 850 3262
rect 862 3258 866 3262
rect 894 3258 898 3262
rect 902 3258 906 3262
rect 966 3258 970 3262
rect 998 3258 1002 3262
rect 1054 3258 1058 3262
rect 1142 3258 1146 3262
rect 1174 3258 1178 3262
rect 1182 3258 1186 3262
rect 1230 3258 1234 3262
rect 1254 3258 1258 3262
rect 1270 3258 1274 3262
rect 1294 3258 1298 3262
rect 1334 3258 1338 3262
rect 1358 3258 1362 3262
rect 1366 3258 1370 3262
rect 1406 3258 1410 3262
rect 1478 3258 1482 3262
rect 1486 3258 1490 3262
rect 1518 3258 1522 3262
rect 1614 3259 1618 3263
rect 1646 3258 1650 3262
rect 1662 3258 1666 3262
rect 1702 3258 1706 3262
rect 1734 3258 1738 3262
rect 1790 3258 1794 3262
rect 1806 3258 1810 3262
rect 1838 3259 1842 3263
rect 3006 3268 3010 3272
rect 3102 3268 3106 3272
rect 3126 3268 3130 3272
rect 3270 3268 3274 3272
rect 3310 3268 3314 3272
rect 3374 3268 3378 3272
rect 3398 3268 3402 3272
rect 3422 3268 3426 3272
rect 3502 3268 3506 3272
rect 3598 3268 3602 3272
rect 3654 3268 3658 3272
rect 3758 3268 3762 3272
rect 3790 3268 3794 3272
rect 3862 3268 3866 3272
rect 3982 3268 3986 3272
rect 4150 3268 4154 3272
rect 4158 3268 4162 3272
rect 4206 3268 4210 3272
rect 4382 3268 4386 3272
rect 4398 3268 4402 3272
rect 4430 3268 4434 3272
rect 4446 3268 4450 3272
rect 4582 3268 4586 3272
rect 4638 3268 4642 3272
rect 4742 3268 4746 3272
rect 4822 3268 4826 3272
rect 4854 3268 4858 3272
rect 4878 3268 4882 3272
rect 4910 3268 4914 3272
rect 4926 3268 4930 3272
rect 5062 3268 5066 3272
rect 1950 3258 1954 3262
rect 2014 3258 2018 3262
rect 2062 3258 2066 3262
rect 2118 3258 2122 3262
rect 2134 3258 2138 3262
rect 2166 3258 2170 3262
rect 2238 3258 2242 3262
rect 2302 3258 2306 3262
rect 2342 3258 2346 3262
rect 2382 3258 2386 3262
rect 2438 3258 2442 3262
rect 2446 3258 2450 3262
rect 2486 3258 2490 3262
rect 2502 3258 2506 3262
rect 2558 3258 2562 3262
rect 2614 3258 2618 3262
rect 2646 3258 2650 3262
rect 2678 3258 2682 3262
rect 2734 3258 2738 3262
rect 2742 3258 2746 3262
rect 2766 3258 2770 3262
rect 2782 3258 2786 3262
rect 2806 3258 2810 3262
rect 2862 3258 2866 3262
rect 2886 3258 2890 3262
rect 2894 3258 2898 3262
rect 2902 3258 2906 3262
rect 2910 3258 2914 3262
rect 2934 3258 2938 3262
rect 2942 3258 2946 3262
rect 2966 3258 2970 3262
rect 2982 3258 2986 3262
rect 2998 3258 3002 3262
rect 3014 3258 3018 3262
rect 3030 3258 3034 3262
rect 3094 3258 3098 3262
rect 3102 3258 3106 3262
rect 3134 3258 3138 3262
rect 3182 3259 3186 3263
rect 3214 3258 3218 3262
rect 3270 3258 3274 3262
rect 3318 3258 3322 3262
rect 3390 3258 3394 3262
rect 3422 3258 3426 3262
rect 3462 3258 3466 3262
rect 3486 3258 3490 3262
rect 3494 3258 3498 3262
rect 3510 3258 3514 3262
rect 3534 3258 3538 3262
rect 3542 3258 3546 3262
rect 3550 3258 3554 3262
rect 3558 3258 3562 3262
rect 3582 3258 3586 3262
rect 3678 3258 3682 3262
rect 3694 3258 3698 3262
rect 3726 3258 3730 3262
rect 3750 3258 3754 3262
rect 3766 3258 3770 3262
rect 3798 3258 3802 3262
rect 3846 3259 3850 3263
rect 3942 3258 3946 3262
rect 3966 3258 3970 3262
rect 3974 3258 3978 3262
rect 3990 3258 3994 3262
rect 4046 3258 4050 3262
rect 4070 3258 4074 3262
rect 4118 3258 4122 3262
rect 4142 3258 4146 3262
rect 4214 3258 4218 3262
rect 4230 3258 4234 3262
rect 4238 3258 4242 3262
rect 4246 3258 4250 3262
rect 4286 3258 4290 3262
rect 4366 3259 4370 3263
rect 4406 3258 4410 3262
rect 4502 3258 4506 3262
rect 4518 3258 4522 3262
rect 4590 3258 4594 3262
rect 4630 3258 4634 3262
rect 4718 3258 4722 3262
rect 4782 3258 4786 3262
rect 4814 3258 4818 3262
rect 4822 3258 4826 3262
rect 4838 3258 4842 3262
rect 4894 3258 4898 3262
rect 4934 3258 4938 3262
rect 4998 3258 5002 3262
rect 5014 3258 5018 3262
rect 5086 3258 5090 3262
rect 5166 3258 5170 3262
rect 5190 3258 5194 3262
rect 102 3248 106 3252
rect 246 3248 250 3252
rect 254 3248 258 3252
rect 366 3248 370 3252
rect 742 3248 746 3252
rect 878 3248 882 3252
rect 1278 3248 1282 3252
rect 1302 3248 1306 3252
rect 1646 3248 1650 3252
rect 1750 3248 1754 3252
rect 1774 3248 1778 3252
rect 2094 3248 2098 3252
rect 2398 3248 2402 3252
rect 2590 3248 2594 3252
rect 2630 3248 2634 3252
rect 2694 3248 2698 3252
rect 2766 3248 2770 3252
rect 2830 3248 2834 3252
rect 2950 3248 2954 3252
rect 2966 3248 2970 3252
rect 2982 3248 2986 3252
rect 3374 3248 3378 3252
rect 3446 3248 3450 3252
rect 3678 3248 3682 3252
rect 3782 3248 3786 3252
rect 3798 3248 3802 3252
rect 3814 3248 3818 3252
rect 3894 3248 3898 3252
rect 4006 3248 4010 3252
rect 4110 3248 4114 3252
rect 4198 3248 4202 3252
rect 4430 3248 4434 3252
rect 4606 3248 4610 3252
rect 4630 3248 4634 3252
rect 4846 3248 4850 3252
rect 4870 3248 4874 3252
rect 4894 3248 4898 3252
rect 5190 3248 5194 3252
rect 6 3238 10 3242
rect 270 3238 274 3242
rect 574 3238 578 3242
rect 630 3238 634 3242
rect 1126 3238 1130 3242
rect 1206 3238 1210 3242
rect 1446 3238 1450 3242
rect 1502 3238 1506 3242
rect 1958 3238 1962 3242
rect 2286 3238 2290 3242
rect 2326 3238 2330 3242
rect 2542 3238 2546 3242
rect 2750 3238 2754 3242
rect 3630 3238 3634 3242
rect 3638 3238 3642 3242
rect 4174 3238 4178 3242
rect 1462 3228 1466 3232
rect 2150 3228 2154 3232
rect 3430 3228 3434 3232
rect 3766 3228 3770 3232
rect 110 3218 114 3222
rect 342 3218 346 3222
rect 478 3218 482 3222
rect 894 3218 898 3222
rect 1110 3218 1114 3222
rect 1190 3218 1194 3222
rect 1246 3218 1250 3222
rect 1550 3218 1554 3222
rect 1686 3218 1690 3222
rect 1734 3218 1738 3222
rect 1918 3218 1922 3222
rect 2430 3218 2434 3222
rect 2718 3218 2722 3222
rect 2878 3218 2882 3222
rect 3478 3218 3482 3222
rect 3566 3218 3570 3222
rect 3670 3218 3674 3222
rect 3950 3218 3954 3222
rect 3990 3218 3994 3222
rect 4262 3218 4266 3222
rect 4294 3218 4298 3222
rect 4302 3218 4306 3222
rect 4566 3218 4570 3222
rect 4798 3218 4802 3222
rect 4886 3218 4890 3222
rect 4958 3218 4962 3222
rect 538 3203 542 3207
rect 545 3203 549 3207
rect 1562 3203 1566 3207
rect 1569 3203 1573 3207
rect 2586 3203 2590 3207
rect 2593 3203 2597 3207
rect 3610 3203 3614 3207
rect 3617 3203 3621 3207
rect 4634 3203 4638 3207
rect 4641 3203 4645 3207
rect 374 3188 378 3192
rect 430 3188 434 3192
rect 886 3188 890 3192
rect 1078 3188 1082 3192
rect 1950 3188 1954 3192
rect 2750 3188 2754 3192
rect 2774 3188 2778 3192
rect 2950 3188 2954 3192
rect 2974 3188 2978 3192
rect 3990 3188 3994 3192
rect 4190 3188 4194 3192
rect 4310 3188 4314 3192
rect 5094 3188 5098 3192
rect 1110 3178 1114 3182
rect 1142 3178 1146 3182
rect 1214 3178 1218 3182
rect 1278 3178 1282 3182
rect 2918 3178 2922 3182
rect 3102 3178 3106 3182
rect 3238 3178 3242 3182
rect 326 3168 330 3172
rect 342 3168 346 3172
rect 454 3168 458 3172
rect 1046 3168 1050 3172
rect 1198 3168 1202 3172
rect 1382 3168 1386 3172
rect 1590 3168 1594 3172
rect 1766 3168 1770 3172
rect 2078 3168 2082 3172
rect 2606 3168 2610 3172
rect 2646 3168 2650 3172
rect 2806 3168 2810 3172
rect 2822 3168 2826 3172
rect 2982 3168 2986 3172
rect 62 3158 66 3162
rect 78 3158 82 3162
rect 118 3158 122 3162
rect 358 3158 362 3162
rect 398 3158 402 3162
rect 22 3148 26 3152
rect 62 3148 66 3152
rect 86 3148 90 3152
rect 102 3148 106 3152
rect 118 3148 122 3152
rect 174 3148 178 3152
rect 198 3148 202 3152
rect 278 3148 282 3152
rect 342 3148 346 3152
rect 390 3148 394 3152
rect 422 3148 426 3152
rect 566 3158 570 3162
rect 686 3158 690 3162
rect 718 3158 722 3162
rect 734 3158 738 3162
rect 830 3158 834 3162
rect 902 3158 906 3162
rect 1126 3158 1130 3162
rect 1158 3158 1162 3162
rect 1254 3158 1258 3162
rect 470 3148 474 3152
rect 486 3148 490 3152
rect 550 3148 554 3152
rect 582 3148 586 3152
rect 630 3148 634 3152
rect 702 3148 706 3152
rect 774 3148 778 3152
rect 798 3148 802 3152
rect 806 3148 810 3152
rect 838 3148 842 3152
rect 870 3148 874 3152
rect 950 3148 954 3152
rect 990 3148 994 3152
rect 1094 3148 1098 3152
rect 1110 3148 1114 3152
rect 1142 3148 1146 3152
rect 1166 3148 1170 3152
rect 1182 3148 1186 3152
rect 1238 3148 1242 3152
rect 1502 3158 1506 3162
rect 1278 3148 1282 3152
rect 54 3138 58 3142
rect 94 3138 98 3142
rect 1318 3147 1322 3151
rect 1350 3148 1354 3152
rect 1454 3147 1458 3151
rect 1534 3148 1538 3152
rect 1574 3158 1578 3162
rect 3742 3168 3746 3172
rect 3758 3168 3762 3172
rect 3830 3168 3834 3172
rect 4006 3168 4010 3172
rect 4486 3168 4490 3172
rect 4830 3168 4834 3172
rect 4918 3168 4922 3172
rect 4958 3168 4962 3172
rect 1678 3158 1682 3162
rect 1694 3158 1698 3162
rect 1606 3148 1610 3152
rect 1614 3148 1618 3152
rect 1630 3148 1634 3152
rect 1638 3148 1642 3152
rect 1662 3148 1666 3152
rect 1702 3148 1706 3152
rect 1718 3148 1722 3152
rect 1734 3148 1738 3152
rect 1830 3147 1834 3151
rect 1886 3148 1890 3152
rect 1902 3148 1906 3152
rect 1942 3148 1946 3152
rect 1966 3148 1970 3152
rect 2006 3148 2010 3152
rect 2318 3158 2322 3162
rect 2358 3158 2362 3162
rect 2110 3148 2114 3152
rect 2126 3148 2130 3152
rect 2158 3148 2162 3152
rect 2166 3148 2170 3152
rect 2214 3148 2218 3152
rect 2254 3148 2258 3152
rect 2366 3148 2370 3152
rect 2422 3148 2426 3152
rect 2446 3148 2450 3152
rect 2486 3148 2490 3152
rect 2518 3148 2522 3152
rect 2526 3148 2530 3152
rect 2534 3148 2538 3152
rect 2574 3148 2578 3152
rect 2790 3158 2794 3162
rect 3014 3158 3018 3162
rect 3046 3158 3050 3162
rect 2630 3148 2634 3152
rect 2702 3148 2706 3152
rect 2742 3148 2746 3152
rect 2774 3148 2778 3152
rect 2806 3148 2810 3152
rect 2854 3147 2858 3151
rect 2886 3148 2890 3152
rect 2942 3148 2946 3152
rect 2998 3148 3002 3152
rect 3022 3148 3026 3152
rect 3214 3158 3218 3162
rect 3062 3148 3066 3152
rect 3070 3148 3074 3152
rect 3158 3148 3162 3152
rect 3350 3158 3354 3162
rect 3390 3158 3394 3162
rect 3470 3158 3474 3162
rect 3790 3158 3794 3162
rect 3238 3148 3242 3152
rect 3278 3147 3282 3151
rect 3374 3148 3378 3152
rect 3398 3148 3402 3152
rect 3446 3148 3450 3152
rect 3534 3148 3538 3152
rect 3574 3148 3578 3152
rect 3606 3148 3610 3152
rect 3622 3148 3626 3152
rect 3702 3148 3706 3152
rect 3758 3148 3762 3152
rect 3950 3158 3954 3162
rect 3806 3148 3810 3152
rect 3814 3148 3818 3152
rect 3862 3148 3866 3152
rect 3886 3148 3890 3152
rect 3934 3148 3938 3152
rect 3966 3148 3970 3152
rect 3974 3148 3978 3152
rect 4046 3148 4050 3152
rect 4134 3148 4138 3152
rect 4158 3148 4162 3152
rect 4198 3148 4202 3152
rect 4246 3148 4250 3152
rect 4262 3148 4266 3152
rect 4286 3148 4290 3152
rect 4294 3148 4298 3152
rect 4686 3158 4690 3162
rect 4742 3158 4746 3162
rect 4934 3158 4938 3162
rect 4966 3158 4970 3162
rect 4982 3158 4986 3162
rect 4398 3147 4402 3151
rect 4510 3148 4514 3152
rect 4550 3148 4554 3152
rect 4614 3148 4618 3152
rect 4686 3148 4690 3152
rect 4702 3148 4706 3152
rect 4726 3148 4730 3152
rect 4782 3148 4786 3152
rect 4870 3148 4874 3152
rect 4918 3148 4922 3152
rect 4982 3148 4986 3152
rect 5030 3148 5034 3152
rect 5054 3148 5058 3152
rect 5134 3148 5138 3152
rect 5150 3148 5154 3152
rect 334 3138 338 3142
rect 414 3138 418 3142
rect 422 3138 426 3142
rect 478 3138 482 3142
rect 526 3138 530 3142
rect 686 3138 690 3142
rect 718 3138 722 3142
rect 734 3138 738 3142
rect 758 3138 762 3142
rect 814 3138 818 3142
rect 862 3138 866 3142
rect 918 3138 922 3142
rect 1102 3138 1106 3142
rect 1134 3138 1138 3142
rect 1166 3138 1170 3142
rect 1190 3138 1194 3142
rect 1230 3138 1234 3142
rect 1286 3138 1290 3142
rect 1446 3138 1450 3142
rect 1502 3138 1506 3142
rect 1518 3138 1522 3142
rect 1526 3138 1530 3142
rect 1590 3138 1594 3142
rect 1622 3138 1626 3142
rect 1694 3138 1698 3142
rect 1726 3138 1730 3142
rect 1846 3138 1850 3142
rect 1862 3138 1866 3142
rect 1910 3138 1914 3142
rect 1926 3138 1930 3142
rect 2014 3138 2018 3142
rect 2086 3138 2090 3142
rect 2134 3138 2138 3142
rect 2150 3138 2154 3142
rect 2198 3138 2202 3142
rect 2206 3138 2210 3142
rect 2246 3138 2250 3142
rect 2334 3138 2338 3142
rect 2542 3138 2546 3142
rect 2566 3138 2570 3142
rect 2606 3138 2610 3142
rect 2638 3138 2642 3142
rect 2726 3138 2730 3142
rect 2766 3138 2770 3142
rect 2798 3138 2802 3142
rect 2934 3138 2938 3142
rect 2966 3138 2970 3142
rect 2990 3138 2994 3142
rect 3022 3138 3026 3142
rect 3078 3138 3082 3142
rect 3182 3138 3186 3142
rect 3198 3138 3202 3142
rect 3246 3138 3250 3142
rect 3294 3138 3298 3142
rect 3366 3138 3370 3142
rect 3382 3138 3386 3142
rect 3438 3138 3442 3142
rect 3454 3138 3458 3142
rect 3558 3138 3562 3142
rect 3582 3138 3586 3142
rect 3702 3138 3706 3142
rect 3742 3138 3746 3142
rect 3766 3138 3770 3142
rect 3822 3138 3826 3142
rect 3894 3138 3898 3142
rect 3926 3138 3930 3142
rect 3982 3138 3986 3142
rect 4070 3138 4074 3142
rect 4206 3138 4210 3142
rect 4366 3138 4370 3142
rect 4382 3138 4386 3142
rect 4414 3138 4418 3142
rect 4470 3138 4474 3142
rect 4518 3138 4522 3142
rect 4670 3138 4674 3142
rect 4758 3138 4762 3142
rect 4774 3138 4778 3142
rect 4894 3138 4898 3142
rect 4910 3138 4914 3142
rect 4942 3138 4946 3142
rect 4990 3138 4994 3142
rect 6 3128 10 3132
rect 126 3128 130 3132
rect 206 3128 210 3132
rect 502 3128 506 3132
rect 614 3128 618 3132
rect 982 3128 986 3132
rect 1486 3128 1490 3132
rect 1886 3128 1890 3132
rect 2110 3128 2114 3132
rect 2182 3128 2186 3132
rect 2550 3128 2554 3132
rect 2558 3128 2562 3132
rect 2758 3128 2762 3132
rect 2958 3128 2962 3132
rect 3414 3128 3418 3132
rect 3430 3128 3434 3132
rect 4230 3128 4234 3132
rect 4622 3128 4626 3132
rect 4710 3128 4714 3132
rect 38 3118 42 3122
rect 406 3118 410 3122
rect 518 3118 522 3122
rect 678 3118 682 3122
rect 726 3118 730 3122
rect 742 3118 746 3122
rect 790 3118 794 3122
rect 822 3118 826 3122
rect 886 3118 890 3122
rect 910 3118 914 3122
rect 934 3118 938 3122
rect 1390 3118 1394 3122
rect 1510 3118 1514 3122
rect 1550 3118 1554 3122
rect 1654 3118 1658 3122
rect 1686 3118 1690 3122
rect 1750 3118 1754 3122
rect 1878 3118 1882 3122
rect 2094 3118 2098 3122
rect 2310 3118 2314 3122
rect 2374 3118 2378 3122
rect 2502 3118 2506 3122
rect 3014 3118 3018 3122
rect 3470 3118 3474 3122
rect 3646 3118 3650 3122
rect 4214 3118 4218 3122
rect 4270 3118 4274 3122
rect 4462 3118 4466 3122
rect 4494 3118 4498 3122
rect 4534 3118 4538 3122
rect 4558 3118 4562 3122
rect 4686 3118 4690 3122
rect 4798 3118 4802 3122
rect 4958 3118 4962 3122
rect 4998 3118 5002 3122
rect 1050 3103 1054 3107
rect 1057 3103 1061 3107
rect 2074 3103 2078 3107
rect 2081 3103 2085 3107
rect 3098 3103 3102 3107
rect 3105 3103 3109 3107
rect 4114 3103 4118 3107
rect 4121 3103 4125 3107
rect 6 3088 10 3092
rect 110 3088 114 3092
rect 174 3088 178 3092
rect 390 3088 394 3092
rect 606 3088 610 3092
rect 694 3088 698 3092
rect 718 3088 722 3092
rect 838 3088 842 3092
rect 894 3088 898 3092
rect 1078 3088 1082 3092
rect 1118 3088 1122 3092
rect 1238 3088 1242 3092
rect 1310 3088 1314 3092
rect 1414 3088 1418 3092
rect 1446 3088 1450 3092
rect 1630 3088 1634 3092
rect 1750 3088 1754 3092
rect 1782 3088 1786 3092
rect 1974 3088 1978 3092
rect 2126 3088 2130 3092
rect 2558 3088 2562 3092
rect 2614 3088 2618 3092
rect 2710 3088 2714 3092
rect 3014 3088 3018 3092
rect 3022 3088 3026 3092
rect 3054 3088 3058 3092
rect 3286 3088 3290 3092
rect 3334 3088 3338 3092
rect 3350 3088 3354 3092
rect 3734 3088 3738 3092
rect 3902 3088 3906 3092
rect 4102 3088 4106 3092
rect 4214 3088 4218 3092
rect 4390 3088 4394 3092
rect 4614 3088 4618 3092
rect 4718 3088 4722 3092
rect 4878 3088 4882 3092
rect 5006 3088 5010 3092
rect 5046 3088 5050 3092
rect 614 3078 618 3082
rect 710 3078 714 3082
rect 726 3078 730 3082
rect 1302 3078 1306 3082
rect 1390 3078 1394 3082
rect 1406 3078 1410 3082
rect 1438 3078 1442 3082
rect 1470 3078 1474 3082
rect 1486 3078 1490 3082
rect 1526 3078 1530 3082
rect 1638 3078 1642 3082
rect 1646 3078 1650 3082
rect 1662 3078 1666 3082
rect 1958 3078 1962 3082
rect 86 3068 90 3072
rect 118 3068 122 3072
rect 270 3068 274 3072
rect 294 3068 298 3072
rect 310 3068 314 3072
rect 46 3058 50 3062
rect 126 3058 130 3062
rect 158 3058 162 3062
rect 166 3058 170 3062
rect 206 3058 210 3062
rect 238 3059 242 3063
rect 286 3058 290 3062
rect 382 3068 386 3072
rect 414 3068 418 3072
rect 454 3068 458 3072
rect 646 3068 650 3072
rect 678 3068 682 3072
rect 702 3068 706 3072
rect 862 3068 866 3072
rect 942 3068 946 3072
rect 958 3068 962 3072
rect 974 3068 978 3072
rect 1038 3068 1042 3072
rect 1094 3068 1098 3072
rect 1182 3068 1186 3072
rect 1206 3068 1210 3072
rect 1286 3068 1290 3072
rect 1334 3068 1338 3072
rect 1350 3068 1354 3072
rect 1358 3068 1362 3072
rect 1438 3068 1442 3072
rect 1454 3068 1458 3072
rect 1622 3068 1626 3072
rect 1670 3068 1674 3072
rect 326 3058 330 3062
rect 334 3058 338 3062
rect 374 3058 378 3062
rect 406 3058 410 3062
rect 422 3058 426 3062
rect 430 3058 434 3062
rect 462 3058 466 3062
rect 470 3058 474 3062
rect 542 3059 546 3063
rect 1702 3068 1706 3072
rect 1846 3068 1850 3072
rect 1902 3068 1906 3072
rect 1918 3068 1922 3072
rect 1942 3068 1946 3072
rect 2070 3068 2074 3072
rect 2078 3068 2082 3072
rect 2126 3068 2130 3072
rect 2142 3068 2146 3072
rect 2150 3068 2154 3072
rect 2246 3068 2250 3072
rect 2262 3068 2266 3072
rect 2310 3068 2314 3072
rect 2414 3068 2418 3072
rect 2430 3068 2434 3072
rect 2470 3078 2474 3082
rect 3446 3078 3450 3082
rect 3502 3078 3506 3082
rect 3590 3078 3594 3082
rect 3702 3078 3706 3082
rect 3830 3078 3834 3082
rect 3918 3078 3922 3082
rect 4422 3078 4426 3082
rect 4678 3078 4682 3082
rect 2486 3068 2490 3072
rect 2510 3068 2514 3072
rect 2518 3068 2522 3072
rect 2566 3068 2570 3072
rect 2574 3068 2578 3072
rect 2694 3068 2698 3072
rect 2774 3068 2778 3072
rect 2806 3068 2810 3072
rect 2830 3068 2834 3072
rect 2846 3068 2850 3072
rect 2862 3068 2866 3072
rect 2886 3068 2890 3072
rect 2894 3068 2898 3072
rect 3038 3068 3042 3072
rect 3046 3068 3050 3072
rect 3310 3068 3314 3072
rect 3326 3068 3330 3072
rect 3406 3068 3410 3072
rect 3462 3068 3466 3072
rect 574 3058 578 3062
rect 670 3058 674 3062
rect 774 3058 778 3062
rect 798 3058 802 3062
rect 854 3058 858 3062
rect 870 3058 874 3062
rect 878 3058 882 3062
rect 902 3058 906 3062
rect 910 3058 914 3062
rect 942 3058 946 3062
rect 950 3058 954 3062
rect 982 3058 986 3062
rect 990 3058 994 3062
rect 998 3058 1002 3062
rect 1022 3058 1026 3062
rect 1030 3058 1034 3062
rect 1102 3058 1106 3062
rect 1142 3058 1146 3062
rect 1166 3058 1170 3062
rect 1174 3058 1178 3062
rect 1182 3058 1186 3062
rect 1214 3058 1218 3062
rect 1222 3058 1226 3062
rect 1230 3058 1234 3062
rect 1254 3058 1258 3062
rect 1270 3058 1274 3062
rect 1318 3058 1322 3062
rect 1342 3058 1346 3062
rect 1358 3058 1362 3062
rect 1390 3058 1394 3062
rect 1406 3058 1410 3062
rect 1462 3058 1466 3062
rect 1534 3058 1538 3062
rect 1598 3058 1602 3062
rect 1662 3058 1666 3062
rect 1678 3058 1682 3062
rect 1694 3058 1698 3062
rect 1710 3058 1714 3062
rect 1734 3058 1738 3062
rect 1766 3058 1770 3062
rect 1806 3058 1810 3062
rect 1830 3058 1834 3062
rect 1838 3058 1842 3062
rect 1854 3058 1858 3062
rect 1878 3058 1882 3062
rect 1886 3058 1890 3062
rect 1910 3058 1914 3062
rect 1990 3058 1994 3062
rect 1998 3058 2002 3062
rect 2006 3058 2010 3062
rect 2030 3058 2034 3062
rect 2054 3058 2058 3062
rect 2062 3058 2066 3062
rect 2118 3058 2122 3062
rect 2230 3059 2234 3063
rect 2262 3058 2266 3062
rect 2310 3058 2314 3062
rect 2350 3058 2354 3062
rect 2374 3058 2378 3062
rect 2454 3058 2458 3062
rect 2486 3058 2490 3062
rect 2526 3058 2530 3062
rect 2534 3058 2538 3062
rect 2550 3058 2554 3062
rect 2574 3058 2578 3062
rect 2654 3058 2658 3062
rect 2766 3058 2770 3062
rect 2822 3058 2826 3062
rect 2854 3058 2858 3062
rect 2870 3058 2874 3062
rect 2902 3058 2906 3062
rect 2950 3059 2954 3063
rect 2982 3058 2986 3062
rect 3070 3058 3074 3062
rect 3086 3058 3090 3062
rect 3102 3058 3106 3062
rect 3110 3058 3114 3062
rect 3134 3058 3138 3062
rect 3142 3058 3146 3062
rect 3166 3058 3170 3062
rect 3214 3058 3218 3062
rect 3238 3058 3242 3062
rect 3302 3058 3306 3062
rect 3414 3059 3418 3063
rect 3494 3068 3498 3072
rect 3518 3068 3522 3072
rect 3534 3068 3538 3072
rect 3622 3068 3626 3072
rect 3718 3068 3722 3072
rect 3814 3068 3818 3072
rect 3854 3068 3858 3072
rect 3870 3068 3874 3072
rect 4030 3068 4034 3072
rect 4046 3068 4050 3072
rect 4062 3068 4066 3072
rect 4086 3068 4090 3072
rect 4158 3068 4162 3072
rect 4270 3068 4274 3072
rect 4294 3068 4298 3072
rect 4382 3068 4386 3072
rect 4454 3068 4458 3072
rect 4486 3068 4490 3072
rect 4494 3068 4498 3072
rect 4518 3068 4522 3072
rect 4574 3068 4578 3072
rect 4606 3068 4610 3072
rect 4638 3068 4642 3072
rect 5014 3078 5018 3082
rect 5142 3078 5146 3082
rect 4702 3068 4706 3072
rect 4798 3068 4802 3072
rect 4814 3068 4818 3072
rect 4870 3068 4874 3072
rect 4998 3068 5002 3072
rect 5022 3068 5026 3072
rect 5070 3068 5074 3072
rect 5078 3068 5082 3072
rect 5094 3068 5098 3072
rect 5174 3068 5178 3072
rect 3462 3058 3466 3062
rect 3470 3058 3474 3062
rect 3486 3058 3490 3062
rect 3526 3058 3530 3062
rect 3566 3058 3570 3062
rect 3574 3058 3578 3062
rect 3590 3058 3594 3062
rect 3694 3058 3698 3062
rect 3774 3058 3778 3062
rect 3798 3059 3802 3063
rect 3846 3058 3850 3062
rect 3878 3058 3882 3062
rect 3886 3058 3890 3062
rect 3934 3058 3938 3062
rect 3942 3058 3946 3062
rect 3982 3058 3986 3062
rect 3990 3058 3994 3062
rect 4014 3058 4018 3062
rect 4022 3058 4026 3062
rect 4038 3058 4042 3062
rect 4166 3058 4170 3062
rect 4230 3058 4234 3062
rect 4254 3058 4258 3062
rect 4262 3058 4266 3062
rect 4302 3058 4306 3062
rect 4318 3058 4322 3062
rect 4326 3058 4330 3062
rect 4334 3058 4338 3062
rect 4358 3058 4362 3062
rect 4374 3058 4378 3062
rect 4406 3058 4410 3062
rect 4430 3058 4434 3062
rect 4478 3058 4482 3062
rect 4526 3058 4530 3062
rect 4566 3058 4570 3062
rect 4606 3058 4610 3062
rect 4630 3058 4634 3062
rect 4654 3058 4658 3062
rect 4710 3058 4714 3062
rect 4774 3058 4778 3062
rect 4814 3058 4818 3062
rect 4862 3058 4866 3062
rect 4910 3058 4914 3062
rect 4926 3058 4930 3062
rect 4982 3058 4986 3062
rect 4990 3058 4994 3062
rect 5062 3058 5066 3062
rect 5118 3058 5122 3062
rect 5126 3058 5130 3062
rect 5142 3058 5146 3062
rect 5166 3058 5170 3062
rect 102 3048 106 3052
rect 390 3048 394 3052
rect 630 3048 634 3052
rect 686 3048 690 3052
rect 838 3048 842 3052
rect 1326 3048 1330 3052
rect 1382 3048 1386 3052
rect 1694 3048 1698 3052
rect 1726 3048 1730 3052
rect 1894 3048 1898 3052
rect 1926 3048 1930 3052
rect 1942 3048 1946 3052
rect 2046 3048 2050 3052
rect 2094 3048 2098 3052
rect 2126 3048 2130 3052
rect 2270 3048 2274 3052
rect 2286 3048 2290 3052
rect 2294 3048 2298 3052
rect 2430 3048 2434 3052
rect 2494 3048 2498 3052
rect 2542 3048 2546 3052
rect 2590 3048 2594 3052
rect 2886 3048 2890 3052
rect 2902 3048 2906 3052
rect 2918 3048 2922 3052
rect 3022 3048 3026 3052
rect 3062 3048 3066 3052
rect 3318 3048 3322 3052
rect 3342 3048 3346 3052
rect 3470 3048 3474 3052
rect 3550 3048 3554 3052
rect 4102 3048 4106 3052
rect 4238 3048 4242 3052
rect 4286 3048 4290 3052
rect 4318 3048 4322 3052
rect 4446 3048 4450 3052
rect 4462 3048 4466 3052
rect 4510 3048 4514 3052
rect 4550 3048 4554 3052
rect 4582 3048 4586 3052
rect 4614 3048 4618 3052
rect 4838 3048 4842 3052
rect 4974 3048 4978 3052
rect 5038 3048 5042 3052
rect 5094 3048 5098 3052
rect 5150 3048 5154 3052
rect 358 3038 362 3042
rect 1078 3038 1082 3042
rect 1470 3038 1474 3042
rect 1590 3038 1594 3042
rect 2406 3038 2410 3042
rect 2510 3038 2514 3042
rect 3502 3038 3506 3042
rect 4086 3038 4090 3042
rect 4278 3038 4282 3042
rect 4342 3038 4346 3042
rect 4494 3038 4498 3042
rect 4734 3038 4738 3042
rect 4862 3038 4866 3042
rect 4894 3038 4898 3042
rect 622 3028 626 3032
rect 4598 3028 4602 3032
rect 4686 3028 4690 3032
rect 150 3018 154 3022
rect 334 3018 338 3022
rect 486 3018 490 3022
rect 670 3018 674 3022
rect 718 3018 722 3022
rect 934 3018 938 3022
rect 958 3018 962 3022
rect 1014 3018 1018 3022
rect 1118 3018 1122 3022
rect 1158 3018 1162 3022
rect 1190 3018 1194 3022
rect 1366 3018 1370 3022
rect 1494 3018 1498 3022
rect 1710 3018 1714 3022
rect 1782 3018 1786 3022
rect 1822 3018 1826 3022
rect 1950 3018 1954 3022
rect 2022 3018 2026 3022
rect 2422 3018 2426 3022
rect 2614 3018 2618 3022
rect 3158 3018 3162 3022
rect 3598 3018 3602 3022
rect 3926 3018 3930 3022
rect 3958 3018 3962 3022
rect 4006 3018 4010 3022
rect 4214 3018 4218 3022
rect 4526 3018 4530 3022
rect 538 3003 542 3007
rect 545 3003 549 3007
rect 1562 3003 1566 3007
rect 1569 3003 1573 3007
rect 2586 3003 2590 3007
rect 2593 3003 2597 3007
rect 3610 3003 3614 3007
rect 3617 3003 3621 3007
rect 4634 3003 4638 3007
rect 4641 3003 4645 3007
rect 830 2988 834 2992
rect 902 2988 906 2992
rect 1038 2988 1042 2992
rect 1486 2988 1490 2992
rect 1766 2988 1770 2992
rect 1982 2988 1986 2992
rect 2278 2988 2282 2992
rect 3718 2988 3722 2992
rect 3750 2988 3754 2992
rect 3950 2988 3954 2992
rect 3982 2988 3986 2992
rect 4022 2988 4026 2992
rect 4054 2988 4058 2992
rect 4238 2988 4242 2992
rect 4278 2988 4282 2992
rect 4814 2988 4818 2992
rect 4886 2988 4890 2992
rect 6 2978 10 2982
rect 798 2978 802 2982
rect 1798 2978 1802 2982
rect 4350 2978 4354 2982
rect 334 2968 338 2972
rect 390 2968 394 2972
rect 566 2968 570 2972
rect 1190 2968 1194 2972
rect 1478 2968 1482 2972
rect 1582 2968 1586 2972
rect 1654 2968 1658 2972
rect 1942 2968 1946 2972
rect 2166 2968 2170 2972
rect 3390 2968 3394 2972
rect 3686 2968 3690 2972
rect 3934 2968 3938 2972
rect 4134 2968 4138 2972
rect 4206 2968 4210 2972
rect 4222 2968 4226 2972
rect 4478 2968 4482 2972
rect 4710 2968 4714 2972
rect 4990 2968 4994 2972
rect 366 2958 370 2962
rect 70 2947 74 2951
rect 118 2948 122 2952
rect 150 2948 154 2952
rect 174 2948 178 2952
rect 206 2948 210 2952
rect 238 2948 242 2952
rect 278 2948 282 2952
rect 358 2948 362 2952
rect 494 2958 498 2962
rect 502 2958 506 2962
rect 518 2958 522 2962
rect 534 2958 538 2962
rect 734 2958 738 2962
rect 750 2958 754 2962
rect 758 2958 762 2962
rect 774 2958 778 2962
rect 806 2958 810 2962
rect 406 2948 410 2952
rect 430 2948 434 2952
rect 454 2948 458 2952
rect 462 2948 466 2952
rect 470 2948 474 2952
rect 518 2948 522 2952
rect 566 2948 570 2952
rect 582 2948 586 2952
rect 638 2948 642 2952
rect 670 2948 674 2952
rect 678 2948 682 2952
rect 686 2948 690 2952
rect 726 2948 730 2952
rect 734 2948 738 2952
rect 774 2948 778 2952
rect 814 2948 818 2952
rect 886 2948 890 2952
rect 910 2948 914 2952
rect 918 2948 922 2952
rect 942 2948 946 2952
rect 982 2948 986 2952
rect 1006 2948 1010 2952
rect 1014 2948 1018 2952
rect 1022 2948 1026 2952
rect 1046 2948 1050 2952
rect 1070 2948 1074 2952
rect 1110 2948 1114 2952
rect 1142 2948 1146 2952
rect 1158 2948 1162 2952
rect 1342 2958 1346 2962
rect 1358 2958 1362 2962
rect 1374 2958 1378 2962
rect 1678 2958 1682 2962
rect 1694 2958 1698 2962
rect 1814 2958 1818 2962
rect 1830 2958 1834 2962
rect 2030 2958 2034 2962
rect 2270 2958 2274 2962
rect 2294 2958 2298 2962
rect 2470 2958 2474 2962
rect 2486 2958 2490 2962
rect 2542 2958 2546 2962
rect 2558 2958 2562 2962
rect 2630 2958 2634 2962
rect 2686 2958 2690 2962
rect 2782 2958 2786 2962
rect 1246 2948 1250 2952
rect 1286 2948 1290 2952
rect 1326 2948 1330 2952
rect 1342 2948 1346 2952
rect 1358 2948 1362 2952
rect 86 2938 90 2942
rect 126 2938 130 2942
rect 142 2938 146 2942
rect 198 2938 202 2942
rect 214 2938 218 2942
rect 254 2938 258 2942
rect 358 2938 362 2942
rect 414 2938 418 2942
rect 470 2938 474 2942
rect 526 2938 530 2942
rect 574 2938 578 2942
rect 606 2938 610 2942
rect 662 2938 666 2942
rect 718 2938 722 2942
rect 782 2938 786 2942
rect 790 2938 794 2942
rect 838 2938 842 2942
rect 966 2938 970 2942
rect 974 2938 978 2942
rect 1118 2938 1122 2942
rect 1142 2938 1146 2942
rect 1182 2938 1186 2942
rect 1270 2938 1274 2942
rect 1318 2938 1322 2942
rect 1406 2947 1410 2951
rect 1534 2948 1538 2952
rect 1614 2948 1618 2952
rect 1678 2948 1682 2952
rect 1694 2948 1698 2952
rect 1710 2948 1714 2952
rect 1726 2948 1730 2952
rect 1782 2948 1786 2952
rect 1798 2948 1802 2952
rect 1830 2948 1834 2952
rect 1846 2948 1850 2952
rect 1350 2938 1354 2942
rect 1422 2938 1426 2942
rect 1606 2938 1610 2942
rect 1638 2938 1642 2942
rect 1686 2938 1690 2942
rect 1878 2947 1882 2951
rect 1998 2948 2002 2952
rect 2006 2948 2010 2952
rect 2038 2948 2042 2952
rect 2102 2947 2106 2951
rect 2134 2948 2138 2952
rect 2174 2948 2178 2952
rect 2182 2948 2186 2952
rect 2206 2948 2210 2952
rect 2222 2948 2226 2952
rect 2230 2948 2234 2952
rect 2262 2948 2266 2952
rect 2334 2948 2338 2952
rect 2382 2948 2386 2952
rect 2446 2948 2450 2952
rect 2462 2948 2466 2952
rect 2494 2948 2498 2952
rect 2502 2948 2506 2952
rect 2526 2948 2530 2952
rect 2614 2948 2618 2952
rect 2670 2948 2674 2952
rect 2678 2948 2682 2952
rect 2702 2948 2706 2952
rect 2726 2948 2730 2952
rect 2734 2948 2738 2952
rect 2750 2948 2754 2952
rect 2758 2948 2762 2952
rect 2934 2958 2938 2962
rect 3126 2958 3130 2962
rect 2798 2948 2802 2952
rect 2814 2948 2818 2952
rect 2830 2948 2834 2952
rect 2894 2948 2898 2952
rect 2958 2948 2962 2952
rect 2974 2948 2978 2952
rect 1718 2938 1722 2942
rect 1790 2938 1794 2942
rect 1822 2938 1826 2942
rect 1966 2938 1970 2942
rect 2014 2938 2018 2942
rect 2286 2938 2290 2942
rect 2310 2938 2314 2942
rect 2342 2938 2346 2942
rect 2374 2938 2378 2942
rect 2382 2938 2386 2942
rect 2542 2938 2546 2942
rect 2558 2938 2562 2942
rect 2582 2938 2586 2942
rect 2606 2938 2610 2942
rect 2694 2938 2698 2942
rect 2710 2938 2714 2942
rect 2766 2938 2770 2942
rect 3070 2947 3074 2951
rect 3126 2948 3130 2952
rect 3150 2958 3154 2962
rect 3550 2958 3554 2962
rect 3734 2958 3738 2962
rect 3790 2958 3794 2962
rect 3198 2948 3202 2952
rect 3214 2948 3218 2952
rect 3246 2948 3250 2952
rect 3254 2948 3258 2952
rect 3262 2948 3266 2952
rect 3286 2948 3290 2952
rect 3326 2947 3330 2951
rect 3430 2948 3434 2952
rect 3462 2947 3466 2951
rect 3518 2948 3522 2952
rect 3534 2948 3538 2952
rect 3542 2948 3546 2952
rect 3582 2947 3586 2951
rect 3718 2948 3722 2952
rect 3766 2948 3770 2952
rect 3814 2958 3818 2962
rect 3942 2958 3946 2962
rect 4574 2958 4578 2962
rect 3814 2948 3818 2952
rect 3870 2947 3874 2951
rect 3966 2948 3970 2952
rect 3974 2948 3978 2952
rect 3998 2948 4002 2952
rect 4038 2948 4042 2952
rect 4070 2948 4074 2952
rect 4102 2948 4106 2952
rect 4150 2948 4154 2952
rect 4254 2948 4258 2952
rect 4310 2948 4314 2952
rect 4326 2948 4330 2952
rect 4342 2948 4346 2952
rect 4406 2948 4410 2952
rect 4614 2958 4618 2962
rect 4702 2958 4706 2962
rect 4526 2947 4530 2951
rect 4598 2948 4602 2952
rect 4678 2948 4682 2952
rect 4766 2948 4770 2952
rect 4830 2948 4834 2952
rect 4838 2948 4842 2952
rect 4870 2948 4874 2952
rect 4902 2948 4906 2952
rect 4966 2958 4970 2962
rect 5070 2958 5074 2962
rect 5030 2948 5034 2952
rect 5086 2948 5090 2952
rect 5166 2948 5170 2952
rect 2870 2938 2874 2942
rect 2918 2938 2922 2942
rect 2950 2938 2954 2942
rect 2990 2938 2994 2942
rect 3054 2938 3058 2942
rect 3110 2938 3114 2942
rect 3166 2938 3170 2942
rect 3174 2938 3178 2942
rect 3190 2938 3194 2942
rect 3238 2938 3242 2942
rect 3494 2938 3498 2942
rect 3510 2938 3514 2942
rect 3526 2938 3530 2942
rect 3566 2938 3570 2942
rect 3614 2938 3618 2942
rect 3686 2938 3690 2942
rect 3702 2938 3706 2942
rect 3710 2938 3714 2942
rect 3774 2938 3778 2942
rect 3854 2938 3858 2942
rect 3958 2938 3962 2942
rect 4094 2938 4098 2942
rect 4110 2938 4114 2942
rect 4182 2938 4186 2942
rect 4206 2938 4210 2942
rect 4334 2938 4338 2942
rect 4382 2938 4386 2942
rect 4414 2938 4418 2942
rect 4542 2938 4546 2942
rect 4558 2938 4562 2942
rect 4582 2938 4586 2942
rect 4606 2938 4610 2942
rect 4630 2938 4634 2942
rect 4670 2938 4674 2942
rect 4686 2938 4690 2942
rect 4702 2938 4706 2942
rect 4790 2938 4794 2942
rect 4846 2938 4850 2942
rect 4902 2938 4906 2942
rect 102 2928 106 2932
rect 158 2928 162 2932
rect 342 2928 346 2932
rect 646 2928 650 2932
rect 654 2928 658 2932
rect 926 2928 930 2932
rect 1158 2928 1162 2932
rect 1478 2928 1482 2932
rect 1518 2928 1522 2932
rect 1878 2928 1882 2932
rect 2070 2928 2074 2932
rect 2238 2928 2242 2932
rect 3198 2928 3202 2932
rect 3326 2928 3330 2932
rect 3494 2928 3498 2932
rect 3838 2928 3842 2932
rect 4078 2928 4082 2932
rect 4294 2928 4298 2932
rect 4446 2928 4450 2932
rect 4654 2928 4658 2932
rect 4862 2928 4866 2932
rect 4942 2938 4946 2942
rect 4950 2938 4954 2942
rect 5054 2938 5058 2942
rect 5086 2938 5090 2942
rect 5158 2938 5162 2942
rect 5174 2938 5178 2942
rect 4918 2928 4922 2932
rect 5190 2928 5194 2932
rect 190 2918 194 2922
rect 350 2918 354 2922
rect 446 2918 450 2922
rect 494 2918 498 2922
rect 598 2918 602 2922
rect 702 2918 706 2922
rect 862 2918 866 2922
rect 958 2918 962 2922
rect 1094 2918 1098 2922
rect 1174 2918 1178 2922
rect 1302 2918 1306 2922
rect 1630 2918 1634 2922
rect 1742 2918 1746 2922
rect 1958 2918 1962 2922
rect 2190 2918 2194 2922
rect 2318 2918 2322 2922
rect 2518 2918 2522 2922
rect 2574 2918 2578 2922
rect 2654 2918 2658 2922
rect 3230 2918 3234 2922
rect 3278 2918 3282 2922
rect 3398 2918 3402 2922
rect 3686 2918 3690 2922
rect 3750 2918 3754 2922
rect 3830 2918 3834 2922
rect 4086 2918 4090 2922
rect 4118 2918 4122 2922
rect 4166 2918 4170 2922
rect 4198 2918 4202 2922
rect 4214 2918 4218 2922
rect 4614 2918 4618 2922
rect 4662 2918 4666 2922
rect 4854 2918 4858 2922
rect 4886 2918 4890 2922
rect 4934 2918 4938 2922
rect 4958 2918 4962 2922
rect 4974 2918 4978 2922
rect 5078 2918 5082 2922
rect 5182 2918 5186 2922
rect 1050 2903 1054 2907
rect 1057 2903 1061 2907
rect 2074 2903 2078 2907
rect 2081 2903 2085 2907
rect 3098 2903 3102 2907
rect 3105 2903 3109 2907
rect 4114 2903 4118 2907
rect 4121 2903 4125 2907
rect 6 2888 10 2892
rect 238 2888 242 2892
rect 334 2888 338 2892
rect 510 2888 514 2892
rect 638 2888 642 2892
rect 654 2888 658 2892
rect 678 2888 682 2892
rect 806 2888 810 2892
rect 998 2888 1002 2892
rect 1446 2888 1450 2892
rect 1910 2888 1914 2892
rect 2014 2888 2018 2892
rect 2078 2888 2082 2892
rect 2158 2888 2162 2892
rect 2278 2888 2282 2892
rect 2318 2888 2322 2892
rect 3030 2888 3034 2892
rect 3070 2888 3074 2892
rect 3350 2888 3354 2892
rect 3470 2888 3474 2892
rect 3534 2888 3538 2892
rect 3550 2888 3554 2892
rect 3598 2888 3602 2892
rect 3758 2888 3762 2892
rect 3918 2888 3922 2892
rect 4022 2888 4026 2892
rect 4182 2888 4186 2892
rect 4246 2888 4250 2892
rect 4302 2888 4306 2892
rect 4406 2888 4410 2892
rect 4678 2888 4682 2892
rect 4718 2888 4722 2892
rect 4774 2888 4778 2892
rect 4918 2888 4922 2892
rect 5038 2888 5042 2892
rect 5086 2888 5090 2892
rect 398 2878 402 2882
rect 414 2878 418 2882
rect 646 2878 650 2882
rect 670 2878 674 2882
rect 1102 2878 1106 2882
rect 1222 2878 1226 2882
rect 2094 2878 2098 2882
rect 2302 2878 2306 2882
rect 2382 2878 2386 2882
rect 3038 2878 3042 2882
rect 3078 2878 3082 2882
rect 3462 2878 3466 2882
rect 3646 2878 3650 2882
rect 4190 2878 4194 2882
rect 4286 2878 4290 2882
rect 4686 2878 4690 2882
rect 4750 2878 4754 2882
rect 4758 2878 4762 2882
rect 5046 2878 5050 2882
rect 5118 2878 5122 2882
rect 86 2868 90 2872
rect 158 2868 162 2872
rect 254 2868 258 2872
rect 342 2868 346 2872
rect 358 2868 362 2872
rect 390 2868 394 2872
rect 430 2868 434 2872
rect 558 2868 562 2872
rect 734 2868 738 2872
rect 766 2868 770 2872
rect 870 2868 874 2872
rect 942 2868 946 2872
rect 990 2868 994 2872
rect 1166 2868 1170 2872
rect 1190 2868 1194 2872
rect 1294 2868 1298 2872
rect 1310 2868 1314 2872
rect 1350 2868 1354 2872
rect 1382 2868 1386 2872
rect 1454 2868 1458 2872
rect 1510 2868 1514 2872
rect 1534 2868 1538 2872
rect 1542 2868 1546 2872
rect 1574 2868 1578 2872
rect 1686 2868 1690 2872
rect 1742 2868 1746 2872
rect 1830 2868 1834 2872
rect 1950 2868 1954 2872
rect 2038 2868 2042 2872
rect 2134 2868 2138 2872
rect 2150 2868 2154 2872
rect 2238 2868 2242 2872
rect 2310 2868 2314 2872
rect 70 2859 74 2863
rect 102 2858 106 2862
rect 110 2858 114 2862
rect 134 2858 138 2862
rect 182 2858 186 2862
rect 278 2858 282 2862
rect 350 2858 354 2862
rect 414 2858 418 2862
rect 454 2858 458 2862
rect 534 2858 538 2862
rect 582 2858 586 2862
rect 662 2858 666 2862
rect 694 2858 698 2862
rect 702 2858 706 2862
rect 758 2858 762 2862
rect 774 2858 778 2862
rect 862 2858 866 2862
rect 902 2858 906 2862
rect 910 2858 914 2862
rect 934 2858 938 2862
rect 950 2858 954 2862
rect 982 2858 986 2862
rect 1014 2858 1018 2862
rect 1030 2858 1034 2862
rect 1054 2858 1058 2862
rect 1062 2858 1066 2862
rect 1070 2858 1074 2862
rect 1094 2858 1098 2862
rect 1118 2858 1122 2862
rect 1158 2858 1162 2862
rect 1182 2858 1186 2862
rect 1230 2858 1234 2862
rect 1302 2858 1306 2862
rect 1342 2858 1346 2862
rect 1390 2858 1394 2862
rect 1462 2858 1466 2862
rect 1502 2858 1506 2862
rect 1534 2858 1538 2862
rect 1550 2858 1554 2862
rect 1590 2858 1594 2862
rect 1598 2858 1602 2862
rect 1622 2858 1626 2862
rect 1638 2858 1642 2862
rect 1646 2858 1650 2862
rect 1670 2858 1674 2862
rect 1678 2858 1682 2862
rect 1734 2858 1738 2862
rect 1798 2858 1802 2862
rect 1846 2858 1850 2862
rect 1854 2858 1858 2862
rect 1878 2858 1882 2862
rect 1894 2858 1898 2862
rect 1918 2858 1922 2862
rect 1942 2858 1946 2862
rect 1958 2858 1962 2862
rect 1990 2858 1994 2862
rect 1998 2858 2002 2862
rect 2030 2858 2034 2862
rect 2046 2858 2050 2862
rect 2110 2858 2114 2862
rect 2214 2858 2218 2862
rect 2254 2858 2258 2862
rect 2286 2858 2290 2862
rect 2302 2858 2306 2862
rect 2350 2858 2354 2862
rect 2382 2859 2386 2863
rect 2462 2868 2466 2872
rect 2486 2868 2490 2872
rect 2518 2868 2522 2872
rect 2678 2868 2682 2872
rect 2766 2868 2770 2872
rect 2414 2858 2418 2862
rect 2422 2858 2426 2862
rect 2486 2858 2490 2862
rect 2510 2858 2514 2862
rect 2526 2858 2530 2862
rect 2534 2858 2538 2862
rect 2558 2858 2562 2862
rect 2598 2858 2602 2862
rect 2622 2858 2626 2862
rect 2630 2858 2634 2862
rect 2654 2858 2658 2862
rect 2750 2859 2754 2863
rect 2830 2868 2834 2872
rect 2838 2868 2842 2872
rect 2894 2868 2898 2872
rect 2918 2868 2922 2872
rect 2982 2868 2986 2872
rect 3206 2868 3210 2872
rect 3262 2868 3266 2872
rect 3310 2868 3314 2872
rect 3334 2868 3338 2872
rect 3342 2868 3346 2872
rect 3566 2868 3570 2872
rect 3574 2868 3578 2872
rect 3702 2868 3706 2872
rect 3886 2868 3890 2872
rect 3902 2868 3906 2872
rect 3926 2868 3930 2872
rect 4006 2868 4010 2872
rect 4022 2868 4026 2872
rect 4078 2868 4082 2872
rect 4150 2868 4154 2872
rect 4158 2868 4162 2872
rect 4222 2868 4226 2872
rect 4230 2868 4234 2872
rect 4294 2868 4298 2872
rect 4382 2868 4386 2872
rect 4430 2868 4434 2872
rect 4446 2868 4450 2872
rect 4606 2868 4610 2872
rect 4670 2868 4674 2872
rect 4742 2868 4746 2872
rect 4798 2868 4802 2872
rect 5022 2868 5026 2872
rect 5134 2868 5138 2872
rect 5182 2868 5186 2872
rect 2782 2858 2786 2862
rect 2790 2858 2794 2862
rect 2846 2858 2850 2862
rect 2886 2858 2890 2862
rect 2902 2858 2906 2862
rect 2942 2858 2946 2862
rect 2966 2858 2970 2862
rect 2974 2858 2978 2862
rect 2990 2858 2994 2862
rect 3014 2858 3018 2862
rect 3022 2858 3026 2862
rect 3046 2858 3050 2862
rect 3142 2858 3146 2862
rect 3166 2858 3170 2862
rect 3214 2858 3218 2862
rect 3230 2858 3234 2862
rect 3270 2858 3274 2862
rect 3278 2858 3282 2862
rect 3310 2858 3314 2862
rect 3366 2858 3370 2862
rect 3374 2858 3378 2862
rect 3398 2858 3402 2862
rect 3422 2858 3426 2862
rect 3446 2858 3450 2862
rect 3454 2858 3458 2862
rect 3478 2858 3482 2862
rect 3510 2858 3514 2862
rect 3518 2858 3522 2862
rect 3630 2858 3634 2862
rect 3638 2858 3642 2862
rect 3694 2858 3698 2862
rect 3742 2858 3746 2862
rect 3798 2858 3802 2862
rect 3838 2858 3842 2862
rect 3870 2858 3874 2862
rect 3926 2858 3930 2862
rect 3966 2858 3970 2862
rect 3990 2858 3994 2862
rect 3998 2858 4002 2862
rect 4038 2858 4042 2862
rect 4062 2858 4066 2862
rect 4070 2858 4074 2862
rect 4086 2858 4090 2862
rect 4110 2858 4114 2862
rect 4142 2858 4146 2862
rect 4214 2858 4218 2862
rect 4262 2858 4266 2862
rect 4270 2858 4274 2862
rect 4358 2858 4362 2862
rect 4422 2858 4426 2862
rect 4438 2858 4442 2862
rect 4462 2858 4466 2862
rect 4470 2858 4474 2862
rect 4494 2858 4498 2862
rect 4510 2858 4514 2862
rect 4518 2858 4522 2862
rect 4542 2858 4546 2862
rect 4566 2858 4570 2862
rect 4590 2858 4594 2862
rect 4598 2858 4602 2862
rect 4662 2858 4666 2862
rect 4702 2858 4706 2862
rect 4790 2858 4794 2862
rect 4806 2858 4810 2862
rect 4814 2858 4818 2862
rect 4854 2859 4858 2863
rect 4886 2858 4890 2862
rect 4982 2858 4986 2862
rect 5062 2858 5066 2862
rect 5070 2858 5074 2862
rect 5134 2858 5138 2862
rect 374 2848 378 2852
rect 718 2848 722 2852
rect 742 2848 746 2852
rect 926 2848 930 2852
rect 1166 2848 1170 2852
rect 1462 2848 1466 2852
rect 1486 2848 1490 2852
rect 1518 2848 1522 2852
rect 1566 2848 1570 2852
rect 1926 2848 1930 2852
rect 2062 2848 2066 2852
rect 2134 2848 2138 2852
rect 2422 2848 2426 2852
rect 2446 2848 2450 2852
rect 2470 2848 2474 2852
rect 2638 2848 2642 2852
rect 2654 2848 2658 2852
rect 2814 2848 2818 2852
rect 3070 2848 3074 2852
rect 3214 2848 3218 2852
rect 3230 2848 3234 2852
rect 3318 2848 3322 2852
rect 3358 2848 3362 2852
rect 3550 2848 3554 2852
rect 3678 2848 3682 2852
rect 3718 2848 3722 2852
rect 3782 2848 3786 2852
rect 3918 2848 3922 2852
rect 3950 2848 3954 2852
rect 4022 2848 4026 2852
rect 4102 2848 4106 2852
rect 4126 2848 4130 2852
rect 4158 2848 4162 2852
rect 4174 2848 4178 2852
rect 4198 2848 4202 2852
rect 4246 2848 4250 2852
rect 4254 2848 4258 2852
rect 4454 2848 4458 2852
rect 4638 2848 4642 2852
rect 4726 2848 4730 2852
rect 4822 2848 4826 2852
rect 5078 2848 5082 2852
rect 494 2838 498 2842
rect 1142 2838 1146 2842
rect 1270 2838 1274 2842
rect 1286 2838 1290 2842
rect 1326 2838 1330 2842
rect 1710 2838 1714 2842
rect 1750 2838 1754 2842
rect 1910 2838 1914 2842
rect 2702 2838 2706 2842
rect 2790 2838 2794 2842
rect 2870 2838 2874 2842
rect 3110 2838 3114 2842
rect 3814 2838 3818 2842
rect 4214 2838 4218 2842
rect 3382 2828 3386 2832
rect 3934 2828 3938 2832
rect 126 2818 130 2822
rect 758 2818 762 2822
rect 790 2818 794 2822
rect 958 2818 962 2822
rect 998 2818 1002 2822
rect 1046 2818 1050 2822
rect 1614 2818 1618 2822
rect 1662 2818 1666 2822
rect 1734 2818 1738 2822
rect 1862 2818 1866 2822
rect 1974 2818 1978 2822
rect 2046 2818 2050 2822
rect 2542 2818 2546 2822
rect 2606 2818 2610 2822
rect 2846 2818 2850 2822
rect 2958 2818 2962 2822
rect 3086 2818 3090 2822
rect 3286 2818 3290 2822
rect 3430 2818 3434 2822
rect 3494 2818 3498 2822
rect 3854 2818 3858 2822
rect 3974 2818 3978 2822
rect 4086 2818 4090 2822
rect 4478 2818 4482 2822
rect 4526 2818 4530 2822
rect 4574 2818 4578 2822
rect 4662 2818 4666 2822
rect 4926 2818 4930 2822
rect 538 2803 542 2807
rect 545 2803 549 2807
rect 1562 2803 1566 2807
rect 1569 2803 1573 2807
rect 2586 2803 2590 2807
rect 2593 2803 2597 2807
rect 3610 2803 3614 2807
rect 3617 2803 3621 2807
rect 4634 2803 4638 2807
rect 4641 2803 4645 2807
rect 606 2788 610 2792
rect 934 2788 938 2792
rect 966 2788 970 2792
rect 1502 2788 1506 2792
rect 1718 2788 1722 2792
rect 2054 2788 2058 2792
rect 2502 2788 2506 2792
rect 2518 2788 2522 2792
rect 2622 2788 2626 2792
rect 3094 2788 3098 2792
rect 3166 2788 3170 2792
rect 3190 2788 3194 2792
rect 3278 2788 3282 2792
rect 3350 2788 3354 2792
rect 3446 2788 3450 2792
rect 3478 2788 3482 2792
rect 3510 2788 3514 2792
rect 3902 2788 3906 2792
rect 4230 2788 4234 2792
rect 4382 2788 4386 2792
rect 4654 2788 4658 2792
rect 4742 2788 4746 2792
rect 4846 2788 4850 2792
rect 4878 2788 4882 2792
rect 4910 2788 4914 2792
rect 4942 2788 4946 2792
rect 4974 2788 4978 2792
rect 5102 2788 5106 2792
rect 5182 2788 5186 2792
rect 222 2768 226 2772
rect 238 2768 242 2772
rect 2254 2768 2258 2772
rect 2758 2768 2762 2772
rect 3574 2768 3578 2772
rect 3622 2768 3626 2772
rect 3662 2768 3666 2772
rect 3734 2768 3738 2772
rect 4014 2768 4018 2772
rect 366 2758 370 2762
rect 486 2758 490 2762
rect 542 2758 546 2762
rect 798 2758 802 2762
rect 1238 2758 1242 2762
rect 134 2748 138 2752
rect 182 2748 186 2752
rect 246 2748 250 2752
rect 294 2747 298 2751
rect 326 2748 330 2752
rect 422 2748 426 2752
rect 502 2748 506 2752
rect 518 2748 522 2752
rect 558 2748 562 2752
rect 662 2748 666 2752
rect 742 2748 746 2752
rect 822 2748 826 2752
rect 870 2748 874 2752
rect 950 2748 954 2752
rect 1102 2748 1106 2752
rect 1166 2748 1170 2752
rect 1214 2748 1218 2752
rect 1262 2758 1266 2762
rect 1390 2758 1394 2762
rect 1462 2758 1466 2762
rect 1262 2748 1266 2752
rect 1350 2748 1354 2752
rect 1438 2748 1442 2752
rect 1486 2758 1490 2762
rect 1686 2758 1690 2762
rect 1790 2758 1794 2762
rect 1486 2748 1490 2752
rect 1566 2748 1570 2752
rect 1590 2748 1594 2752
rect 1630 2748 1634 2752
rect 1662 2748 1666 2752
rect 1734 2748 1738 2752
rect 1742 2748 1746 2752
rect 1750 2748 1754 2752
rect 1774 2748 1778 2752
rect 1790 2748 1794 2752
rect 1814 2748 1818 2752
rect 1822 2748 1826 2752
rect 1846 2748 1850 2752
rect 1854 2748 1858 2752
rect 1886 2748 1890 2752
rect 6 2738 10 2742
rect 78 2738 82 2742
rect 158 2738 162 2742
rect 382 2738 386 2742
rect 398 2738 402 2742
rect 550 2738 554 2742
rect 582 2738 586 2742
rect 654 2738 658 2742
rect 710 2738 714 2742
rect 814 2738 818 2742
rect 822 2738 826 2742
rect 878 2738 882 2742
rect 982 2738 986 2742
rect 1054 2738 1058 2742
rect 1078 2738 1082 2742
rect 1174 2738 1178 2742
rect 1182 2738 1186 2742
rect 1222 2738 1226 2742
rect 1342 2738 1346 2742
rect 1406 2738 1410 2742
rect 1414 2738 1418 2742
rect 1446 2738 1450 2742
rect 1614 2738 1618 2742
rect 1638 2738 1642 2742
rect 1702 2738 1706 2742
rect 1918 2747 1922 2751
rect 1990 2748 1994 2752
rect 2006 2748 2010 2752
rect 2030 2758 2034 2762
rect 2134 2758 2138 2762
rect 2038 2748 2042 2752
rect 2086 2748 2090 2752
rect 2094 2748 2098 2752
rect 2150 2748 2154 2752
rect 2206 2748 2210 2752
rect 2230 2758 2234 2762
rect 2582 2758 2586 2762
rect 2774 2758 2778 2762
rect 2310 2748 2314 2752
rect 2350 2748 2354 2752
rect 2358 2748 2362 2752
rect 2382 2748 2386 2752
rect 2430 2748 2434 2752
rect 2446 2748 2450 2752
rect 2534 2748 2538 2752
rect 2566 2748 2570 2752
rect 2606 2748 2610 2752
rect 2638 2748 2642 2752
rect 2710 2748 2714 2752
rect 2774 2748 2778 2752
rect 2798 2758 2802 2762
rect 2830 2758 2834 2762
rect 2878 2758 2882 2762
rect 2894 2758 2898 2762
rect 3086 2758 3090 2762
rect 3142 2758 3146 2762
rect 2814 2748 2818 2752
rect 2846 2748 2850 2752
rect 2878 2748 2882 2752
rect 2966 2748 2970 2752
rect 3550 2758 3554 2762
rect 3830 2758 3834 2762
rect 3862 2758 3866 2762
rect 3942 2758 3946 2762
rect 3974 2758 3978 2762
rect 3166 2748 3170 2752
rect 3222 2748 3226 2752
rect 3254 2748 3258 2752
rect 3262 2748 3266 2752
rect 3494 2748 3498 2752
rect 3526 2748 3530 2752
rect 3534 2748 3538 2752
rect 3590 2748 3594 2752
rect 3622 2748 3626 2752
rect 3662 2748 3666 2752
rect 3694 2748 3698 2752
rect 1806 2738 1810 2742
rect 1862 2738 1866 2742
rect 1870 2738 1874 2742
rect 2030 2738 2034 2742
rect 2118 2738 2122 2742
rect 2158 2738 2162 2742
rect 2174 2738 2178 2742
rect 2230 2738 2234 2742
rect 2246 2738 2250 2742
rect 2334 2738 2338 2742
rect 2390 2738 2394 2742
rect 2662 2738 2666 2742
rect 2702 2738 2706 2742
rect 2766 2738 2770 2742
rect 2822 2738 2826 2742
rect 2846 2738 2850 2742
rect 2854 2738 2858 2742
rect 2886 2738 2890 2742
rect 2998 2738 3002 2742
rect 3014 2738 3018 2742
rect 3078 2738 3082 2742
rect 3118 2738 3122 2742
rect 3126 2738 3130 2742
rect 3798 2747 3802 2751
rect 3846 2748 3850 2752
rect 3878 2748 3882 2752
rect 3886 2748 3890 2752
rect 3902 2748 3906 2752
rect 3942 2748 3946 2752
rect 4534 2758 4538 2762
rect 4614 2758 4618 2762
rect 4862 2758 4866 2762
rect 4926 2758 4930 2762
rect 4990 2758 4994 2762
rect 3998 2748 4002 2752
rect 4062 2748 4066 2752
rect 4126 2748 4130 2752
rect 4134 2748 4138 2752
rect 4182 2748 4186 2752
rect 4206 2748 4210 2752
rect 4214 2748 4218 2752
rect 4230 2748 4234 2752
rect 3294 2738 3298 2742
rect 3366 2738 3370 2742
rect 3430 2738 3434 2742
rect 3470 2738 3474 2742
rect 3598 2738 3602 2742
rect 3646 2738 3650 2742
rect 3726 2738 3730 2742
rect 3798 2738 3802 2742
rect 3838 2738 3842 2742
rect 3854 2738 3858 2742
rect 3886 2738 3890 2742
rect 3926 2738 3930 2742
rect 3950 2738 3954 2742
rect 3990 2738 3994 2742
rect 4006 2738 4010 2742
rect 4342 2747 4346 2751
rect 4398 2748 4402 2752
rect 4462 2747 4466 2751
rect 4590 2748 4594 2752
rect 4646 2748 4650 2752
rect 4670 2748 4674 2752
rect 4678 2748 4682 2752
rect 4686 2748 4690 2752
rect 4734 2748 4738 2752
rect 4798 2748 4802 2752
rect 4838 2748 4842 2752
rect 4894 2748 4898 2752
rect 4910 2748 4914 2752
rect 4958 2748 4962 2752
rect 4974 2748 4978 2752
rect 5022 2747 5026 2751
rect 5054 2748 5058 2752
rect 5118 2748 5122 2752
rect 4222 2738 4226 2742
rect 4254 2738 4258 2742
rect 4326 2738 4330 2742
rect 4374 2738 4378 2742
rect 4446 2738 4450 2742
rect 4542 2738 4546 2742
rect 4558 2738 4562 2742
rect 4582 2738 4586 2742
rect 4598 2738 4602 2742
rect 4614 2738 4618 2742
rect 4726 2738 4730 2742
rect 4822 2738 4826 2742
rect 4838 2738 4842 2742
rect 4902 2738 4906 2742
rect 4966 2738 4970 2742
rect 5126 2738 5130 2742
rect 262 2728 266 2732
rect 574 2728 578 2732
rect 846 2728 850 2732
rect 854 2728 858 2732
rect 870 2728 874 2732
rect 1198 2728 1202 2732
rect 1678 2728 1682 2732
rect 1886 2728 1890 2732
rect 1918 2728 1922 2732
rect 1990 2728 1994 2732
rect 2006 2728 2010 2732
rect 2182 2728 2186 2732
rect 2190 2728 2194 2732
rect 2542 2728 2546 2732
rect 2878 2728 2882 2732
rect 2934 2728 2938 2732
rect 3182 2728 3186 2732
rect 3862 2728 3866 2732
rect 4078 2728 4082 2732
rect 4294 2728 4298 2732
rect 4566 2728 4570 2732
rect 4702 2728 4706 2732
rect 62 2718 66 2722
rect 254 2718 258 2722
rect 358 2718 362 2722
rect 374 2718 378 2722
rect 798 2718 802 2722
rect 838 2718 842 2722
rect 1158 2718 1162 2722
rect 1278 2718 1282 2722
rect 1398 2718 1402 2722
rect 1646 2718 1650 2722
rect 1694 2718 1698 2722
rect 1798 2718 1802 2722
rect 1982 2718 1986 2722
rect 2166 2718 2170 2722
rect 2366 2718 2370 2722
rect 2590 2718 2594 2722
rect 2838 2718 2842 2722
rect 3206 2718 3210 2722
rect 3478 2718 3482 2722
rect 3686 2718 3690 2722
rect 4142 2718 4146 2722
rect 4382 2718 4386 2722
rect 4422 2718 4426 2722
rect 4526 2718 4530 2722
rect 4718 2718 4722 2722
rect 4878 2718 4882 2722
rect 4942 2718 4946 2722
rect 5086 2718 5090 2722
rect 5102 2718 5106 2722
rect 1050 2703 1054 2707
rect 1057 2703 1061 2707
rect 2074 2703 2078 2707
rect 2081 2703 2085 2707
rect 3098 2703 3102 2707
rect 3105 2703 3109 2707
rect 4114 2703 4118 2707
rect 4121 2703 4125 2707
rect 246 2688 250 2692
rect 278 2688 282 2692
rect 542 2688 546 2692
rect 582 2688 586 2692
rect 702 2688 706 2692
rect 1678 2688 1682 2692
rect 1710 2688 1714 2692
rect 1942 2688 1946 2692
rect 2110 2688 2114 2692
rect 2206 2688 2210 2692
rect 2294 2688 2298 2692
rect 2526 2688 2530 2692
rect 2534 2688 2538 2692
rect 2566 2688 2570 2692
rect 2686 2688 2690 2692
rect 2822 2688 2826 2692
rect 2950 2688 2954 2692
rect 3062 2688 3066 2692
rect 3150 2688 3154 2692
rect 3798 2688 3802 2692
rect 3926 2688 3930 2692
rect 3950 2688 3954 2692
rect 4198 2688 4202 2692
rect 4254 2688 4258 2692
rect 4350 2688 4354 2692
rect 4422 2688 4426 2692
rect 4462 2688 4466 2692
rect 4582 2688 4586 2692
rect 4606 2688 4610 2692
rect 4926 2688 4930 2692
rect 4982 2688 4986 2692
rect 4990 2688 4994 2692
rect 5166 2688 5170 2692
rect 102 2678 106 2682
rect 198 2678 202 2682
rect 254 2678 258 2682
rect 310 2678 314 2682
rect 318 2678 322 2682
rect 398 2678 402 2682
rect 646 2678 650 2682
rect 726 2678 730 2682
rect 870 2678 874 2682
rect 950 2678 954 2682
rect 1102 2678 1106 2682
rect 1406 2678 1410 2682
rect 1470 2678 1474 2682
rect 1494 2678 1498 2682
rect 1526 2678 1530 2682
rect 1614 2678 1618 2682
rect 1766 2678 1770 2682
rect 2078 2678 2082 2682
rect 2246 2678 2250 2682
rect 2262 2678 2266 2682
rect 2918 2678 2922 2682
rect 2934 2678 2938 2682
rect 2998 2678 3002 2682
rect 3134 2678 3138 2682
rect 3198 2678 3202 2682
rect 3430 2678 3434 2682
rect 3742 2678 3746 2682
rect 3910 2678 3914 2682
rect 126 2668 130 2672
rect 142 2668 146 2672
rect 238 2668 242 2672
rect 270 2668 274 2672
rect 358 2668 362 2672
rect 518 2668 522 2672
rect 534 2668 538 2672
rect 574 2668 578 2672
rect 662 2668 666 2672
rect 806 2668 810 2672
rect 838 2668 842 2672
rect 966 2668 970 2672
rect 982 2668 986 2672
rect 1030 2668 1034 2672
rect 1062 2668 1066 2672
rect 1086 2668 1090 2672
rect 1118 2668 1122 2672
rect 1222 2668 1226 2672
rect 1254 2668 1258 2672
rect 1286 2668 1290 2672
rect 1366 2668 1370 2672
rect 1422 2668 1426 2672
rect 1550 2668 1554 2672
rect 1566 2668 1570 2672
rect 1686 2668 1690 2672
rect 1822 2668 1826 2672
rect 1894 2668 1898 2672
rect 1950 2668 1954 2672
rect 2022 2668 2026 2672
rect 2038 2668 2042 2672
rect 2062 2668 2066 2672
rect 2102 2668 2106 2672
rect 2190 2668 2194 2672
rect 2222 2668 2226 2672
rect 2270 2668 2274 2672
rect 2294 2668 2298 2672
rect 2366 2668 2370 2672
rect 2374 2668 2378 2672
rect 2430 2668 2434 2672
rect 2446 2668 2450 2672
rect 2550 2668 2554 2672
rect 2726 2668 2730 2672
rect 38 2658 42 2662
rect 62 2658 66 2662
rect 118 2658 122 2662
rect 150 2658 154 2662
rect 182 2658 186 2662
rect 190 2658 194 2662
rect 214 2658 218 2662
rect 222 2658 226 2662
rect 230 2658 234 2662
rect 262 2658 266 2662
rect 294 2658 298 2662
rect 334 2658 338 2662
rect 366 2658 370 2662
rect 406 2658 410 2662
rect 494 2658 498 2662
rect 646 2659 650 2663
rect 686 2658 690 2662
rect 710 2658 714 2662
rect 718 2658 722 2662
rect 798 2658 802 2662
rect 846 2658 850 2662
rect 950 2659 954 2663
rect 990 2658 994 2662
rect 1046 2658 1050 2662
rect 1086 2658 1090 2662
rect 1134 2659 1138 2663
rect 1238 2658 1242 2662
rect 1246 2658 1250 2662
rect 1294 2658 1298 2662
rect 1382 2658 1386 2662
rect 1446 2658 1450 2662
rect 1478 2658 1482 2662
rect 1510 2658 1514 2662
rect 1534 2658 1538 2662
rect 1542 2658 1546 2662
rect 1638 2658 1642 2662
rect 1686 2658 1690 2662
rect 1718 2658 1722 2662
rect 1726 2658 1730 2662
rect 1750 2658 1754 2662
rect 1782 2658 1786 2662
rect 1854 2658 1858 2662
rect 1926 2658 1930 2662
rect 1958 2658 1962 2662
rect 1966 2658 1970 2662
rect 1974 2658 1978 2662
rect 1998 2658 2002 2662
rect 2014 2658 2018 2662
rect 2046 2658 2050 2662
rect 2158 2658 2162 2662
rect 2382 2658 2386 2662
rect 2414 2658 2418 2662
rect 2422 2658 2426 2662
rect 2462 2659 2466 2663
rect 2854 2668 2858 2672
rect 2862 2668 2866 2672
rect 2902 2668 2906 2672
rect 3070 2668 3074 2672
rect 3086 2668 3090 2672
rect 3302 2668 3306 2672
rect 3334 2668 3338 2672
rect 3366 2668 3370 2672
rect 3398 2668 3402 2672
rect 3606 2668 3610 2672
rect 3646 2668 3650 2672
rect 3694 2668 3698 2672
rect 3718 2668 3722 2672
rect 3782 2668 3786 2672
rect 3862 2668 3866 2672
rect 4046 2678 4050 2682
rect 4230 2678 4234 2682
rect 4318 2678 4322 2682
rect 4534 2678 4538 2682
rect 4590 2678 4594 2682
rect 5062 2678 5066 2682
rect 3934 2668 3938 2672
rect 4014 2668 4018 2672
rect 4030 2668 4034 2672
rect 4086 2668 4090 2672
rect 4310 2668 4314 2672
rect 4358 2668 4362 2672
rect 4438 2668 4442 2672
rect 2494 2658 2498 2662
rect 2598 2658 2602 2662
rect 2662 2658 2666 2662
rect 2702 2658 2706 2662
rect 2766 2658 2770 2662
rect 2790 2658 2794 2662
rect 2830 2658 2834 2662
rect 2846 2658 2850 2662
rect 2862 2658 2866 2662
rect 2894 2658 2898 2662
rect 2910 2658 2914 2662
rect 2934 2658 2938 2662
rect 2966 2658 2970 2662
rect 3022 2658 3026 2662
rect 3110 2658 3114 2662
rect 3166 2658 3170 2662
rect 3214 2658 3218 2662
rect 3294 2658 3298 2662
rect 3374 2658 3378 2662
rect 3390 2658 3394 2662
rect 3430 2659 3434 2663
rect 4494 2668 4498 2672
rect 4526 2668 4530 2672
rect 4590 2668 4594 2672
rect 4662 2668 4666 2672
rect 4670 2668 4674 2672
rect 4702 2668 4706 2672
rect 4774 2668 4778 2672
rect 4870 2668 4874 2672
rect 4918 2668 4922 2672
rect 4942 2668 4946 2672
rect 4966 2668 4970 2672
rect 5022 2668 5026 2672
rect 5062 2668 5066 2672
rect 5070 2668 5074 2672
rect 5086 2668 5090 2672
rect 5158 2678 5162 2682
rect 5134 2668 5138 2672
rect 5182 2668 5186 2672
rect 3518 2658 3522 2662
rect 3542 2658 3546 2662
rect 3558 2658 3562 2662
rect 3582 2658 3586 2662
rect 3590 2658 3594 2662
rect 3598 2658 3602 2662
rect 3678 2658 3682 2662
rect 3686 2658 3690 2662
rect 3758 2658 3762 2662
rect 3774 2658 3778 2662
rect 3790 2658 3794 2662
rect 3854 2658 3858 2662
rect 3894 2658 3898 2662
rect 3942 2658 3946 2662
rect 3998 2658 4002 2662
rect 4062 2658 4066 2662
rect 4094 2658 4098 2662
rect 4134 2658 4138 2662
rect 4166 2658 4170 2662
rect 4182 2658 4186 2662
rect 4206 2658 4210 2662
rect 4334 2658 4338 2662
rect 4366 2658 4370 2662
rect 4398 2658 4402 2662
rect 4406 2658 4410 2662
rect 4478 2658 4482 2662
rect 4486 2658 4490 2662
rect 4518 2658 4522 2662
rect 4566 2658 4570 2662
rect 4574 2658 4578 2662
rect 4622 2658 4626 2662
rect 4662 2658 4666 2662
rect 4670 2658 4674 2662
rect 4734 2658 4738 2662
rect 4750 2658 4754 2662
rect 4790 2658 4794 2662
rect 4862 2658 4866 2662
rect 4966 2658 4970 2662
rect 5006 2658 5010 2662
rect 5030 2658 5034 2662
rect 5110 2658 5114 2662
rect 5142 2658 5146 2662
rect 518 2648 522 2652
rect 558 2648 562 2652
rect 846 2648 850 2652
rect 862 2648 866 2652
rect 990 2648 994 2652
rect 1014 2648 1018 2652
rect 1206 2648 1210 2652
rect 1382 2648 1386 2652
rect 1398 2648 1402 2652
rect 1550 2648 1554 2652
rect 1710 2648 1714 2652
rect 1806 2648 1810 2652
rect 2078 2648 2082 2652
rect 2254 2648 2258 2652
rect 2294 2648 2298 2652
rect 2398 2648 2402 2652
rect 2830 2648 2834 2652
rect 2886 2648 2890 2652
rect 3086 2648 3090 2652
rect 3318 2648 3322 2652
rect 3334 2648 3338 2652
rect 3374 2648 3378 2652
rect 3390 2648 3394 2652
rect 3638 2648 3642 2652
rect 3710 2648 3714 2652
rect 3734 2648 3738 2652
rect 4142 2648 4146 2652
rect 4174 2648 4178 2652
rect 4454 2648 4458 2652
rect 4614 2648 4618 2652
rect 4638 2648 4642 2652
rect 4934 2648 4938 2652
rect 4958 2648 4962 2652
rect 4982 2648 4986 2652
rect 4990 2648 4994 2652
rect 5030 2648 5034 2652
rect 5046 2648 5050 2652
rect 5070 2648 5074 2652
rect 5086 2648 5090 2652
rect 5166 2648 5170 2652
rect 158 2638 162 2642
rect 758 2638 762 2642
rect 902 2638 906 2642
rect 1182 2638 1186 2642
rect 1198 2638 1202 2642
rect 1470 2638 1474 2642
rect 1662 2638 1666 2642
rect 2206 2638 2210 2642
rect 2246 2638 2250 2642
rect 2534 2638 2538 2642
rect 3694 2638 3698 2642
rect 4158 2638 4162 2642
rect 3134 2628 3138 2632
rect 4806 2628 4810 2632
rect 342 2618 346 2622
rect 478 2618 482 2622
rect 726 2618 730 2622
rect 870 2618 874 2622
rect 1446 2618 1450 2622
rect 1742 2618 1746 2622
rect 1790 2618 1794 2622
rect 1982 2618 1986 2622
rect 2622 2618 2626 2622
rect 2646 2618 2650 2622
rect 2870 2618 2874 2622
rect 3078 2618 3082 2622
rect 3278 2618 3282 2622
rect 3358 2618 3362 2622
rect 3526 2618 3530 2622
rect 3566 2618 3570 2622
rect 3726 2618 3730 2622
rect 4070 2618 4074 2622
rect 4110 2618 4114 2622
rect 4198 2618 4202 2622
rect 4254 2618 4258 2622
rect 4382 2618 4386 2622
rect 4422 2618 4426 2622
rect 4550 2618 4554 2622
rect 4822 2618 4826 2622
rect 5118 2618 5122 2622
rect 5150 2618 5154 2622
rect 538 2603 542 2607
rect 545 2603 549 2607
rect 1562 2603 1566 2607
rect 1569 2603 1573 2607
rect 2586 2603 2590 2607
rect 2593 2603 2597 2607
rect 3610 2603 3614 2607
rect 3617 2603 3621 2607
rect 4634 2603 4638 2607
rect 4641 2603 4645 2607
rect 246 2588 250 2592
rect 606 2588 610 2592
rect 750 2588 754 2592
rect 774 2588 778 2592
rect 1430 2588 1434 2592
rect 1518 2588 1522 2592
rect 1702 2588 1706 2592
rect 2350 2588 2354 2592
rect 2406 2588 2410 2592
rect 3742 2588 3746 2592
rect 3974 2588 3978 2592
rect 4078 2588 4082 2592
rect 4766 2588 4770 2592
rect 4862 2588 4866 2592
rect 1806 2578 1810 2582
rect 4462 2578 4466 2582
rect 526 2568 530 2572
rect 1342 2568 1346 2572
rect 2158 2568 2162 2572
rect 2414 2568 2418 2572
rect 2558 2568 2562 2572
rect 2654 2568 2658 2572
rect 2774 2568 2778 2572
rect 3086 2568 3090 2572
rect 3854 2568 3858 2572
rect 4646 2568 4650 2572
rect 4918 2568 4922 2572
rect 5110 2568 5114 2572
rect 470 2558 474 2562
rect 486 2558 490 2562
rect 502 2558 506 2562
rect 622 2558 626 2562
rect 758 2558 762 2562
rect 38 2548 42 2552
rect 62 2548 66 2552
rect 126 2548 130 2552
rect 134 2548 138 2552
rect 190 2548 194 2552
rect 278 2548 282 2552
rect 318 2548 322 2552
rect 382 2548 386 2552
rect 398 2548 402 2552
rect 430 2548 434 2552
rect 438 2548 442 2552
rect 494 2548 498 2552
rect 534 2548 538 2552
rect 574 2548 578 2552
rect 582 2548 586 2552
rect 590 2548 594 2552
rect 710 2547 714 2551
rect 774 2548 778 2552
rect 798 2558 802 2562
rect 830 2558 834 2562
rect 1038 2558 1042 2562
rect 1054 2558 1058 2562
rect 1134 2558 1138 2562
rect 1150 2558 1154 2562
rect 1366 2558 1370 2562
rect 798 2548 802 2552
rect 814 2548 818 2552
rect 846 2548 850 2552
rect 862 2548 866 2552
rect 910 2548 914 2552
rect 966 2548 970 2552
rect 998 2547 1002 2551
rect 1038 2548 1042 2552
rect 1070 2548 1074 2552
rect 1110 2548 1114 2552
rect 1158 2548 1162 2552
rect 1190 2548 1194 2552
rect 1198 2548 1202 2552
rect 1206 2548 1210 2552
rect 1230 2548 1234 2552
rect 1278 2548 1282 2552
rect 1302 2548 1306 2552
rect 1366 2548 1370 2552
rect 1390 2558 1394 2562
rect 1462 2558 1466 2562
rect 1414 2548 1418 2552
rect 1486 2558 1490 2562
rect 1678 2558 1682 2562
rect 1486 2548 1490 2552
rect 1502 2548 1506 2552
rect 1510 2548 1514 2552
rect 1534 2548 1538 2552
rect 1598 2548 1602 2552
rect 1894 2558 1898 2562
rect 2070 2558 2074 2562
rect 2150 2558 2154 2562
rect 2270 2558 2274 2562
rect 2310 2558 2314 2562
rect 2430 2558 2434 2562
rect 2446 2558 2450 2562
rect 2462 2558 2466 2562
rect 2638 2558 2642 2562
rect 2742 2558 2746 2562
rect 2758 2558 2762 2562
rect 2790 2558 2794 2562
rect 1702 2548 1706 2552
rect 1742 2548 1746 2552
rect 1782 2548 1786 2552
rect 1790 2548 1794 2552
rect 1814 2548 1818 2552
rect 1822 2548 1826 2552
rect 1830 2548 1834 2552
rect 1838 2548 1842 2552
rect 1862 2548 1866 2552
rect 1902 2548 1906 2552
rect 1934 2548 1938 2552
rect 1942 2548 1946 2552
rect 1974 2548 1978 2552
rect 1982 2548 1986 2552
rect 2014 2548 2018 2552
rect 2022 2548 2026 2552
rect 2094 2548 2098 2552
rect 2126 2548 2130 2552
rect 2134 2548 2138 2552
rect 2214 2548 2218 2552
rect 2270 2548 2274 2552
rect 2334 2548 2338 2552
rect 2366 2548 2370 2552
rect 2382 2548 2386 2552
rect 2398 2548 2402 2552
rect 2422 2548 2426 2552
rect 2446 2548 2450 2552
rect 2510 2548 2514 2552
rect 2566 2548 2570 2552
rect 2630 2548 2634 2552
rect 2662 2548 2666 2552
rect 2694 2548 2698 2552
rect 2702 2548 2706 2552
rect 2742 2548 2746 2552
rect 2782 2548 2786 2552
rect 2798 2548 2802 2552
rect 2814 2548 2818 2552
rect 2830 2548 2834 2552
rect 2846 2548 2850 2552
rect 2910 2548 2914 2552
rect 2958 2548 2962 2552
rect 2982 2558 2986 2562
rect 3006 2548 3010 2552
rect 3134 2547 3138 2551
rect 3174 2548 3178 2552
rect 3182 2548 3186 2552
rect 3198 2558 3202 2562
rect 3486 2558 3490 2562
rect 3294 2548 3298 2552
rect 3326 2548 3330 2552
rect 3342 2548 3346 2552
rect 3510 2558 3514 2562
rect 3718 2558 3722 2562
rect 3726 2558 3730 2562
rect 3774 2558 3778 2562
rect 3374 2547 3378 2551
rect 3510 2548 3514 2552
rect 3550 2547 3554 2551
rect 3654 2548 3658 2552
rect 3686 2548 3690 2552
rect 3702 2548 3706 2552
rect 3710 2548 3714 2552
rect 3750 2548 3754 2552
rect 3774 2548 3778 2552
rect 3790 2548 3794 2552
rect 3814 2558 3818 2562
rect 4454 2558 4458 2562
rect 4574 2558 4578 2562
rect 4878 2558 4882 2562
rect 5126 2558 5130 2562
rect 5150 2558 5154 2562
rect 3910 2548 3914 2552
rect 4014 2548 4018 2552
rect 102 2538 106 2542
rect 134 2538 138 2542
rect 166 2538 170 2542
rect 270 2538 274 2542
rect 294 2538 298 2542
rect 326 2538 330 2542
rect 390 2538 394 2542
rect 446 2538 450 2542
rect 494 2538 498 2542
rect 518 2538 522 2542
rect 638 2538 642 2542
rect 726 2538 730 2542
rect 742 2538 746 2542
rect 766 2538 770 2542
rect 822 2538 826 2542
rect 854 2538 858 2542
rect 878 2538 882 2542
rect 902 2538 906 2542
rect 982 2538 986 2542
rect 1030 2538 1034 2542
rect 1062 2538 1066 2542
rect 1078 2538 1082 2542
rect 1102 2538 1106 2542
rect 1150 2538 1154 2542
rect 1166 2538 1170 2542
rect 1182 2538 1186 2542
rect 1406 2538 1410 2542
rect 1430 2538 1434 2542
rect 1446 2538 1450 2542
rect 1494 2538 1498 2542
rect 1574 2538 1578 2542
rect 1662 2538 1666 2542
rect 1710 2538 1714 2542
rect 1870 2538 1874 2542
rect 1878 2538 1882 2542
rect 1910 2538 1914 2542
rect 1926 2538 1930 2542
rect 1950 2538 1954 2542
rect 1966 2538 1970 2542
rect 1990 2538 1994 2542
rect 1998 2538 2002 2542
rect 2014 2538 2018 2542
rect 2046 2538 2050 2542
rect 2054 2538 2058 2542
rect 2094 2538 2098 2542
rect 2102 2538 2106 2542
rect 2118 2538 2122 2542
rect 2134 2538 2138 2542
rect 2254 2538 2258 2542
rect 2374 2538 2378 2542
rect 2390 2538 2394 2542
rect 2438 2538 2442 2542
rect 2574 2538 2578 2542
rect 2654 2538 2658 2542
rect 2662 2538 2666 2542
rect 2686 2538 2690 2542
rect 2694 2538 2698 2542
rect 2726 2538 2730 2542
rect 2758 2538 2762 2542
rect 2806 2538 2810 2542
rect 2822 2538 2826 2542
rect 2934 2538 2938 2542
rect 2950 2538 2954 2542
rect 2966 2538 2970 2542
rect 2998 2538 3002 2542
rect 3150 2538 3154 2542
rect 3166 2538 3170 2542
rect 3214 2538 3218 2542
rect 3222 2538 3226 2542
rect 3286 2538 3290 2542
rect 3334 2538 3338 2542
rect 3462 2538 3466 2542
rect 3470 2538 3474 2542
rect 3518 2538 3522 2542
rect 3654 2538 3658 2542
rect 3662 2538 3666 2542
rect 3678 2538 3682 2542
rect 3694 2538 3698 2542
rect 3750 2538 3754 2542
rect 3758 2538 3762 2542
rect 4038 2547 4042 2551
rect 4094 2548 4098 2552
rect 4126 2548 4130 2552
rect 4150 2548 4154 2552
rect 4158 2548 4162 2552
rect 4166 2548 4170 2552
rect 4198 2548 4202 2552
rect 4246 2547 4250 2551
rect 4342 2548 4346 2552
rect 4406 2548 4410 2552
rect 4430 2548 4434 2552
rect 3814 2538 3818 2542
rect 3830 2538 3834 2542
rect 3846 2538 3850 2542
rect 3918 2538 3922 2542
rect 3950 2538 3954 2542
rect 4110 2538 4114 2542
rect 4174 2538 4178 2542
rect 4190 2538 4194 2542
rect 4214 2538 4218 2542
rect 4254 2538 4258 2542
rect 4334 2538 4338 2542
rect 4366 2538 4370 2542
rect 4526 2547 4530 2551
rect 4598 2548 4602 2552
rect 4614 2548 4618 2552
rect 4638 2548 4642 2552
rect 4710 2548 4714 2552
rect 4750 2548 4754 2552
rect 4782 2548 4786 2552
rect 4814 2548 4818 2552
rect 4862 2548 4866 2552
rect 4910 2548 4914 2552
rect 4982 2547 4986 2551
rect 5046 2548 5050 2552
rect 5158 2548 5162 2552
rect 5190 2548 5194 2552
rect 4438 2538 4442 2542
rect 4542 2538 4546 2542
rect 4558 2538 4562 2542
rect 4622 2538 4626 2542
rect 4734 2538 4738 2542
rect 4790 2538 4794 2542
rect 4806 2538 4810 2542
rect 4902 2538 4906 2542
rect 4974 2538 4978 2542
rect 5054 2538 5058 2542
rect 5110 2538 5114 2542
rect 5134 2538 5138 2542
rect 102 2528 106 2532
rect 142 2528 146 2532
rect 150 2528 154 2532
rect 254 2528 258 2532
rect 414 2528 418 2532
rect 462 2528 466 2532
rect 862 2528 866 2532
rect 886 2528 890 2532
rect 918 2528 922 2532
rect 1126 2528 1130 2532
rect 1214 2528 1218 2532
rect 2110 2528 2114 2532
rect 2222 2528 2226 2532
rect 2278 2528 2282 2532
rect 2294 2528 2298 2532
rect 2494 2528 2498 2532
rect 2598 2528 2602 2532
rect 2838 2528 2842 2532
rect 3022 2528 3026 2532
rect 3310 2528 3314 2532
rect 3374 2528 3378 2532
rect 3550 2528 3554 2532
rect 3838 2528 3842 2532
rect 4078 2528 4082 2532
rect 4582 2528 4586 2532
rect 4830 2528 4834 2532
rect 4838 2528 4842 2532
rect 4886 2528 4890 2532
rect 5174 2528 5178 2532
rect 94 2518 98 2522
rect 262 2518 266 2522
rect 374 2518 378 2522
rect 454 2518 458 2522
rect 566 2518 570 2522
rect 630 2518 634 2522
rect 646 2518 650 2522
rect 798 2518 802 2522
rect 830 2518 834 2522
rect 894 2518 898 2522
rect 1174 2518 1178 2522
rect 1654 2518 1658 2522
rect 1726 2518 1730 2522
rect 1758 2518 1762 2522
rect 1886 2518 1890 2522
rect 1926 2518 1930 2522
rect 1958 2518 1962 2522
rect 2286 2518 2290 2522
rect 2582 2518 2586 2522
rect 2678 2518 2682 2522
rect 2710 2518 2714 2522
rect 2782 2518 2786 2522
rect 2854 2518 2858 2522
rect 3038 2518 3042 2522
rect 3438 2518 3442 2522
rect 3454 2518 3458 2522
rect 3662 2518 3666 2522
rect 3766 2518 3770 2522
rect 3958 2518 3962 2522
rect 4310 2518 4314 2522
rect 4318 2518 4322 2522
rect 4382 2518 4386 2522
rect 4414 2518 4418 2522
rect 4454 2518 4458 2522
rect 4566 2518 4570 2522
rect 4766 2518 4770 2522
rect 4846 2518 4850 2522
rect 4894 2518 4898 2522
rect 5118 2518 5122 2522
rect 5142 2518 5146 2522
rect 1050 2503 1054 2507
rect 1057 2503 1061 2507
rect 2074 2503 2078 2507
rect 2081 2503 2085 2507
rect 3098 2503 3102 2507
rect 3105 2503 3109 2507
rect 4114 2503 4118 2507
rect 4121 2503 4125 2507
rect 150 2488 154 2492
rect 254 2488 258 2492
rect 374 2488 378 2492
rect 494 2488 498 2492
rect 918 2488 922 2492
rect 1046 2488 1050 2492
rect 1158 2488 1162 2492
rect 1182 2488 1186 2492
rect 1342 2488 1346 2492
rect 1382 2488 1386 2492
rect 1486 2488 1490 2492
rect 1510 2488 1514 2492
rect 1574 2488 1578 2492
rect 1686 2488 1690 2492
rect 1702 2488 1706 2492
rect 1742 2488 1746 2492
rect 1774 2488 1778 2492
rect 1806 2488 1810 2492
rect 1862 2488 1866 2492
rect 2006 2488 2010 2492
rect 2030 2488 2034 2492
rect 2142 2488 2146 2492
rect 2214 2488 2218 2492
rect 2238 2488 2242 2492
rect 2278 2488 2282 2492
rect 2310 2488 2314 2492
rect 2550 2488 2554 2492
rect 3046 2488 3050 2492
rect 3086 2488 3090 2492
rect 3182 2488 3186 2492
rect 3270 2488 3274 2492
rect 3382 2488 3386 2492
rect 3470 2488 3474 2492
rect 3542 2488 3546 2492
rect 3742 2488 3746 2492
rect 3806 2488 3810 2492
rect 4078 2488 4082 2492
rect 4310 2488 4314 2492
rect 4622 2488 4626 2492
rect 4742 2488 4746 2492
rect 4814 2488 4818 2492
rect 4878 2488 4882 2492
rect 4894 2488 4898 2492
rect 4910 2488 4914 2492
rect 5006 2488 5010 2492
rect 5134 2488 5138 2492
rect 5174 2488 5178 2492
rect 366 2478 370 2482
rect 510 2478 514 2482
rect 702 2478 706 2482
rect 854 2478 858 2482
rect 6 2468 10 2472
rect 30 2468 34 2472
rect 134 2468 138 2472
rect 230 2468 234 2472
rect 398 2468 402 2472
rect 590 2468 594 2472
rect 638 2468 642 2472
rect 646 2468 650 2472
rect 774 2468 778 2472
rect 886 2468 890 2472
rect 902 2468 906 2472
rect 934 2478 938 2482
rect 982 2478 986 2482
rect 1094 2478 1098 2482
rect 1422 2478 1426 2482
rect 1246 2468 1250 2472
rect 22 2458 26 2462
rect 86 2458 90 2462
rect 118 2459 122 2463
rect 182 2458 186 2462
rect 214 2459 218 2463
rect 246 2458 250 2462
rect 302 2458 306 2462
rect 310 2458 314 2462
rect 382 2458 386 2462
rect 422 2458 426 2462
rect 502 2458 506 2462
rect 526 2458 530 2462
rect 542 2458 546 2462
rect 550 2458 554 2462
rect 574 2458 578 2462
rect 598 2458 602 2462
rect 654 2458 658 2462
rect 670 2458 674 2462
rect 702 2459 706 2463
rect 782 2458 786 2462
rect 806 2458 810 2462
rect 814 2458 818 2462
rect 838 2458 842 2462
rect 870 2458 874 2462
rect 902 2458 906 2462
rect 950 2458 954 2462
rect 982 2459 986 2463
rect 1502 2468 1506 2472
rect 1526 2478 1530 2482
rect 1598 2478 1602 2482
rect 1670 2478 1674 2482
rect 1678 2478 1682 2482
rect 1710 2478 1714 2482
rect 1734 2478 1738 2482
rect 2054 2478 2058 2482
rect 2286 2478 2290 2482
rect 2390 2478 2394 2482
rect 2574 2478 2578 2482
rect 2790 2478 2794 2482
rect 3510 2478 3514 2482
rect 3798 2478 3802 2482
rect 3974 2478 3978 2482
rect 4158 2478 4162 2482
rect 4358 2478 4362 2482
rect 4646 2478 4650 2482
rect 4782 2478 4786 2482
rect 4974 2478 4978 2482
rect 5102 2478 5106 2482
rect 5182 2478 5186 2482
rect 1654 2468 1658 2472
rect 1670 2468 1674 2472
rect 1758 2468 1762 2472
rect 1798 2468 1802 2472
rect 1830 2468 1834 2472
rect 1854 2468 1858 2472
rect 1878 2468 1882 2472
rect 1894 2468 1898 2472
rect 1910 2468 1914 2472
rect 1934 2468 1938 2472
rect 1942 2468 1946 2472
rect 1990 2468 1994 2472
rect 2006 2468 2010 2472
rect 2038 2468 2042 2472
rect 2046 2468 2050 2472
rect 2070 2468 2074 2472
rect 2118 2468 2122 2472
rect 2126 2468 2130 2472
rect 2158 2468 2162 2472
rect 2166 2468 2170 2472
rect 2182 2468 2186 2472
rect 2198 2468 2202 2472
rect 2230 2468 2234 2472
rect 2246 2468 2250 2472
rect 2270 2468 2274 2472
rect 2302 2468 2306 2472
rect 2318 2468 2322 2472
rect 2342 2468 2346 2472
rect 2358 2468 2362 2472
rect 2430 2468 2434 2472
rect 2446 2468 2450 2472
rect 2502 2468 2506 2472
rect 2526 2468 2530 2472
rect 2566 2468 2570 2472
rect 2574 2468 2578 2472
rect 2590 2468 2594 2472
rect 2646 2468 2650 2472
rect 2710 2468 2714 2472
rect 2726 2468 2730 2472
rect 2742 2468 2746 2472
rect 2894 2468 2898 2472
rect 2902 2468 2906 2472
rect 2950 2468 2954 2472
rect 2958 2468 2962 2472
rect 3014 2468 3018 2472
rect 3038 2468 3042 2472
rect 3054 2468 3058 2472
rect 3078 2468 3082 2472
rect 3094 2468 3098 2472
rect 3134 2468 3138 2472
rect 3142 2468 3146 2472
rect 3158 2468 3162 2472
rect 3166 2468 3170 2472
rect 3198 2468 3202 2472
rect 3214 2468 3218 2472
rect 3238 2468 3242 2472
rect 3254 2468 3258 2472
rect 3286 2468 3290 2472
rect 3294 2468 3298 2472
rect 3334 2468 3338 2472
rect 3358 2468 3362 2472
rect 3366 2468 3370 2472
rect 3390 2468 3394 2472
rect 3414 2468 3418 2472
rect 3430 2468 3434 2472
rect 3446 2468 3450 2472
rect 3462 2468 3466 2472
rect 3566 2468 3570 2472
rect 3590 2468 3594 2472
rect 3678 2468 3682 2472
rect 3758 2468 3762 2472
rect 3782 2468 3786 2472
rect 3862 2468 3866 2472
rect 3894 2468 3898 2472
rect 3902 2468 3906 2472
rect 3918 2468 3922 2472
rect 3958 2468 3962 2472
rect 3966 2468 3970 2472
rect 3982 2468 3986 2472
rect 4014 2468 4018 2472
rect 4038 2468 4042 2472
rect 4054 2468 4058 2472
rect 4086 2468 4090 2472
rect 4102 2468 4106 2472
rect 4110 2468 4114 2472
rect 4118 2468 4122 2472
rect 4142 2468 4146 2472
rect 4174 2468 4178 2472
rect 4254 2468 4258 2472
rect 4414 2468 4418 2472
rect 4478 2468 4482 2472
rect 4534 2468 4538 2472
rect 4550 2468 4554 2472
rect 4582 2468 4586 2472
rect 4686 2468 4690 2472
rect 4750 2468 4754 2472
rect 4822 2468 4826 2472
rect 4854 2468 4858 2472
rect 4862 2468 4866 2472
rect 4886 2468 4890 2472
rect 5054 2468 5058 2472
rect 5142 2468 5146 2472
rect 5166 2468 5170 2472
rect 1102 2458 1106 2462
rect 1166 2458 1170 2462
rect 1206 2458 1210 2462
rect 1230 2458 1234 2462
rect 1238 2458 1242 2462
rect 1278 2458 1282 2462
rect 1294 2458 1298 2462
rect 1302 2458 1306 2462
rect 1358 2458 1362 2462
rect 1430 2458 1434 2462
rect 1494 2458 1498 2462
rect 1542 2458 1546 2462
rect 1590 2458 1594 2462
rect 1614 2458 1618 2462
rect 1694 2458 1698 2462
rect 1718 2458 1722 2462
rect 1790 2458 1794 2462
rect 1822 2458 1826 2462
rect 1854 2458 1858 2462
rect 1902 2458 1906 2462
rect 1974 2458 1978 2462
rect 2014 2458 2018 2462
rect 2110 2458 2114 2462
rect 2150 2458 2154 2462
rect 2158 2458 2162 2462
rect 2174 2458 2178 2462
rect 2190 2458 2194 2462
rect 2222 2458 2226 2462
rect 2254 2458 2258 2462
rect 2262 2458 2266 2462
rect 2294 2458 2298 2462
rect 2326 2458 2330 2462
rect 2334 2458 2338 2462
rect 2366 2458 2370 2462
rect 2374 2458 2378 2462
rect 2406 2458 2410 2462
rect 2438 2458 2442 2462
rect 2470 2458 2474 2462
rect 2502 2458 2506 2462
rect 2534 2458 2538 2462
rect 2558 2458 2562 2462
rect 2598 2458 2602 2462
rect 2638 2458 2642 2462
rect 2646 2458 2650 2462
rect 2686 2458 2690 2462
rect 2694 2458 2698 2462
rect 2702 2458 2706 2462
rect 2734 2458 2738 2462
rect 2766 2458 2770 2462
rect 2774 2458 2778 2462
rect 2782 2458 2786 2462
rect 2814 2458 2818 2462
rect 2822 2458 2826 2462
rect 2830 2458 2834 2462
rect 2886 2458 2890 2462
rect 2926 2458 2930 2462
rect 2966 2458 2970 2462
rect 2990 2458 2994 2462
rect 3022 2458 3026 2462
rect 3030 2458 3034 2462
rect 3062 2458 3066 2462
rect 3070 2458 3074 2462
rect 3102 2458 3106 2462
rect 3118 2458 3122 2462
rect 3166 2458 3170 2462
rect 3190 2458 3194 2462
rect 3206 2458 3210 2462
rect 3222 2458 3226 2462
rect 3262 2458 3266 2462
rect 3302 2458 3306 2462
rect 3326 2458 3330 2462
rect 3358 2458 3362 2462
rect 3366 2458 3370 2462
rect 3398 2458 3402 2462
rect 3406 2458 3410 2462
rect 3422 2458 3426 2462
rect 3446 2458 3450 2462
rect 3494 2458 3498 2462
rect 3526 2458 3530 2462
rect 3598 2458 3602 2462
rect 3622 2458 3626 2462
rect 3670 2459 3674 2463
rect 3766 2458 3770 2462
rect 3814 2458 3818 2462
rect 3822 2458 3826 2462
rect 3846 2458 3850 2462
rect 3886 2458 3890 2462
rect 3910 2458 3914 2462
rect 3934 2458 3938 2462
rect 3958 2458 3962 2462
rect 3990 2458 3994 2462
rect 3998 2458 4002 2462
rect 4030 2458 4034 2462
rect 4070 2458 4074 2462
rect 4086 2458 4090 2462
rect 4126 2458 4130 2462
rect 4150 2458 4154 2462
rect 4190 2458 4194 2462
rect 4214 2458 4218 2462
rect 4262 2458 4266 2462
rect 4334 2458 4338 2462
rect 4374 2458 4378 2462
rect 4422 2458 4426 2462
rect 4446 2458 4450 2462
rect 4462 2458 4466 2462
rect 4470 2458 4474 2462
rect 4486 2458 4490 2462
rect 4494 2458 4498 2462
rect 4526 2458 4530 2462
rect 4574 2458 4578 2462
rect 4606 2458 4610 2462
rect 4678 2459 4682 2463
rect 4758 2458 4762 2462
rect 4798 2458 4802 2462
rect 4830 2458 4834 2462
rect 4902 2458 4906 2462
rect 4942 2458 4946 2462
rect 4966 2458 4970 2462
rect 5062 2458 5066 2462
rect 5118 2458 5122 2462
rect 5150 2458 5154 2462
rect 5158 2458 5162 2462
rect 286 2448 290 2452
rect 598 2448 602 2452
rect 622 2448 626 2452
rect 670 2448 674 2452
rect 798 2448 802 2452
rect 830 2448 834 2452
rect 894 2448 898 2452
rect 1142 2448 1146 2452
rect 1278 2448 1282 2452
rect 1622 2448 1626 2452
rect 1742 2448 1746 2452
rect 1814 2448 1818 2452
rect 1846 2448 1850 2452
rect 1862 2448 1866 2452
rect 1886 2448 1890 2452
rect 1918 2448 1922 2452
rect 2022 2448 2026 2452
rect 2078 2448 2082 2452
rect 2430 2448 2434 2452
rect 2462 2448 2466 2452
rect 2478 2448 2482 2452
rect 2510 2448 2514 2452
rect 2622 2448 2626 2452
rect 2638 2448 2642 2452
rect 2870 2448 2874 2452
rect 2918 2448 2922 2452
rect 2934 2448 2938 2452
rect 2982 2448 2986 2452
rect 3182 2448 3186 2452
rect 3270 2448 3274 2452
rect 3302 2448 3306 2452
rect 3318 2448 3322 2452
rect 3446 2448 3450 2452
rect 3462 2448 3466 2452
rect 3550 2448 3554 2452
rect 3574 2448 3578 2452
rect 3742 2448 3746 2452
rect 3934 2448 3938 2452
rect 4038 2448 4042 2452
rect 4070 2448 4074 2452
rect 4318 2448 4322 2452
rect 4334 2448 4338 2452
rect 4374 2448 4378 2452
rect 4398 2448 4402 2452
rect 4454 2448 4458 2452
rect 4550 2448 4554 2452
rect 4558 2448 4562 2452
rect 4590 2448 4594 2452
rect 4606 2448 4610 2452
rect 4774 2448 4778 2452
rect 4838 2448 4842 2452
rect 4854 2448 4858 2452
rect 4878 2448 4882 2452
rect 1934 2438 1938 2442
rect 2214 2438 2218 2442
rect 2358 2438 2362 2442
rect 3238 2438 3242 2442
rect 3630 2438 3634 2442
rect 3734 2438 3738 2442
rect 3942 2438 3946 2442
rect 1950 2428 1954 2432
rect 4502 2428 4506 2432
rect 4542 2428 4546 2432
rect 478 2418 482 2422
rect 566 2418 570 2422
rect 766 2418 770 2422
rect 782 2418 786 2422
rect 1214 2418 1218 2422
rect 1286 2418 1290 2422
rect 1318 2418 1322 2422
rect 1382 2418 1386 2422
rect 1654 2418 1658 2422
rect 1718 2418 1722 2422
rect 2518 2418 2522 2422
rect 2670 2418 2674 2422
rect 2710 2418 2714 2422
rect 2838 2418 2842 2422
rect 2998 2418 3002 2422
rect 3334 2418 3338 2422
rect 3582 2418 3586 2422
rect 3638 2418 3642 2422
rect 3878 2418 3882 2422
rect 4198 2418 4202 2422
rect 4758 2418 4762 2422
rect 538 2403 542 2407
rect 545 2403 549 2407
rect 1562 2403 1566 2407
rect 1569 2403 1573 2407
rect 2586 2403 2590 2407
rect 2593 2403 2597 2407
rect 3610 2403 3614 2407
rect 3617 2403 3621 2407
rect 4634 2403 4638 2407
rect 4641 2403 4645 2407
rect 758 2388 762 2392
rect 862 2388 866 2392
rect 950 2388 954 2392
rect 1190 2388 1194 2392
rect 1294 2388 1298 2392
rect 1422 2388 1426 2392
rect 1710 2388 1714 2392
rect 1966 2388 1970 2392
rect 2678 2388 2682 2392
rect 2710 2388 2714 2392
rect 2750 2388 2754 2392
rect 2782 2388 2786 2392
rect 3118 2388 3122 2392
rect 3150 2388 3154 2392
rect 3190 2388 3194 2392
rect 3278 2388 3282 2392
rect 3430 2388 3434 2392
rect 4094 2388 4098 2392
rect 4182 2388 4186 2392
rect 4366 2388 4370 2392
rect 4854 2388 4858 2392
rect 3014 2378 3018 2382
rect 4766 2378 4770 2382
rect 6 2368 10 2372
rect 182 2368 186 2372
rect 278 2368 282 2372
rect 374 2368 378 2372
rect 486 2368 490 2372
rect 534 2368 538 2372
rect 838 2368 842 2372
rect 1446 2368 1450 2372
rect 1638 2368 1642 2372
rect 1854 2368 1858 2372
rect 1918 2368 1922 2372
rect 2382 2368 2386 2372
rect 2534 2368 2538 2372
rect 4222 2368 4226 2372
rect 4342 2368 4346 2372
rect 4926 2368 4930 2372
rect 5134 2368 5138 2372
rect 5150 2368 5154 2372
rect 150 2358 154 2362
rect 166 2358 170 2362
rect 358 2358 362 2362
rect 390 2358 394 2362
rect 502 2358 506 2362
rect 62 2348 66 2352
rect 94 2347 98 2351
rect 134 2348 138 2352
rect 150 2348 154 2352
rect 166 2348 170 2352
rect 214 2347 218 2351
rect 286 2348 290 2352
rect 318 2348 322 2352
rect 326 2348 330 2352
rect 342 2348 346 2352
rect 374 2348 378 2352
rect 430 2348 434 2352
rect 502 2348 506 2352
rect 814 2358 818 2362
rect 822 2358 826 2362
rect 854 2358 858 2362
rect 1142 2358 1146 2362
rect 1214 2358 1218 2362
rect 1318 2358 1322 2362
rect 558 2348 562 2352
rect 574 2348 578 2352
rect 606 2348 610 2352
rect 614 2348 618 2352
rect 630 2348 634 2352
rect 638 2348 642 2352
rect 646 2348 650 2352
rect 694 2348 698 2352
rect 766 2348 770 2352
rect 790 2348 794 2352
rect 798 2348 802 2352
rect 838 2348 842 2352
rect 878 2348 882 2352
rect 886 2348 890 2352
rect 910 2348 914 2352
rect 918 2348 922 2352
rect 926 2348 930 2352
rect 934 2348 938 2352
rect 958 2348 962 2352
rect 1006 2348 1010 2352
rect 1102 2348 1106 2352
rect 86 2338 90 2342
rect 126 2338 130 2342
rect 158 2338 162 2342
rect 230 2338 234 2342
rect 334 2338 338 2342
rect 366 2338 370 2342
rect 406 2338 410 2342
rect 494 2338 498 2342
rect 566 2338 570 2342
rect 622 2338 626 2342
rect 662 2338 666 2342
rect 790 2338 794 2342
rect 846 2338 850 2342
rect 870 2338 874 2342
rect 1134 2348 1138 2352
rect 1174 2348 1178 2352
rect 1198 2348 1202 2352
rect 1206 2348 1210 2352
rect 1270 2348 1274 2352
rect 1278 2348 1282 2352
rect 1302 2348 1306 2352
rect 1310 2348 1314 2352
rect 1318 2348 1322 2352
rect 1334 2348 1338 2352
rect 1350 2348 1354 2352
rect 1358 2348 1362 2352
rect 1382 2348 1386 2352
rect 1390 2348 1394 2352
rect 1398 2348 1402 2352
rect 1406 2348 1410 2352
rect 1430 2348 1434 2352
rect 1494 2348 1498 2352
rect 1518 2348 1522 2352
rect 1582 2348 1586 2352
rect 1606 2358 1610 2362
rect 1670 2358 1674 2362
rect 2174 2358 2178 2362
rect 2190 2358 2194 2362
rect 1630 2348 1634 2352
rect 1662 2348 1666 2352
rect 1710 2348 1714 2352
rect 1718 2348 1722 2352
rect 1750 2348 1754 2352
rect 1798 2348 1802 2352
rect 1006 2338 1010 2342
rect 1110 2338 1114 2342
rect 1126 2338 1130 2342
rect 1134 2338 1138 2342
rect 1158 2338 1162 2342
rect 1230 2338 1234 2342
rect 1238 2338 1242 2342
rect 1342 2338 1346 2342
rect 1822 2347 1826 2351
rect 1878 2348 1882 2352
rect 1894 2348 1898 2352
rect 1958 2348 1962 2352
rect 1990 2348 1994 2352
rect 2022 2348 2026 2352
rect 2030 2348 2034 2352
rect 2070 2348 2074 2352
rect 2110 2348 2114 2352
rect 2142 2348 2146 2352
rect 2150 2348 2154 2352
rect 2182 2348 2186 2352
rect 2206 2348 2210 2352
rect 2254 2348 2258 2352
rect 2278 2348 2282 2352
rect 2286 2348 2290 2352
rect 2318 2348 2322 2352
rect 2334 2348 2338 2352
rect 2358 2358 2362 2362
rect 2486 2358 2490 2362
rect 2550 2358 2554 2362
rect 2822 2358 2826 2362
rect 2950 2358 2954 2362
rect 2422 2348 2426 2352
rect 2502 2348 2506 2352
rect 2510 2348 2514 2352
rect 2542 2348 2546 2352
rect 2582 2348 2586 2352
rect 2622 2348 2626 2352
rect 2662 2348 2666 2352
rect 2686 2348 2690 2352
rect 2694 2348 2698 2352
rect 2726 2348 2730 2352
rect 2766 2348 2770 2352
rect 2774 2348 2778 2352
rect 2798 2348 2802 2352
rect 2838 2348 2842 2352
rect 2878 2348 2882 2352
rect 2950 2348 2954 2352
rect 2974 2358 2978 2362
rect 3206 2358 3210 2362
rect 2998 2348 3002 2352
rect 3030 2348 3034 2352
rect 3086 2348 3090 2352
rect 3142 2348 3146 2352
rect 3166 2348 3170 2352
rect 3174 2348 3178 2352
rect 3230 2348 3234 2352
rect 3262 2348 3266 2352
rect 3270 2348 3274 2352
rect 3310 2348 3314 2352
rect 3342 2348 3346 2352
rect 3350 2348 3354 2352
rect 3382 2348 3386 2352
rect 3398 2348 3402 2352
rect 3742 2358 3746 2362
rect 3782 2358 3786 2362
rect 3846 2358 3850 2362
rect 3462 2348 3466 2352
rect 3486 2348 3490 2352
rect 3526 2348 3530 2352
rect 3534 2348 3538 2352
rect 3558 2348 3562 2352
rect 3574 2348 3578 2352
rect 3638 2348 3642 2352
rect 3702 2348 3706 2352
rect 3790 2348 3794 2352
rect 3830 2348 3834 2352
rect 3870 2358 3874 2362
rect 4022 2358 4026 2362
rect 4054 2358 4058 2362
rect 4166 2358 4170 2362
rect 4502 2358 4506 2362
rect 4534 2358 4538 2362
rect 4806 2358 4810 2362
rect 4822 2358 4826 2362
rect 4870 2358 4874 2362
rect 4878 2358 4882 2362
rect 4894 2358 4898 2362
rect 5110 2358 5114 2362
rect 3870 2348 3874 2352
rect 3910 2347 3914 2351
rect 3934 2348 3938 2352
rect 3982 2348 3986 2352
rect 3998 2348 4002 2352
rect 4014 2348 4018 2352
rect 4046 2348 4050 2352
rect 4086 2348 4090 2352
rect 4134 2348 4138 2352
rect 4182 2348 4186 2352
rect 4198 2348 4202 2352
rect 4246 2348 4250 2352
rect 4278 2347 4282 2351
rect 4350 2348 4354 2352
rect 4358 2348 4362 2352
rect 4382 2348 4386 2352
rect 4398 2348 4402 2352
rect 4446 2348 4450 2352
rect 4478 2348 4482 2352
rect 4518 2348 4522 2352
rect 4526 2348 4530 2352
rect 4598 2348 4602 2352
rect 4710 2348 4714 2352
rect 4750 2348 4754 2352
rect 4758 2348 4762 2352
rect 4782 2348 4786 2352
rect 4806 2348 4810 2352
rect 4854 2348 4858 2352
rect 4990 2347 4994 2351
rect 5054 2348 5058 2352
rect 5070 2348 5074 2352
rect 5102 2348 5106 2352
rect 5150 2348 5154 2352
rect 5174 2348 5178 2352
rect 1558 2338 1562 2342
rect 1590 2338 1594 2342
rect 1622 2338 1626 2342
rect 1638 2338 1642 2342
rect 1654 2338 1658 2342
rect 1686 2338 1690 2342
rect 1710 2338 1714 2342
rect 1742 2338 1746 2342
rect 1870 2338 1874 2342
rect 1942 2338 1946 2342
rect 1998 2338 2002 2342
rect 2022 2338 2026 2342
rect 2038 2338 2042 2342
rect 2054 2338 2058 2342
rect 2086 2338 2090 2342
rect 2150 2338 2154 2342
rect 2174 2338 2178 2342
rect 2206 2338 2210 2342
rect 2214 2338 2218 2342
rect 2230 2338 2234 2342
rect 2246 2338 2250 2342
rect 2294 2338 2298 2342
rect 2310 2338 2314 2342
rect 2326 2338 2330 2342
rect 2358 2338 2362 2342
rect 2374 2338 2378 2342
rect 2438 2338 2442 2342
rect 2518 2338 2522 2342
rect 2534 2338 2538 2342
rect 2566 2338 2570 2342
rect 2614 2338 2618 2342
rect 2854 2338 2858 2342
rect 2942 2338 2946 2342
rect 2990 2338 2994 2342
rect 3198 2338 3202 2342
rect 3222 2338 3226 2342
rect 3238 2338 3242 2342
rect 3246 2338 3250 2342
rect 3254 2338 3258 2342
rect 3278 2338 3282 2342
rect 3294 2338 3298 2342
rect 3302 2338 3306 2342
rect 3318 2338 3322 2342
rect 3334 2338 3338 2342
rect 3358 2338 3362 2342
rect 3422 2338 3426 2342
rect 3630 2338 3634 2342
rect 3758 2338 3762 2342
rect 3766 2338 3770 2342
rect 3814 2338 3818 2342
rect 3830 2338 3834 2342
rect 3878 2338 3882 2342
rect 3990 2338 3994 2342
rect 4006 2338 4010 2342
rect 4022 2338 4026 2342
rect 4038 2338 4042 2342
rect 4046 2338 4050 2342
rect 4070 2338 4074 2342
rect 4190 2338 4194 2342
rect 4238 2338 4242 2342
rect 4262 2338 4266 2342
rect 4454 2338 4458 2342
rect 4470 2338 4474 2342
rect 4486 2338 4490 2342
rect 4510 2338 4514 2342
rect 4590 2338 4594 2342
rect 4622 2338 4626 2342
rect 4734 2338 4738 2342
rect 4798 2338 4802 2342
rect 4846 2338 4850 2342
rect 4894 2338 4898 2342
rect 4902 2338 4906 2342
rect 4918 2338 4922 2342
rect 4982 2338 4986 2342
rect 5094 2338 5098 2342
rect 5126 2338 5130 2342
rect 5134 2338 5138 2342
rect 5158 2338 5162 2342
rect 782 2328 786 2332
rect 1694 2328 1698 2332
rect 1854 2328 1858 2332
rect 1886 2328 1890 2332
rect 1918 2328 1922 2332
rect 1926 2328 1930 2332
rect 1942 2328 1946 2332
rect 1982 2328 1986 2332
rect 2294 2328 2298 2332
rect 3070 2328 3074 2332
rect 3366 2328 3370 2332
rect 3398 2328 3402 2332
rect 3542 2328 3546 2332
rect 3598 2328 3602 2332
rect 3710 2328 3714 2332
rect 4214 2328 4218 2332
rect 4222 2328 4226 2332
rect 4430 2328 4434 2332
rect 4838 2328 4842 2332
rect 5022 2328 5026 2332
rect 5038 2328 5042 2332
rect 5054 2328 5058 2332
rect 5070 2328 5074 2332
rect 5078 2328 5082 2332
rect 5182 2328 5186 2332
rect 310 2318 314 2322
rect 358 2318 362 2322
rect 590 2318 594 2322
rect 742 2318 746 2322
rect 814 2318 818 2322
rect 1070 2318 1074 2322
rect 1214 2318 1218 2322
rect 1670 2318 1674 2322
rect 1742 2318 1746 2322
rect 1758 2318 1762 2322
rect 1950 2318 1954 2322
rect 2006 2318 2010 2322
rect 2046 2318 2050 2322
rect 2126 2318 2130 2322
rect 2198 2318 2202 2322
rect 2550 2318 2554 2322
rect 2638 2318 2642 2322
rect 2750 2318 2754 2322
rect 2934 2318 2938 2322
rect 3046 2318 3050 2322
rect 3118 2318 3122 2322
rect 3206 2318 3210 2322
rect 3326 2318 3330 2322
rect 3406 2318 3410 2322
rect 3622 2318 3626 2322
rect 3646 2318 3650 2322
rect 3742 2318 3746 2322
rect 3798 2318 3802 2322
rect 3974 2318 3978 2322
rect 4150 2318 4154 2322
rect 4206 2318 4210 2322
rect 4414 2318 4418 2322
rect 4502 2318 4506 2322
rect 4542 2318 4546 2322
rect 4654 2318 4658 2322
rect 4830 2318 4834 2322
rect 5030 2318 5034 2322
rect 5062 2318 5066 2322
rect 5110 2318 5114 2322
rect 1050 2303 1054 2307
rect 1057 2303 1061 2307
rect 2074 2303 2078 2307
rect 2081 2303 2085 2307
rect 3098 2303 3102 2307
rect 3105 2303 3109 2307
rect 4114 2303 4118 2307
rect 4121 2303 4125 2307
rect 6 2288 10 2292
rect 286 2288 290 2292
rect 446 2288 450 2292
rect 502 2288 506 2292
rect 542 2288 546 2292
rect 694 2288 698 2292
rect 822 2288 826 2292
rect 1046 2288 1050 2292
rect 1510 2288 1514 2292
rect 1574 2288 1578 2292
rect 1646 2288 1650 2292
rect 1702 2288 1706 2292
rect 1798 2288 1802 2292
rect 1814 2288 1818 2292
rect 1894 2288 1898 2292
rect 2102 2288 2106 2292
rect 2286 2288 2290 2292
rect 2318 2288 2322 2292
rect 2430 2288 2434 2292
rect 2502 2288 2506 2292
rect 2630 2288 2634 2292
rect 2694 2288 2698 2292
rect 2734 2288 2738 2292
rect 2790 2288 2794 2292
rect 2886 2288 2890 2292
rect 3070 2288 3074 2292
rect 3398 2288 3402 2292
rect 3558 2288 3562 2292
rect 3662 2288 3666 2292
rect 3822 2288 3826 2292
rect 3902 2288 3906 2292
rect 4054 2288 4058 2292
rect 4238 2288 4242 2292
rect 4326 2288 4330 2292
rect 4358 2288 4362 2292
rect 4398 2288 4402 2292
rect 4486 2288 4490 2292
rect 4510 2288 4514 2292
rect 4830 2288 4834 2292
rect 454 2278 458 2282
rect 470 2278 474 2282
rect 478 2278 482 2282
rect 1102 2278 1106 2282
rect 1206 2278 1210 2282
rect 1478 2278 1482 2282
rect 1806 2278 1810 2282
rect 1854 2278 1858 2282
rect 1950 2278 1954 2282
rect 1966 2278 1970 2282
rect 1998 2278 2002 2282
rect 2054 2278 2058 2282
rect 2238 2278 2242 2282
rect 2342 2278 2346 2282
rect 2902 2278 2906 2282
rect 2918 2278 2922 2282
rect 2926 2278 2930 2282
rect 2966 2278 2970 2282
rect 2974 2278 2978 2282
rect 2990 2278 2994 2282
rect 3014 2278 3018 2282
rect 3046 2278 3050 2282
rect 3382 2278 3386 2282
rect 3462 2278 3466 2282
rect 3550 2278 3554 2282
rect 3574 2278 3578 2282
rect 3846 2278 3850 2282
rect 3910 2278 3914 2282
rect 4318 2278 4322 2282
rect 4478 2278 4482 2282
rect 4590 2278 4594 2282
rect 4838 2278 4842 2282
rect 62 2268 66 2272
rect 102 2268 106 2272
rect 118 2268 122 2272
rect 158 2268 162 2272
rect 166 2268 170 2272
rect 294 2268 298 2272
rect 350 2268 354 2272
rect 390 2268 394 2272
rect 406 2268 410 2272
rect 518 2268 522 2272
rect 566 2268 570 2272
rect 582 2268 586 2272
rect 670 2268 674 2272
rect 702 2268 706 2272
rect 766 2268 770 2272
rect 830 2268 834 2272
rect 846 2268 850 2272
rect 902 2268 906 2272
rect 1110 2268 1114 2272
rect 1118 2268 1122 2272
rect 1150 2268 1154 2272
rect 1182 2268 1186 2272
rect 1230 2268 1234 2272
rect 1238 2268 1242 2272
rect 1294 2268 1298 2272
rect 1302 2268 1306 2272
rect 1326 2268 1330 2272
rect 1366 2268 1370 2272
rect 1486 2268 1490 2272
rect 1494 2268 1498 2272
rect 1518 2268 1522 2272
rect 1550 2268 1554 2272
rect 1654 2268 1658 2272
rect 1670 2268 1674 2272
rect 1686 2268 1690 2272
rect 1726 2268 1730 2272
rect 1750 2268 1754 2272
rect 1758 2268 1762 2272
rect 1838 2268 1842 2272
rect 1846 2268 1850 2272
rect 1862 2268 1866 2272
rect 1870 2268 1874 2272
rect 1902 2268 1906 2272
rect 1990 2268 1994 2272
rect 2014 2268 2018 2272
rect 2078 2268 2082 2272
rect 2158 2268 2162 2272
rect 2166 2268 2170 2272
rect 2230 2268 2234 2272
rect 2262 2268 2266 2272
rect 2326 2268 2330 2272
rect 2366 2268 2370 2272
rect 2446 2268 2450 2272
rect 2486 2268 2490 2272
rect 2518 2268 2522 2272
rect 2566 2268 2570 2272
rect 2766 2268 2770 2272
rect 2814 2268 2818 2272
rect 2894 2268 2898 2272
rect 2942 2268 2946 2272
rect 3182 2268 3186 2272
rect 3294 2268 3298 2272
rect 3342 2268 3346 2272
rect 3494 2268 3498 2272
rect 3542 2268 3546 2272
rect 3590 2268 3594 2272
rect 3678 2268 3682 2272
rect 3726 2268 3730 2272
rect 3782 2268 3786 2272
rect 3814 2268 3818 2272
rect 3838 2268 3842 2272
rect 3886 2268 3890 2272
rect 3998 2268 4002 2272
rect 4078 2268 4082 2272
rect 4158 2268 4162 2272
rect 4286 2268 4290 2272
rect 4294 2268 4298 2272
rect 4382 2268 4386 2272
rect 4422 2268 4426 2272
rect 4478 2268 4482 2272
rect 4502 2268 4506 2272
rect 4686 2268 4690 2272
rect 4734 2268 4738 2272
rect 4750 2268 4754 2272
rect 4854 2268 4858 2272
rect 4934 2268 4938 2272
rect 4942 2268 4946 2272
rect 5054 2268 5058 2272
rect 5070 2268 5074 2272
rect 5086 2268 5090 2272
rect 5118 2268 5122 2272
rect 5190 2268 5194 2272
rect 70 2259 74 2263
rect 110 2258 114 2262
rect 190 2258 194 2262
rect 230 2258 234 2262
rect 254 2258 258 2262
rect 302 2258 306 2262
rect 342 2258 346 2262
rect 382 2259 386 2263
rect 470 2258 474 2262
rect 486 2258 490 2262
rect 526 2258 530 2262
rect 598 2258 602 2262
rect 622 2258 626 2262
rect 630 2258 634 2262
rect 654 2258 658 2262
rect 678 2258 682 2262
rect 710 2258 714 2262
rect 782 2258 786 2262
rect 854 2258 858 2262
rect 894 2258 898 2262
rect 910 2258 914 2262
rect 918 2258 922 2262
rect 942 2258 946 2262
rect 982 2259 986 2263
rect 1006 2258 1010 2262
rect 1094 2258 1098 2262
rect 1118 2258 1122 2262
rect 1158 2258 1162 2262
rect 1190 2258 1194 2262
rect 1238 2258 1242 2262
rect 1294 2258 1298 2262
rect 1302 2258 1306 2262
rect 1334 2258 1338 2262
rect 1342 2258 1346 2262
rect 1374 2258 1378 2262
rect 1406 2259 1410 2263
rect 1430 2258 1434 2262
rect 1526 2258 1530 2262
rect 1550 2258 1554 2262
rect 1590 2258 1594 2262
rect 1598 2258 1602 2262
rect 1622 2258 1626 2262
rect 1662 2258 1666 2262
rect 1694 2258 1698 2262
rect 1718 2258 1722 2262
rect 1782 2258 1786 2262
rect 1790 2258 1794 2262
rect 1838 2258 1842 2262
rect 1870 2258 1874 2262
rect 1878 2258 1882 2262
rect 1910 2258 1914 2262
rect 1942 2258 1946 2262
rect 1966 2258 1970 2262
rect 1998 2258 2002 2262
rect 2014 2258 2018 2262
rect 2054 2258 2058 2262
rect 2070 2258 2074 2262
rect 2118 2258 2122 2262
rect 2158 2258 2162 2262
rect 2198 2258 2202 2262
rect 2206 2258 2210 2262
rect 2254 2258 2258 2262
rect 2270 2258 2274 2262
rect 2302 2258 2306 2262
rect 2350 2258 2354 2262
rect 2406 2258 2410 2262
rect 2510 2258 2514 2262
rect 2542 2258 2546 2262
rect 2646 2258 2650 2262
rect 2678 2258 2682 2262
rect 2710 2258 2714 2262
rect 2750 2258 2754 2262
rect 2806 2258 2810 2262
rect 2822 2258 2826 2262
rect 2846 2258 2850 2262
rect 2854 2258 2858 2262
rect 2902 2258 2906 2262
rect 2942 2258 2946 2262
rect 2974 2258 2978 2262
rect 2998 2258 3002 2262
rect 3030 2258 3034 2262
rect 3062 2258 3066 2262
rect 3086 2258 3090 2262
rect 3094 2258 3098 2262
rect 3102 2258 3106 2262
rect 3158 2258 3162 2262
rect 3174 2258 3178 2262
rect 3230 2258 3234 2262
rect 3262 2259 3266 2263
rect 3294 2258 3298 2262
rect 3358 2258 3362 2262
rect 3366 2258 3370 2262
rect 3462 2259 3466 2263
rect 3502 2258 3506 2262
rect 3566 2258 3570 2262
rect 3574 2258 3578 2262
rect 3638 2258 3642 2262
rect 3646 2258 3650 2262
rect 3726 2258 3730 2262
rect 3750 2258 3754 2262
rect 3758 2258 3762 2262
rect 3782 2258 3786 2262
rect 3806 2258 3810 2262
rect 3862 2258 3866 2262
rect 3894 2258 3898 2262
rect 3974 2258 3978 2262
rect 4046 2258 4050 2262
rect 4070 2258 4074 2262
rect 4198 2258 4202 2262
rect 4254 2258 4258 2262
rect 4278 2258 4282 2262
rect 4342 2258 4346 2262
rect 4414 2258 4418 2262
rect 4462 2258 4466 2262
rect 4502 2258 4506 2262
rect 4582 2258 4586 2262
rect 4638 2258 4642 2262
rect 4646 2258 4650 2262
rect 4670 2258 4674 2262
rect 4726 2258 4730 2262
rect 4766 2259 4770 2263
rect 4798 2258 4802 2262
rect 4862 2258 4866 2262
rect 4966 2258 4970 2262
rect 5006 2258 5010 2262
rect 5030 2258 5034 2262
rect 5078 2258 5082 2262
rect 134 2248 138 2252
rect 302 2248 306 2252
rect 326 2248 330 2252
rect 542 2248 546 2252
rect 574 2248 578 2252
rect 582 2248 586 2252
rect 614 2248 618 2252
rect 694 2248 698 2252
rect 710 2248 714 2252
rect 726 2248 730 2252
rect 870 2248 874 2252
rect 894 2248 898 2252
rect 1142 2248 1146 2252
rect 1158 2248 1162 2252
rect 1206 2248 1210 2252
rect 1214 2248 1218 2252
rect 1262 2248 1266 2252
rect 1286 2248 1290 2252
rect 1510 2248 1514 2252
rect 1542 2248 1546 2252
rect 1582 2248 1586 2252
rect 1638 2248 1642 2252
rect 1702 2248 1706 2252
rect 1734 2248 1738 2252
rect 1814 2248 1818 2252
rect 1974 2248 1978 2252
rect 2214 2248 2218 2252
rect 2502 2248 2506 2252
rect 2534 2248 2538 2252
rect 2550 2248 2554 2252
rect 3134 2248 3138 2252
rect 3150 2248 3154 2252
rect 3302 2248 3306 2252
rect 3326 2248 3330 2252
rect 3350 2248 3354 2252
rect 3390 2248 3394 2252
rect 3526 2248 3530 2252
rect 3766 2248 3770 2252
rect 3790 2248 3794 2252
rect 3822 2248 3826 2252
rect 4262 2248 4266 2252
rect 4294 2248 4298 2252
rect 4318 2248 4322 2252
rect 4366 2248 4370 2252
rect 4438 2248 4442 2252
rect 4702 2248 4706 2252
rect 5094 2248 5098 2252
rect 5102 2248 5106 2252
rect 1078 2238 1082 2242
rect 1174 2238 1178 2242
rect 1454 2238 1458 2242
rect 1750 2238 1754 2242
rect 2134 2238 2138 2242
rect 2886 2238 2890 2242
rect 3502 2238 3506 2242
rect 3870 2238 3874 2242
rect 3918 2238 3922 2242
rect 3934 2238 3938 2242
rect 4462 2238 4466 2242
rect 3014 2228 3018 2232
rect 3558 2228 3562 2232
rect 4214 2228 4218 2232
rect 598 2218 602 2222
rect 646 2218 650 2222
rect 838 2218 842 2222
rect 934 2218 938 2222
rect 1126 2218 1130 2222
rect 1222 2218 1226 2222
rect 1310 2218 1314 2222
rect 1366 2218 1370 2222
rect 1614 2218 1618 2222
rect 1686 2218 1690 2222
rect 1926 2218 1930 2222
rect 1958 2218 1962 2222
rect 2062 2218 2066 2222
rect 2390 2218 2394 2222
rect 2430 2218 2434 2222
rect 2470 2218 2474 2222
rect 2598 2218 2602 2222
rect 2662 2218 2666 2222
rect 2734 2218 2738 2222
rect 2790 2218 2794 2222
rect 2966 2218 2970 2222
rect 3030 2218 3034 2222
rect 3702 2218 3706 2222
rect 3774 2218 3778 2222
rect 4022 2218 4026 2222
rect 4054 2218 4058 2222
rect 4174 2218 4178 2222
rect 4278 2218 4282 2222
rect 4398 2218 4402 2222
rect 4662 2218 4666 2222
rect 4726 2218 4730 2222
rect 4838 2218 4842 2222
rect 4878 2218 4882 2222
rect 5110 2218 5114 2222
rect 5134 2218 5138 2222
rect 538 2203 542 2207
rect 545 2203 549 2207
rect 1562 2203 1566 2207
rect 1569 2203 1573 2207
rect 2586 2203 2590 2207
rect 2593 2203 2597 2207
rect 3610 2203 3614 2207
rect 3617 2203 3621 2207
rect 4634 2203 4638 2207
rect 4641 2203 4645 2207
rect 374 2188 378 2192
rect 622 2188 626 2192
rect 638 2188 642 2192
rect 686 2188 690 2192
rect 1302 2188 1306 2192
rect 1342 2188 1346 2192
rect 1934 2188 1938 2192
rect 2182 2188 2186 2192
rect 2318 2188 2322 2192
rect 2350 2188 2354 2192
rect 3054 2188 3058 2192
rect 3150 2188 3154 2192
rect 3470 2188 3474 2192
rect 3742 2188 3746 2192
rect 4086 2188 4090 2192
rect 4206 2188 4210 2192
rect 4326 2188 4330 2192
rect 4806 2188 4810 2192
rect 918 2178 922 2182
rect 1246 2178 1250 2182
rect 2590 2178 2594 2182
rect 3398 2178 3402 2182
rect 3630 2178 3634 2182
rect 3718 2178 3722 2182
rect 4686 2178 4690 2182
rect 214 2168 218 2172
rect 254 2168 258 2172
rect 470 2168 474 2172
rect 510 2168 514 2172
rect 582 2168 586 2172
rect 798 2168 802 2172
rect 1086 2168 1090 2172
rect 1390 2168 1394 2172
rect 3166 2168 3170 2172
rect 3406 2168 3410 2172
rect 3678 2168 3682 2172
rect 3886 2168 3890 2172
rect 4062 2168 4066 2172
rect 4886 2168 4890 2172
rect 4982 2168 4986 2172
rect 62 2148 66 2152
rect 94 2147 98 2151
rect 158 2148 162 2152
rect 230 2148 234 2152
rect 238 2148 242 2152
rect 270 2148 274 2152
rect 310 2147 314 2151
rect 414 2148 418 2152
rect 486 2148 490 2152
rect 494 2148 498 2152
rect 590 2158 594 2162
rect 614 2158 618 2162
rect 526 2148 530 2152
rect 638 2148 642 2152
rect 670 2148 674 2152
rect 694 2148 698 2152
rect 702 2148 706 2152
rect 742 2148 746 2152
rect 766 2148 770 2152
rect 814 2148 818 2152
rect 822 2148 826 2152
rect 838 2158 842 2162
rect 886 2158 890 2162
rect 910 2158 914 2162
rect 926 2158 930 2162
rect 854 2148 858 2152
rect 966 2158 970 2162
rect 1150 2158 1154 2162
rect 1254 2158 1258 2162
rect 1422 2158 1426 2162
rect 942 2148 946 2152
rect 958 2148 962 2152
rect 974 2148 978 2152
rect 982 2148 986 2152
rect 1022 2147 1026 2151
rect 1134 2148 1138 2152
rect 1182 2147 1186 2151
rect 1278 2148 1282 2152
rect 1286 2148 1290 2152
rect 1310 2148 1314 2152
rect 1334 2148 1338 2152
rect 1358 2148 1362 2152
rect 1366 2148 1370 2152
rect 1382 2148 1386 2152
rect 1406 2148 1410 2152
rect 1414 2148 1418 2152
rect 1446 2148 1450 2152
rect 1462 2148 1466 2152
rect 1502 2148 1506 2152
rect 1526 2158 1530 2162
rect 1662 2158 1666 2162
rect 1686 2158 1690 2162
rect 1902 2158 1906 2162
rect 1598 2148 1602 2152
rect 1622 2148 1626 2152
rect 1710 2148 1714 2152
rect 1734 2148 1738 2152
rect 1742 2148 1746 2152
rect 1774 2148 1778 2152
rect 1830 2148 1834 2152
rect 6 2138 10 2142
rect 222 2138 226 2142
rect 278 2138 282 2142
rect 294 2138 298 2142
rect 390 2138 394 2142
rect 478 2138 482 2142
rect 558 2138 562 2142
rect 606 2138 610 2142
rect 630 2138 634 2142
rect 718 2138 722 2142
rect 806 2138 810 2142
rect 862 2138 866 2142
rect 870 2138 874 2142
rect 910 2138 914 2142
rect 934 2138 938 2142
rect 958 2138 962 2142
rect 990 2138 994 2142
rect 1006 2138 1010 2142
rect 1126 2138 1130 2142
rect 1142 2138 1146 2142
rect 1166 2138 1170 2142
rect 1270 2138 1274 2142
rect 1438 2138 1442 2142
rect 1526 2138 1530 2142
rect 1542 2138 1546 2142
rect 1678 2138 1682 2142
rect 1862 2147 1866 2151
rect 1902 2148 1906 2152
rect 1926 2158 1930 2162
rect 1990 2158 1994 2162
rect 2046 2158 2050 2162
rect 2086 2158 2090 2162
rect 2166 2158 2170 2162
rect 2334 2158 2338 2162
rect 2366 2158 2370 2162
rect 1926 2148 1930 2152
rect 1950 2148 1954 2152
rect 1982 2148 1986 2152
rect 2038 2148 2042 2152
rect 2102 2148 2106 2152
rect 2142 2148 2146 2152
rect 2174 2148 2178 2152
rect 2206 2148 2210 2152
rect 2230 2148 2234 2152
rect 2270 2148 2274 2152
rect 2294 2148 2298 2152
rect 2302 2148 2306 2152
rect 2350 2148 2354 2152
rect 2438 2148 2442 2152
rect 2478 2148 2482 2152
rect 2494 2148 2498 2152
rect 2510 2158 2514 2162
rect 3006 2158 3010 2162
rect 3062 2158 3066 2162
rect 3382 2158 3386 2162
rect 3422 2158 3426 2162
rect 3438 2158 3442 2162
rect 2622 2148 2626 2152
rect 2646 2148 2650 2152
rect 2718 2148 2722 2152
rect 2782 2148 2786 2152
rect 2886 2148 2890 2152
rect 1750 2138 1754 2142
rect 1766 2138 1770 2142
rect 1790 2138 1794 2142
rect 1894 2138 1898 2142
rect 1942 2138 1946 2142
rect 1958 2138 1962 2142
rect 1974 2138 1978 2142
rect 2006 2138 2010 2142
rect 2070 2138 2074 2142
rect 2118 2138 2122 2142
rect 2126 2138 2130 2142
rect 2134 2138 2138 2142
rect 2150 2138 2154 2142
rect 2198 2138 2202 2142
rect 2278 2138 2282 2142
rect 2446 2138 2450 2142
rect 2478 2138 2482 2142
rect 2526 2138 2530 2142
rect 2534 2138 2538 2142
rect 2918 2148 2922 2152
rect 2926 2148 2930 2152
rect 2958 2148 2962 2152
rect 2982 2148 2986 2152
rect 2998 2148 3002 2152
rect 3022 2148 3026 2152
rect 3102 2148 3106 2152
rect 3134 2148 3138 2152
rect 3222 2148 3226 2152
rect 3262 2148 3266 2152
rect 3310 2148 3314 2152
rect 3318 2148 3322 2152
rect 3350 2148 3354 2152
rect 3366 2148 3370 2152
rect 3398 2148 3402 2152
rect 3446 2148 3450 2152
rect 3454 2148 3458 2152
rect 3478 2148 3482 2152
rect 3486 2148 3490 2152
rect 3510 2148 3514 2152
rect 3550 2148 3554 2152
rect 3574 2158 3578 2162
rect 3726 2158 3730 2162
rect 3614 2148 3618 2152
rect 3622 2148 3626 2152
rect 3646 2148 3650 2152
rect 3654 2148 3658 2152
rect 3670 2148 3674 2152
rect 3694 2148 3698 2152
rect 3742 2148 3746 2152
rect 3766 2148 3770 2152
rect 3790 2158 3794 2162
rect 3814 2158 3818 2162
rect 3862 2158 3866 2162
rect 3838 2148 3842 2152
rect 3910 2158 3914 2162
rect 4150 2158 4154 2162
rect 4230 2158 4234 2162
rect 4302 2158 4306 2162
rect 4638 2158 4642 2162
rect 4734 2158 4738 2162
rect 3886 2148 3890 2152
rect 3974 2148 3978 2152
rect 4022 2148 4026 2152
rect 4038 2148 4042 2152
rect 4078 2148 4082 2152
rect 4102 2148 4106 2152
rect 4110 2148 4114 2152
rect 4142 2148 4146 2152
rect 4166 2148 4170 2152
rect 4174 2148 4178 2152
rect 4190 2148 4194 2152
rect 4214 2148 4218 2152
rect 4222 2148 4226 2152
rect 4254 2148 4258 2152
rect 4286 2148 4290 2152
rect 4342 2148 4346 2152
rect 4350 2148 4354 2152
rect 2758 2138 2762 2142
rect 2862 2138 2866 2142
rect 2894 2138 2898 2142
rect 2926 2138 2930 2142
rect 2934 2138 2938 2142
rect 2942 2138 2946 2142
rect 2950 2138 2954 2142
rect 2974 2138 2978 2142
rect 2990 2138 2994 2142
rect 3022 2138 3026 2142
rect 3038 2138 3042 2142
rect 3054 2138 3058 2142
rect 3078 2138 3082 2142
rect 3086 2138 3090 2142
rect 3134 2138 3138 2142
rect 3142 2138 3146 2142
rect 3230 2138 3234 2142
rect 3270 2138 3274 2142
rect 3326 2138 3330 2142
rect 3342 2138 3346 2142
rect 3358 2138 3362 2142
rect 3422 2138 3426 2142
rect 3494 2138 3498 2142
rect 3590 2138 3594 2142
rect 3750 2138 3754 2142
rect 3774 2138 3778 2142
rect 3806 2138 3810 2142
rect 3822 2138 3826 2142
rect 3838 2138 3842 2142
rect 3846 2138 3850 2142
rect 3998 2138 4002 2142
rect 4014 2138 4018 2142
rect 4446 2147 4450 2151
rect 4478 2148 4482 2152
rect 4494 2148 4498 2152
rect 4526 2148 4530 2152
rect 4582 2148 4586 2152
rect 4662 2148 4666 2152
rect 4702 2148 4706 2152
rect 4710 2148 4714 2152
rect 4790 2158 4794 2162
rect 4846 2158 4850 2162
rect 4750 2148 4754 2152
rect 4758 2148 4762 2152
rect 4766 2148 4770 2152
rect 4806 2148 4810 2152
rect 4918 2148 4922 2152
rect 4998 2148 5002 2152
rect 5022 2148 5026 2152
rect 5086 2148 5090 2152
rect 5134 2148 5138 2152
rect 5150 2148 5154 2152
rect 4046 2138 4050 2142
rect 4358 2138 4362 2142
rect 4374 2138 4378 2142
rect 4462 2138 4466 2142
rect 4486 2138 4490 2142
rect 4590 2138 4594 2142
rect 4662 2138 4666 2142
rect 4718 2138 4722 2142
rect 4774 2138 4778 2142
rect 4798 2138 4802 2142
rect 4830 2138 4834 2142
rect 4854 2138 4858 2142
rect 4950 2138 4954 2142
rect 182 2128 186 2132
rect 374 2128 378 2132
rect 654 2128 658 2132
rect 894 2128 898 2132
rect 1118 2128 1122 2132
rect 1486 2128 1490 2132
rect 1670 2128 1674 2132
rect 1966 2128 1970 2132
rect 2094 2128 2098 2132
rect 2214 2128 2218 2132
rect 2838 2128 2842 2132
rect 2870 2128 2874 2132
rect 3054 2128 3058 2132
rect 3110 2128 3114 2132
rect 3294 2128 3298 2132
rect 3526 2128 3530 2132
rect 3710 2128 3714 2132
rect 4262 2128 4266 2132
rect 4414 2128 4418 2132
rect 4510 2128 4514 2132
rect 582 2118 586 2122
rect 598 2118 602 2122
rect 886 2118 890 2122
rect 1102 2118 1106 2122
rect 1246 2118 1250 2122
rect 1254 2118 1258 2122
rect 1558 2118 1562 2122
rect 1694 2118 1698 2122
rect 1718 2118 1722 2122
rect 1750 2118 1754 2122
rect 1990 2118 1994 2122
rect 2022 2118 2026 2122
rect 2046 2118 2050 2122
rect 2222 2118 2226 2122
rect 2246 2118 2250 2122
rect 2638 2118 2642 2122
rect 2670 2118 2674 2122
rect 2702 2118 2706 2122
rect 2734 2118 2738 2122
rect 2846 2118 2850 2122
rect 3006 2118 3010 2122
rect 3278 2118 3282 2122
rect 3326 2118 3330 2122
rect 3566 2118 3570 2122
rect 4230 2118 4234 2122
rect 4534 2118 4538 2122
rect 4646 2118 4650 2122
rect 4790 2118 4794 2122
rect 4966 2118 4970 2122
rect 5070 2118 5074 2122
rect 5094 2118 5098 2122
rect 1050 2103 1054 2107
rect 1057 2103 1061 2107
rect 2074 2103 2078 2107
rect 2081 2103 2085 2107
rect 3098 2103 3102 2107
rect 3105 2103 3109 2107
rect 4114 2103 4118 2107
rect 4121 2103 4125 2107
rect 6 2088 10 2092
rect 118 2088 122 2092
rect 230 2088 234 2092
rect 326 2088 330 2092
rect 422 2088 426 2092
rect 814 2088 818 2092
rect 854 2088 858 2092
rect 1222 2088 1226 2092
rect 1462 2088 1466 2092
rect 1510 2088 1514 2092
rect 1534 2088 1538 2092
rect 1582 2088 1586 2092
rect 1694 2088 1698 2092
rect 1806 2088 1810 2092
rect 1886 2088 1890 2092
rect 2014 2088 2018 2092
rect 2094 2088 2098 2092
rect 2214 2088 2218 2092
rect 2262 2088 2266 2092
rect 2294 2088 2298 2092
rect 2334 2088 2338 2092
rect 2462 2088 2466 2092
rect 2518 2088 2522 2092
rect 2558 2088 2562 2092
rect 2710 2088 2714 2092
rect 3286 2088 3290 2092
rect 3446 2088 3450 2092
rect 3486 2088 3490 2092
rect 3502 2088 3506 2092
rect 3702 2088 3706 2092
rect 3726 2088 3730 2092
rect 3886 2088 3890 2092
rect 3966 2088 3970 2092
rect 4166 2088 4170 2092
rect 4174 2088 4178 2092
rect 4518 2088 4522 2092
rect 4582 2088 4586 2092
rect 4614 2088 4618 2092
rect 4822 2088 4826 2092
rect 4990 2088 4994 2092
rect 5054 2088 5058 2092
rect 5118 2088 5122 2092
rect 150 2078 154 2082
rect 158 2078 162 2082
rect 222 2078 226 2082
rect 526 2078 530 2082
rect 1270 2078 1274 2082
rect 1630 2078 1634 2082
rect 2222 2078 2226 2082
rect 2230 2078 2234 2082
rect 2438 2078 2442 2082
rect 2502 2078 2506 2082
rect 2910 2078 2914 2082
rect 3254 2078 3258 2082
rect 3262 2078 3266 2082
rect 3382 2078 3386 2082
rect 3862 2078 3866 2082
rect 3910 2078 3914 2082
rect 4126 2078 4130 2082
rect 86 2068 90 2072
rect 110 2068 114 2072
rect 182 2068 186 2072
rect 214 2068 218 2072
rect 262 2068 266 2072
rect 342 2068 346 2072
rect 390 2068 394 2072
rect 430 2068 434 2072
rect 462 2068 466 2072
rect 494 2068 498 2072
rect 686 2068 690 2072
rect 702 2068 706 2072
rect 718 2068 722 2072
rect 750 2068 754 2072
rect 766 2068 770 2072
rect 774 2068 778 2072
rect 822 2068 826 2072
rect 870 2068 874 2072
rect 886 2068 890 2072
rect 974 2068 978 2072
rect 1030 2068 1034 2072
rect 1054 2068 1058 2072
rect 1102 2068 1106 2072
rect 1150 2068 1154 2072
rect 1190 2068 1194 2072
rect 1238 2068 1242 2072
rect 1310 2068 1314 2072
rect 1326 2068 1330 2072
rect 1342 2068 1346 2072
rect 1366 2068 1370 2072
rect 1486 2068 1490 2072
rect 1502 2068 1506 2072
rect 1518 2068 1522 2072
rect 1550 2068 1554 2072
rect 1582 2068 1586 2072
rect 1598 2068 1602 2072
rect 1662 2068 1666 2072
rect 1710 2068 1714 2072
rect 1742 2068 1746 2072
rect 1750 2068 1754 2072
rect 1782 2068 1786 2072
rect 1798 2068 1802 2072
rect 1814 2068 1818 2072
rect 1926 2068 1930 2072
rect 1934 2068 1938 2072
rect 2086 2068 2090 2072
rect 2094 2068 2098 2072
rect 2110 2068 2114 2072
rect 2238 2068 2242 2072
rect 2318 2068 2322 2072
rect 2382 2068 2386 2072
rect 2422 2068 2426 2072
rect 2486 2068 2490 2072
rect 2518 2068 2522 2072
rect 2534 2068 2538 2072
rect 2542 2068 2546 2072
rect 2590 2068 2594 2072
rect 2630 2068 2634 2072
rect 2718 2068 2722 2072
rect 2766 2068 2770 2072
rect 2790 2068 2794 2072
rect 2798 2068 2802 2072
rect 2822 2068 2826 2072
rect 2878 2068 2882 2072
rect 2982 2068 2986 2072
rect 3030 2068 3034 2072
rect 3078 2068 3082 2072
rect 3126 2068 3130 2072
rect 3142 2068 3146 2072
rect 3334 2068 3338 2072
rect 3422 2068 3426 2072
rect 3446 2068 3450 2072
rect 3462 2068 3466 2072
rect 3478 2068 3482 2072
rect 3710 2068 3714 2072
rect 3726 2068 3730 2072
rect 3870 2068 3874 2072
rect 3902 2068 3906 2072
rect 3950 2068 3954 2072
rect 4062 2068 4066 2072
rect 4086 2068 4090 2072
rect 4134 2068 4138 2072
rect 4294 2068 4298 2072
rect 4382 2068 4386 2072
rect 4406 2068 4410 2072
rect 4430 2068 4434 2072
rect 4438 2068 4442 2072
rect 4470 2068 4474 2072
rect 4494 2068 4498 2072
rect 4526 2068 4530 2072
rect 4542 2068 4546 2072
rect 4958 2078 4962 2082
rect 5086 2078 5090 2082
rect 5190 2078 5194 2082
rect 4590 2068 4594 2072
rect 4606 2068 4610 2072
rect 4670 2068 4674 2072
rect 4782 2068 4786 2072
rect 4918 2068 4922 2072
rect 4934 2068 4938 2072
rect 4998 2068 5002 2072
rect 5014 2068 5018 2072
rect 5046 2068 5050 2072
rect 5094 2068 5098 2072
rect 5142 2068 5146 2072
rect 5174 2068 5178 2072
rect 70 2059 74 2063
rect 102 2058 106 2062
rect 134 2058 138 2062
rect 174 2058 178 2062
rect 222 2058 226 2062
rect 270 2058 274 2062
rect 366 2058 370 2062
rect 438 2058 442 2062
rect 470 2058 474 2062
rect 502 2058 506 2062
rect 566 2058 570 2062
rect 622 2058 626 2062
rect 646 2058 650 2062
rect 694 2058 698 2062
rect 718 2058 722 2062
rect 734 2058 738 2062
rect 766 2058 770 2062
rect 782 2058 786 2062
rect 798 2058 802 2062
rect 830 2058 834 2062
rect 838 2058 842 2062
rect 862 2058 866 2062
rect 910 2058 914 2062
rect 982 2058 986 2062
rect 1022 2058 1026 2062
rect 1094 2058 1098 2062
rect 1110 2058 1114 2062
rect 1118 2058 1122 2062
rect 1142 2058 1146 2062
rect 1158 2058 1162 2062
rect 1166 2058 1170 2062
rect 1190 2058 1194 2062
rect 1206 2058 1210 2062
rect 1238 2058 1242 2062
rect 1262 2058 1266 2062
rect 1294 2058 1298 2062
rect 1302 2058 1306 2062
rect 1310 2058 1314 2062
rect 1350 2058 1354 2062
rect 1382 2059 1386 2063
rect 1494 2058 1498 2062
rect 1534 2058 1538 2062
rect 1574 2058 1578 2062
rect 1606 2058 1610 2062
rect 1614 2058 1618 2062
rect 1622 2058 1626 2062
rect 1646 2058 1650 2062
rect 1686 2058 1690 2062
rect 1742 2058 1746 2062
rect 1782 2058 1786 2062
rect 1790 2058 1794 2062
rect 1822 2058 1826 2062
rect 1838 2058 1842 2062
rect 1862 2058 1866 2062
rect 1870 2058 1874 2062
rect 1910 2058 1914 2062
rect 1974 2058 1978 2062
rect 2038 2058 2042 2062
rect 2062 2058 2066 2062
rect 2118 2058 2122 2062
rect 2158 2058 2162 2062
rect 2182 2058 2186 2062
rect 2246 2058 2250 2062
rect 2278 2058 2282 2062
rect 2310 2058 2314 2062
rect 2342 2058 2346 2062
rect 2350 2058 2354 2062
rect 2374 2058 2378 2062
rect 2382 2058 2386 2062
rect 2398 2058 2402 2062
rect 2438 2058 2442 2062
rect 2462 2058 2466 2062
rect 2510 2058 2514 2062
rect 2542 2058 2546 2062
rect 2550 2058 2554 2062
rect 2582 2058 2586 2062
rect 2654 2058 2658 2062
rect 2758 2058 2762 2062
rect 2822 2058 2826 2062
rect 2830 2058 2834 2062
rect 2870 2058 2874 2062
rect 2910 2059 2914 2063
rect 2998 2058 3002 2062
rect 3038 2058 3042 2062
rect 3062 2058 3066 2062
rect 3070 2058 3074 2062
rect 3142 2058 3146 2062
rect 3182 2058 3186 2062
rect 3206 2058 3210 2062
rect 3278 2058 3282 2062
rect 3350 2059 3354 2063
rect 3398 2058 3402 2062
rect 3430 2058 3434 2062
rect 3438 2058 3442 2062
rect 3470 2058 3474 2062
rect 3566 2059 3570 2063
rect 3646 2058 3650 2062
rect 3670 2058 3674 2062
rect 3782 2058 3786 2062
rect 3790 2058 3794 2062
rect 3846 2058 3850 2062
rect 3878 2058 3882 2062
rect 3926 2058 3930 2062
rect 3942 2058 3946 2062
rect 3958 2058 3962 2062
rect 3998 2058 4002 2062
rect 4022 2058 4026 2062
rect 4078 2058 4082 2062
rect 4110 2058 4114 2062
rect 4230 2058 4234 2062
rect 4302 2058 4306 2062
rect 4390 2058 4394 2062
rect 4446 2058 4450 2062
rect 4502 2058 4506 2062
rect 4566 2058 4570 2062
rect 4598 2058 4602 2062
rect 4670 2058 4674 2062
rect 4702 2059 4706 2063
rect 4734 2058 4738 2062
rect 4806 2058 4810 2062
rect 4894 2058 4898 2062
rect 4974 2058 4978 2062
rect 5006 2058 5010 2062
rect 5038 2058 5042 2062
rect 5070 2058 5074 2062
rect 5134 2058 5138 2062
rect 5142 2058 5146 2062
rect 5174 2058 5178 2062
rect 158 2048 162 2052
rect 190 2048 194 2052
rect 454 2048 458 2052
rect 470 2048 474 2052
rect 486 2048 490 2052
rect 502 2048 506 2052
rect 526 2048 530 2052
rect 582 2048 586 2052
rect 710 2048 714 2052
rect 750 2048 754 2052
rect 798 2048 802 2052
rect 806 2048 810 2052
rect 1038 2048 1042 2052
rect 1286 2048 1290 2052
rect 1534 2048 1538 2052
rect 1678 2048 1682 2052
rect 1726 2048 1730 2052
rect 1846 2048 1850 2052
rect 2334 2048 2338 2052
rect 2734 2048 2738 2052
rect 2774 2048 2778 2052
rect 2814 2048 2818 2052
rect 2846 2048 2850 2052
rect 2854 2048 2858 2052
rect 2870 2048 2874 2052
rect 3094 2048 3098 2052
rect 3270 2048 3274 2052
rect 3494 2048 3498 2052
rect 3726 2048 3730 2052
rect 3886 2048 3890 2052
rect 4166 2048 4170 2052
rect 4414 2048 4418 2052
rect 4486 2048 4490 2052
rect 4542 2048 4546 2052
rect 4622 2048 4626 2052
rect 4646 2048 4650 2052
rect 4662 2048 4666 2052
rect 4790 2048 4794 2052
rect 4806 2048 4810 2052
rect 4950 2048 4954 2052
rect 5110 2048 5114 2052
rect 5150 2048 5154 2052
rect 206 2038 210 2042
rect 438 2038 442 2042
rect 678 2038 682 2042
rect 966 2038 970 2042
rect 1006 2038 1010 2042
rect 1094 2038 1098 2042
rect 1270 2038 1274 2042
rect 1430 2038 1434 2042
rect 1446 2038 1450 2042
rect 3406 2038 3410 2042
rect 3982 2038 3986 2042
rect 4446 2038 4450 2042
rect 4942 2038 4946 2042
rect 5030 2038 5034 2042
rect 982 2028 986 2032
rect 566 2018 570 2022
rect 1278 2018 1282 2022
rect 1342 2018 1346 2022
rect 1758 2018 1762 2022
rect 1990 2018 1994 2022
rect 2014 2018 2018 2022
rect 2054 2018 2058 2022
rect 2294 2018 2298 2022
rect 2758 2018 2762 2022
rect 2782 2018 2786 2022
rect 2830 2018 2834 2022
rect 3054 2018 3058 2022
rect 3822 2018 3826 2022
rect 4070 2018 4074 2022
rect 4102 2018 4106 2022
rect 5022 2018 5026 2022
rect 538 2003 542 2007
rect 545 2003 549 2007
rect 1562 2003 1566 2007
rect 1569 2003 1573 2007
rect 2586 2003 2590 2007
rect 2593 2003 2597 2007
rect 3610 2003 3614 2007
rect 3617 2003 3621 2007
rect 4634 2003 4638 2007
rect 4641 2003 4645 2007
rect 62 1988 66 1992
rect 134 1988 138 1992
rect 862 1988 866 1992
rect 1014 1988 1018 1992
rect 1134 1988 1138 1992
rect 1182 1988 1186 1992
rect 1382 1988 1386 1992
rect 1510 1988 1514 1992
rect 1790 1988 1794 1992
rect 2038 1988 2042 1992
rect 2102 1988 2106 1992
rect 2142 1988 2146 1992
rect 2174 1988 2178 1992
rect 2214 1988 2218 1992
rect 2518 1988 2522 1992
rect 2686 1988 2690 1992
rect 2734 1988 2738 1992
rect 3446 1988 3450 1992
rect 3646 1988 3650 1992
rect 3686 1988 3690 1992
rect 3798 1988 3802 1992
rect 3878 1988 3882 1992
rect 4118 1988 4122 1992
rect 4390 1988 4394 1992
rect 4518 1988 4522 1992
rect 4718 1988 4722 1992
rect 5182 1988 5186 1992
rect 254 1978 258 1982
rect 2246 1978 2250 1982
rect 4886 1978 4890 1982
rect 238 1968 242 1972
rect 278 1968 282 1972
rect 598 1968 602 1972
rect 638 1968 642 1972
rect 798 1968 802 1972
rect 1310 1968 1314 1972
rect 2014 1968 2018 1972
rect 2294 1968 2298 1972
rect 2310 1968 2314 1972
rect 2774 1968 2778 1972
rect 3158 1968 3162 1972
rect 3766 1968 3770 1972
rect 3814 1968 3818 1972
rect 4350 1968 4354 1972
rect 4470 1968 4474 1972
rect 4782 1968 4786 1972
rect 5022 1968 5026 1972
rect 182 1948 186 1952
rect 246 1948 250 1952
rect 486 1958 490 1962
rect 614 1958 618 1962
rect 294 1948 298 1952
rect 342 1948 346 1952
rect 422 1948 426 1952
rect 454 1948 458 1952
rect 470 1948 474 1952
rect 494 1948 498 1952
rect 542 1948 546 1952
rect 614 1948 618 1952
rect 766 1958 770 1962
rect 654 1948 658 1952
rect 702 1948 706 1952
rect 790 1948 794 1952
rect 822 1958 826 1962
rect 918 1958 922 1962
rect 958 1958 962 1962
rect 966 1958 970 1962
rect 1038 1958 1042 1962
rect 1246 1958 1250 1962
rect 854 1948 858 1952
rect 878 1948 882 1952
rect 886 1948 890 1952
rect 894 1948 898 1952
rect 902 1948 906 1952
rect 926 1948 930 1952
rect 990 1948 994 1952
rect 998 1948 1002 1952
rect 1030 1948 1034 1952
rect 1102 1948 1106 1952
rect 1110 1948 1114 1952
rect 1118 1948 1122 1952
rect 1142 1948 1146 1952
rect 1158 1948 1162 1952
rect 1166 1948 1170 1952
rect 1190 1948 1194 1952
rect 1230 1948 1234 1952
rect 1286 1948 1290 1952
rect 1294 1948 1298 1952
rect 1310 1948 1314 1952
rect 1334 1958 1338 1962
rect 1358 1948 1362 1952
rect 1366 1948 1370 1952
rect 1390 1948 1394 1952
rect 1430 1948 1434 1952
rect 1454 1958 1458 1962
rect 1502 1948 1506 1952
rect 1566 1948 1570 1952
rect 1662 1948 1666 1952
rect 1686 1947 1690 1951
rect 1726 1948 1730 1952
rect 1734 1948 1738 1952
rect 1750 1958 1754 1962
rect 1822 1958 1826 1962
rect 1870 1958 1874 1962
rect 1774 1948 1778 1952
rect 1782 1948 1786 1952
rect 1838 1948 1842 1952
rect 1894 1958 1898 1962
rect 2542 1958 2546 1962
rect 2566 1958 2570 1962
rect 2662 1958 2666 1962
rect 2758 1958 2762 1962
rect 2982 1958 2986 1962
rect 3110 1958 3114 1962
rect 3230 1958 3234 1962
rect 3350 1958 3354 1962
rect 1902 1948 1906 1952
rect 1950 1947 1954 1951
rect 1982 1948 1986 1952
rect 2022 1948 2026 1952
rect 2030 1948 2034 1952
rect 2054 1948 2058 1952
rect 2070 1948 2074 1952
rect 2094 1948 2098 1952
rect 2126 1948 2130 1952
rect 2158 1948 2162 1952
rect 2198 1948 2202 1952
rect 2230 1948 2234 1952
rect 2286 1948 2290 1952
rect 2358 1947 2362 1951
rect 2406 1948 2410 1952
rect 2438 1948 2442 1952
rect 2454 1948 2458 1952
rect 2478 1948 2482 1952
rect 2486 1948 2490 1952
rect 2494 1948 2498 1952
rect 2502 1948 2506 1952
rect 2526 1948 2530 1952
rect 2638 1948 2642 1952
rect 2646 1948 2650 1952
rect 2702 1948 2706 1952
rect 2710 1948 2714 1952
rect 2718 1948 2722 1952
rect 2806 1948 2810 1952
rect 6 1938 10 1942
rect 78 1938 82 1942
rect 182 1938 186 1942
rect 246 1938 250 1942
rect 302 1938 306 1942
rect 446 1938 450 1942
rect 462 1938 466 1942
rect 518 1938 522 1942
rect 606 1938 610 1942
rect 662 1938 666 1942
rect 678 1938 682 1942
rect 782 1938 786 1942
rect 790 1938 794 1942
rect 838 1938 842 1942
rect 934 1938 938 1942
rect 982 1938 986 1942
rect 1054 1938 1058 1942
rect 1302 1938 1306 1942
rect 1350 1938 1354 1942
rect 1454 1938 1458 1942
rect 1470 1938 1474 1942
rect 1590 1938 1594 1942
rect 1718 1938 1722 1942
rect 1766 1938 1770 1942
rect 1846 1938 1850 1942
rect 1854 1938 1858 1942
rect 1902 1938 1906 1942
rect 2414 1938 2418 1942
rect 2430 1938 2434 1942
rect 2558 1938 2562 1942
rect 2582 1938 2586 1942
rect 2638 1938 2642 1942
rect 2838 1947 2842 1951
rect 2886 1948 2890 1952
rect 2918 1948 2922 1952
rect 2942 1948 2946 1952
rect 2974 1948 2978 1952
rect 3030 1947 3034 1951
rect 3102 1948 3106 1952
rect 3134 1948 3138 1952
rect 3174 1948 3178 1952
rect 3230 1948 3234 1952
rect 2750 1938 2754 1942
rect 2894 1938 2898 1942
rect 2910 1938 2914 1942
rect 2966 1938 2970 1942
rect 2998 1938 3002 1942
rect 3150 1938 3154 1942
rect 3214 1938 3218 1942
rect 3318 1947 3322 1951
rect 3382 1948 3386 1952
rect 3406 1958 3410 1962
rect 3606 1958 3610 1962
rect 3782 1958 3786 1962
rect 3830 1958 3834 1962
rect 3838 1958 3842 1962
rect 3894 1958 3898 1962
rect 3910 1958 3914 1962
rect 4022 1958 4026 1962
rect 3438 1948 3442 1952
rect 3462 1948 3466 1952
rect 3470 1948 3474 1952
rect 3478 1948 3482 1952
rect 3486 1948 3490 1952
rect 3502 1948 3506 1952
rect 3510 1948 3514 1952
rect 3518 1948 3522 1952
rect 3558 1948 3562 1952
rect 3574 1948 3578 1952
rect 3590 1948 3594 1952
rect 3622 1948 3626 1952
rect 3630 1948 3634 1952
rect 3662 1948 3666 1952
rect 3670 1948 3674 1952
rect 3718 1948 3722 1952
rect 3742 1948 3746 1952
rect 3750 1948 3754 1952
rect 3766 1948 3770 1952
rect 3806 1948 3810 1952
rect 3862 1948 3866 1952
rect 3918 1948 3922 1952
rect 3334 1938 3338 1942
rect 3366 1938 3370 1942
rect 3374 1938 3378 1942
rect 3390 1938 3394 1942
rect 3422 1938 3426 1942
rect 3534 1938 3538 1942
rect 3558 1938 3562 1942
rect 3582 1938 3586 1942
rect 3950 1947 3954 1951
rect 3982 1948 3986 1952
rect 4038 1948 4042 1952
rect 4086 1948 4090 1952
rect 4094 1948 4098 1952
rect 4102 1948 4106 1952
rect 4126 1948 4130 1952
rect 4158 1948 4162 1952
rect 4166 1948 4170 1952
rect 4190 1948 4194 1952
rect 4206 1948 4210 1952
rect 4222 1948 4226 1952
rect 4238 1958 4242 1962
rect 4438 1958 4442 1962
rect 4454 1958 4458 1962
rect 4286 1947 4290 1951
rect 4382 1948 4386 1952
rect 4414 1948 4418 1952
rect 4470 1948 4474 1952
rect 4494 1958 4498 1962
rect 4654 1958 4658 1962
rect 4598 1947 4602 1951
rect 4654 1948 4658 1952
rect 4678 1958 4682 1962
rect 4766 1958 4770 1962
rect 4822 1958 4826 1962
rect 4846 1958 4850 1962
rect 4702 1948 4706 1952
rect 4710 1948 4714 1952
rect 4734 1948 4738 1952
rect 4782 1948 4786 1952
rect 4870 1958 4874 1962
rect 5190 1958 5194 1962
rect 4870 1948 4874 1952
rect 4958 1948 4962 1952
rect 4998 1948 5002 1952
rect 5054 1948 5058 1952
rect 5078 1948 5082 1952
rect 5118 1948 5122 1952
rect 5150 1948 5154 1952
rect 3758 1938 3762 1942
rect 3830 1938 3834 1942
rect 3854 1938 3858 1942
rect 3918 1938 3922 1942
rect 4046 1938 4050 1942
rect 4198 1938 4202 1942
rect 4254 1938 4258 1942
rect 4270 1938 4274 1942
rect 4374 1938 4378 1942
rect 4406 1938 4410 1942
rect 4438 1938 4442 1942
rect 4462 1938 4466 1942
rect 4510 1938 4514 1942
rect 4566 1938 4570 1942
rect 4614 1938 4618 1942
rect 4638 1938 4642 1942
rect 4694 1938 4698 1942
rect 4750 1938 4754 1942
rect 4774 1938 4778 1942
rect 4806 1938 4810 1942
rect 4830 1938 4834 1942
rect 4934 1938 4938 1942
rect 4982 1938 4986 1942
rect 5126 1938 5130 1942
rect 5174 1938 5178 1942
rect 334 1928 338 1932
rect 406 1928 410 1932
rect 566 1928 570 1932
rect 1206 1928 1210 1932
rect 1414 1928 1418 1932
rect 1486 1928 1490 1932
rect 1918 1928 1922 1932
rect 2358 1928 2362 1932
rect 2390 1928 2394 1932
rect 2470 1928 2474 1932
rect 2870 1928 2874 1932
rect 2926 1928 2930 1932
rect 2958 1928 2962 1932
rect 3030 1928 3034 1932
rect 3550 1928 3554 1932
rect 3790 1928 3794 1932
rect 4070 1928 4074 1932
rect 4174 1928 4178 1932
rect 4358 1928 4362 1932
rect 4390 1928 4394 1932
rect 4422 1928 4426 1932
rect 5166 1928 5170 1932
rect 398 1918 402 1922
rect 438 1918 442 1922
rect 758 1918 762 1922
rect 766 1918 770 1922
rect 958 1918 962 1922
rect 974 1918 978 1922
rect 1038 1918 1042 1922
rect 1086 1918 1090 1922
rect 1278 1918 1282 1922
rect 1406 1918 1410 1922
rect 1614 1918 1618 1922
rect 2142 1918 2146 1922
rect 2214 1918 2218 1922
rect 2270 1918 2274 1922
rect 2542 1918 2546 1922
rect 2574 1918 2578 1922
rect 2614 1918 2618 1922
rect 2734 1918 2738 1922
rect 2990 1918 2994 1922
rect 3094 1918 3098 1922
rect 3198 1918 3202 1922
rect 3230 1918 3234 1922
rect 3350 1918 3354 1922
rect 3542 1918 3546 1922
rect 3646 1918 3650 1922
rect 3838 1918 3842 1922
rect 3878 1918 3882 1922
rect 4054 1918 4058 1922
rect 4366 1918 4370 1922
rect 4430 1918 4434 1922
rect 4766 1918 4770 1922
rect 5006 1918 5010 1922
rect 5134 1918 5138 1922
rect 1050 1903 1054 1907
rect 1057 1903 1061 1907
rect 2074 1903 2078 1907
rect 2081 1903 2085 1907
rect 3098 1903 3102 1907
rect 3105 1903 3109 1907
rect 4114 1903 4118 1907
rect 4121 1903 4125 1907
rect 6 1888 10 1892
rect 246 1888 250 1892
rect 366 1888 370 1892
rect 382 1888 386 1892
rect 414 1888 418 1892
rect 446 1888 450 1892
rect 486 1888 490 1892
rect 742 1888 746 1892
rect 782 1888 786 1892
rect 1190 1888 1194 1892
rect 1486 1888 1490 1892
rect 1550 1888 1554 1892
rect 1590 1888 1594 1892
rect 1830 1888 1834 1892
rect 1902 1888 1906 1892
rect 1974 1888 1978 1892
rect 2158 1888 2162 1892
rect 2206 1888 2210 1892
rect 2374 1888 2378 1892
rect 2430 1888 2434 1892
rect 2494 1888 2498 1892
rect 2782 1888 2786 1892
rect 2870 1888 2874 1892
rect 2910 1888 2914 1892
rect 3038 1888 3042 1892
rect 3438 1888 3442 1892
rect 3534 1888 3538 1892
rect 3574 1888 3578 1892
rect 3606 1888 3610 1892
rect 3862 1888 3866 1892
rect 3870 1888 3874 1892
rect 4318 1888 4322 1892
rect 4422 1888 4426 1892
rect 4542 1888 4546 1892
rect 4854 1888 4858 1892
rect 4966 1888 4970 1892
rect 5086 1888 5090 1892
rect 5190 1888 5194 1892
rect 166 1878 170 1882
rect 174 1878 178 1882
rect 374 1878 378 1882
rect 734 1878 738 1882
rect 870 1878 874 1882
rect 1430 1878 1434 1882
rect 1446 1878 1450 1882
rect 1598 1878 1602 1882
rect 2030 1878 2034 1882
rect 2902 1878 2906 1882
rect 3006 1878 3010 1882
rect 3542 1878 3546 1882
rect 3670 1878 3674 1882
rect 3998 1878 4002 1882
rect 4062 1878 4066 1882
rect 4310 1878 4314 1882
rect 4614 1878 4618 1882
rect 4798 1878 4802 1882
rect 4974 1878 4978 1882
rect 5166 1878 5170 1882
rect 62 1868 66 1872
rect 102 1868 106 1872
rect 126 1868 130 1872
rect 158 1868 162 1872
rect 190 1868 194 1872
rect 214 1868 218 1872
rect 270 1868 274 1872
rect 302 1868 306 1872
rect 334 1868 338 1872
rect 390 1868 394 1872
rect 438 1868 442 1872
rect 462 1868 466 1872
rect 502 1868 506 1872
rect 590 1868 594 1872
rect 70 1859 74 1863
rect 118 1858 122 1862
rect 142 1858 146 1862
rect 150 1858 154 1862
rect 206 1858 210 1862
rect 222 1858 226 1862
rect 262 1858 266 1862
rect 310 1858 314 1862
rect 398 1858 402 1862
rect 470 1858 474 1862
rect 574 1858 578 1862
rect 638 1858 642 1862
rect 670 1859 674 1863
rect 750 1868 754 1872
rect 806 1868 810 1872
rect 814 1868 818 1872
rect 838 1868 842 1872
rect 1014 1868 1018 1872
rect 1022 1868 1026 1872
rect 1094 1868 1098 1872
rect 1198 1868 1202 1872
rect 1230 1868 1234 1872
rect 1262 1868 1266 1872
rect 1326 1868 1330 1872
rect 1342 1868 1346 1872
rect 1366 1868 1370 1872
rect 1494 1868 1498 1872
rect 1734 1868 1738 1872
rect 1766 1868 1770 1872
rect 1806 1868 1810 1872
rect 1822 1868 1826 1872
rect 1846 1868 1850 1872
rect 2182 1868 2186 1872
rect 2230 1868 2234 1872
rect 2398 1868 2402 1872
rect 2406 1868 2410 1872
rect 2438 1868 2442 1872
rect 2590 1868 2594 1872
rect 2622 1868 2626 1872
rect 2686 1868 2690 1872
rect 2702 1868 2706 1872
rect 2806 1868 2810 1872
rect 2814 1868 2818 1872
rect 2862 1868 2866 1872
rect 3022 1868 3026 1872
rect 3078 1868 3082 1872
rect 3110 1868 3114 1872
rect 3142 1868 3146 1872
rect 3166 1868 3170 1872
rect 3182 1868 3186 1872
rect 3230 1868 3234 1872
rect 3358 1868 3362 1872
rect 3582 1868 3586 1872
rect 3614 1868 3618 1872
rect 3638 1868 3642 1872
rect 3846 1868 3850 1872
rect 3982 1868 3986 1872
rect 4086 1868 4090 1872
rect 4102 1868 4106 1872
rect 4158 1868 4162 1872
rect 4174 1868 4178 1872
rect 4294 1868 4298 1872
rect 4342 1868 4346 1872
rect 4430 1868 4434 1872
rect 4446 1868 4450 1872
rect 4478 1868 4482 1872
rect 4534 1868 4538 1872
rect 4582 1868 4586 1872
rect 4590 1868 4594 1872
rect 4726 1868 4730 1872
rect 4742 1868 4746 1872
rect 4774 1868 4778 1872
rect 4838 1868 4842 1872
rect 4934 1868 4938 1872
rect 4958 1868 4962 1872
rect 4990 1868 4994 1872
rect 5102 1868 5106 1872
rect 702 1858 706 1862
rect 710 1858 714 1862
rect 726 1858 730 1862
rect 750 1858 754 1862
rect 798 1858 802 1862
rect 830 1858 834 1862
rect 878 1858 882 1862
rect 966 1858 970 1862
rect 982 1858 986 1862
rect 1006 1858 1010 1862
rect 1030 1858 1034 1862
rect 1078 1858 1082 1862
rect 1086 1858 1090 1862
rect 1126 1859 1130 1863
rect 1150 1858 1154 1862
rect 1206 1858 1210 1862
rect 1222 1858 1226 1862
rect 1238 1858 1242 1862
rect 1358 1859 1362 1863
rect 1470 1858 1474 1862
rect 1502 1858 1506 1862
rect 1518 1858 1522 1862
rect 1526 1858 1530 1862
rect 1534 1858 1538 1862
rect 1558 1858 1562 1862
rect 1638 1858 1642 1862
rect 1662 1858 1666 1862
rect 1726 1858 1730 1862
rect 1774 1858 1778 1862
rect 1782 1858 1786 1862
rect 1806 1858 1810 1862
rect 1854 1858 1858 1862
rect 1910 1858 1914 1862
rect 1918 1858 1922 1862
rect 1950 1858 1954 1862
rect 1958 1858 1962 1862
rect 2014 1858 2018 1862
rect 2054 1858 2058 1862
rect 2102 1858 2106 1862
rect 2134 1858 2138 1862
rect 2142 1858 2146 1862
rect 2166 1858 2170 1862
rect 2190 1858 2194 1862
rect 2270 1858 2274 1862
rect 2294 1858 2298 1862
rect 2350 1858 2354 1862
rect 2358 1858 2362 1862
rect 2414 1858 2418 1862
rect 2486 1858 2490 1862
rect 2566 1858 2570 1862
rect 2726 1858 2730 1862
rect 2854 1858 2858 1862
rect 2886 1858 2890 1862
rect 2950 1858 2954 1862
rect 2974 1859 2978 1863
rect 3022 1858 3026 1862
rect 3062 1858 3066 1862
rect 3134 1858 3138 1862
rect 3158 1858 3162 1862
rect 3238 1858 3242 1862
rect 3318 1858 3322 1862
rect 3326 1858 3330 1862
rect 3334 1858 3338 1862
rect 3382 1858 3386 1862
rect 3478 1858 3482 1862
rect 3502 1858 3506 1862
rect 3558 1858 3562 1862
rect 3590 1858 3594 1862
rect 3638 1858 3642 1862
rect 3662 1858 3666 1862
rect 3718 1858 3722 1862
rect 3742 1858 3746 1862
rect 3806 1858 3810 1862
rect 3814 1858 3818 1862
rect 3902 1858 3906 1862
rect 3934 1859 3938 1863
rect 4022 1858 4026 1862
rect 4086 1858 4090 1862
rect 4166 1858 4170 1862
rect 4206 1858 4210 1862
rect 4278 1859 4282 1863
rect 4326 1858 4330 1862
rect 4366 1858 4370 1862
rect 4382 1858 4386 1862
rect 4430 1858 4434 1862
rect 4486 1858 4490 1862
rect 4494 1858 4498 1862
rect 4518 1858 4522 1862
rect 4574 1858 4578 1862
rect 4710 1859 4714 1863
rect 4750 1858 4754 1862
rect 4814 1858 4818 1862
rect 4846 1858 4850 1862
rect 4910 1858 4914 1862
rect 4950 1858 4954 1862
rect 5014 1858 5018 1862
rect 5134 1858 5138 1862
rect 102 1848 106 1852
rect 134 1848 138 1852
rect 238 1848 242 1852
rect 422 1848 426 1852
rect 446 1848 450 1852
rect 726 1848 730 1852
rect 774 1848 778 1852
rect 782 1848 786 1852
rect 982 1848 986 1852
rect 990 1848 994 1852
rect 1062 1848 1066 1852
rect 1222 1848 1226 1852
rect 1238 1848 1242 1852
rect 1486 1848 1490 1852
rect 1518 1848 1522 1852
rect 1750 1848 1754 1852
rect 1870 1848 1874 1852
rect 2214 1848 2218 1852
rect 2382 1848 2386 1852
rect 2430 1848 2434 1852
rect 2454 1848 2458 1852
rect 2478 1848 2482 1852
rect 3078 1848 3082 1852
rect 3094 1848 3098 1852
rect 3342 1848 3346 1852
rect 3598 1848 3602 1852
rect 3662 1848 3666 1852
rect 3862 1848 3866 1852
rect 3966 1848 3970 1852
rect 4102 1848 4106 1852
rect 4150 1848 4154 1852
rect 4462 1848 4466 1852
rect 4550 1848 4554 1852
rect 4558 1848 4562 1852
rect 4606 1848 4610 1852
rect 4766 1848 4770 1852
rect 4790 1848 4794 1852
rect 814 1838 818 1842
rect 942 1838 946 1842
rect 1254 1838 1258 1842
rect 1422 1838 1426 1842
rect 1838 1838 1842 1842
rect 1934 1838 1938 1842
rect 2118 1838 2122 1842
rect 2310 1838 2314 1842
rect 3038 1838 3042 1842
rect 3054 1838 3058 1842
rect 3198 1838 3202 1842
rect 4110 1838 4114 1842
rect 4142 1838 4146 1842
rect 4214 1838 4218 1842
rect 4574 1838 4578 1842
rect 4750 1838 4754 1842
rect 4822 1838 4826 1842
rect 5054 1838 5058 1842
rect 1438 1828 1442 1832
rect 758 1818 762 1822
rect 1006 1818 1010 1822
rect 1710 1818 1714 1822
rect 1974 1818 1978 1822
rect 1998 1818 2002 1822
rect 2062 1818 2066 1822
rect 2798 1818 2802 1822
rect 2838 1818 2842 1822
rect 3062 1818 3066 1822
rect 3790 1818 3794 1822
rect 3830 1818 3834 1822
rect 3974 1818 3978 1822
rect 4038 1818 4042 1822
rect 4094 1818 4098 1822
rect 4190 1818 4194 1822
rect 4502 1818 4506 1822
rect 4598 1818 4602 1822
rect 4782 1818 4786 1822
rect 538 1803 542 1807
rect 545 1803 549 1807
rect 1562 1803 1566 1807
rect 1569 1803 1573 1807
rect 2586 1803 2590 1807
rect 2593 1803 2597 1807
rect 3610 1803 3614 1807
rect 3617 1803 3621 1807
rect 4634 1803 4638 1807
rect 4641 1803 4645 1807
rect 62 1788 66 1792
rect 166 1788 170 1792
rect 838 1788 842 1792
rect 918 1788 922 1792
rect 1174 1788 1178 1792
rect 1222 1788 1226 1792
rect 1934 1788 1938 1792
rect 2246 1788 2250 1792
rect 2446 1788 2450 1792
rect 2742 1788 2746 1792
rect 2934 1788 2938 1792
rect 3150 1788 3154 1792
rect 3190 1788 3194 1792
rect 3278 1788 3282 1792
rect 3486 1788 3490 1792
rect 3550 1788 3554 1792
rect 3582 1788 3586 1792
rect 3870 1788 3874 1792
rect 3974 1788 3978 1792
rect 4078 1788 4082 1792
rect 4214 1788 4218 1792
rect 4278 1788 4282 1792
rect 4318 1788 4322 1792
rect 4366 1788 4370 1792
rect 5102 1788 5106 1792
rect 5182 1788 5186 1792
rect 318 1778 322 1782
rect 1966 1778 1970 1782
rect 3414 1778 3418 1782
rect 3654 1778 3658 1782
rect 4638 1778 4642 1782
rect 4926 1778 4930 1782
rect 302 1768 306 1772
rect 358 1768 362 1772
rect 478 1768 482 1772
rect 710 1768 714 1772
rect 1318 1768 1322 1772
rect 3054 1768 3058 1772
rect 3782 1768 3786 1772
rect 4438 1768 4442 1772
rect 4478 1768 4482 1772
rect 4774 1768 4778 1772
rect 334 1758 338 1762
rect 102 1747 106 1751
rect 198 1748 202 1752
rect 6 1738 10 1742
rect 70 1738 74 1742
rect 86 1738 90 1742
rect 190 1738 194 1742
rect 262 1748 266 1752
rect 326 1748 330 1752
rect 542 1758 546 1762
rect 694 1758 698 1762
rect 742 1758 746 1762
rect 886 1758 890 1762
rect 966 1758 970 1762
rect 1086 1758 1090 1762
rect 1422 1758 1426 1762
rect 1742 1758 1746 1762
rect 1766 1758 1770 1762
rect 374 1748 378 1752
rect 430 1748 434 1752
rect 486 1748 490 1752
rect 502 1748 506 1752
rect 518 1748 522 1752
rect 622 1748 626 1752
rect 686 1748 690 1752
rect 726 1748 730 1752
rect 742 1748 746 1752
rect 326 1738 330 1742
rect 382 1738 386 1742
rect 398 1738 402 1742
rect 494 1738 498 1742
rect 574 1738 578 1742
rect 614 1738 618 1742
rect 710 1738 714 1742
rect 718 1738 722 1742
rect 774 1747 778 1751
rect 870 1748 874 1752
rect 878 1748 882 1752
rect 894 1748 898 1752
rect 902 1748 906 1752
rect 926 1748 930 1752
rect 950 1748 954 1752
rect 958 1748 962 1752
rect 998 1747 1002 1751
rect 1070 1748 1074 1752
rect 1102 1748 1106 1752
rect 1118 1748 1122 1752
rect 1158 1748 1162 1752
rect 1182 1748 1186 1752
rect 1198 1748 1202 1752
rect 1206 1748 1210 1752
rect 1230 1748 1234 1752
rect 1238 1748 1242 1752
rect 1246 1748 1250 1752
rect 1294 1748 1298 1752
rect 1334 1748 1338 1752
rect 1358 1748 1362 1752
rect 1398 1748 1402 1752
rect 1430 1748 1434 1752
rect 1526 1748 1530 1752
rect 1550 1748 1554 1752
rect 1654 1748 1658 1752
rect 1686 1747 1690 1751
rect 1718 1748 1722 1752
rect 1726 1748 1730 1752
rect 1734 1748 1738 1752
rect 2206 1758 2210 1762
rect 2374 1758 2378 1762
rect 2398 1758 2402 1762
rect 2414 1758 2418 1762
rect 1782 1748 1786 1752
rect 1790 1748 1794 1752
rect 1862 1748 1866 1752
rect 1918 1748 1922 1752
rect 1926 1748 1930 1752
rect 1958 1748 1962 1752
rect 2022 1748 2026 1752
rect 2102 1748 2106 1752
rect 2134 1748 2138 1752
rect 2142 1748 2146 1752
rect 2222 1748 2226 1752
rect 2238 1748 2242 1752
rect 2262 1748 2266 1752
rect 2310 1748 2314 1752
rect 2318 1748 2322 1752
rect 2414 1748 2418 1752
rect 2430 1748 2434 1752
rect 2438 1748 2442 1752
rect 2462 1748 2466 1752
rect 2470 1748 2474 1752
rect 2534 1758 2538 1762
rect 2566 1758 2570 1762
rect 2718 1758 2722 1762
rect 2782 1758 2786 1762
rect 2798 1758 2802 1762
rect 2902 1758 2906 1762
rect 2918 1758 2922 1762
rect 2974 1758 2978 1762
rect 3038 1758 3042 1762
rect 3430 1758 3434 1762
rect 3446 1758 3450 1762
rect 3526 1758 3530 1762
rect 3566 1758 3570 1762
rect 3646 1758 3650 1762
rect 2494 1748 2498 1752
rect 2518 1748 2522 1752
rect 2550 1748 2554 1752
rect 2558 1748 2562 1752
rect 2574 1748 2578 1752
rect 2662 1748 2666 1752
rect 2726 1748 2730 1752
rect 2734 1748 2738 1752
rect 2774 1748 2778 1752
rect 2782 1748 2786 1752
rect 2854 1748 2858 1752
rect 2934 1748 2938 1752
rect 2958 1748 2962 1752
rect 2982 1748 2986 1752
rect 3014 1748 3018 1752
rect 3054 1748 3058 1752
rect 3070 1748 3074 1752
rect 3078 1748 3082 1752
rect 3102 1748 3106 1752
rect 3174 1748 3178 1752
rect 3206 1748 3210 1752
rect 3214 1748 3218 1752
rect 3238 1748 3242 1752
rect 3270 1748 3274 1752
rect 3310 1748 3314 1752
rect 942 1738 946 1742
rect 982 1738 986 1742
rect 1030 1738 1034 1742
rect 1110 1738 1114 1742
rect 1254 1738 1258 1742
rect 1270 1738 1274 1742
rect 1406 1738 1410 1742
rect 1470 1738 1474 1742
rect 1486 1738 1490 1742
rect 1574 1738 1578 1742
rect 1606 1738 1610 1742
rect 1750 1738 1754 1742
rect 1798 1738 1802 1742
rect 1878 1738 1882 1742
rect 2046 1738 2050 1742
rect 2158 1738 2162 1742
rect 3342 1747 3346 1751
rect 3398 1748 3402 1752
rect 3422 1748 3426 1752
rect 3446 1748 3450 1752
rect 3462 1748 3466 1752
rect 3470 1748 3474 1752
rect 3494 1748 3498 1752
rect 3534 1748 3538 1752
rect 3590 1748 3594 1752
rect 3686 1748 3690 1752
rect 3710 1748 3714 1752
rect 3758 1748 3762 1752
rect 3766 1748 3770 1752
rect 4222 1758 4226 1762
rect 4294 1758 4298 1762
rect 3798 1748 3802 1752
rect 3814 1748 3818 1752
rect 3918 1748 3922 1752
rect 3982 1748 3986 1752
rect 4030 1748 4034 1752
rect 4038 1748 4042 1752
rect 4062 1748 4066 1752
rect 4142 1748 4146 1752
rect 4222 1748 4226 1752
rect 4238 1748 4242 1752
rect 4270 1748 4274 1752
rect 4302 1748 4306 1752
rect 4310 1748 4314 1752
rect 4334 1748 4338 1752
rect 4350 1748 4354 1752
rect 4382 1748 4386 1752
rect 4422 1748 4426 1752
rect 4462 1758 4466 1762
rect 4590 1758 4594 1762
rect 4462 1748 4466 1752
rect 4534 1748 4538 1752
rect 4758 1758 4762 1762
rect 4790 1758 4794 1762
rect 4806 1758 4810 1762
rect 4934 1758 4938 1762
rect 5078 1758 5082 1762
rect 4614 1748 4618 1752
rect 4718 1748 4722 1752
rect 4790 1748 4794 1752
rect 4806 1748 4810 1752
rect 4862 1747 4866 1751
rect 4934 1748 4938 1752
rect 4950 1748 4954 1752
rect 5022 1748 5026 1752
rect 5102 1748 5106 1752
rect 5134 1748 5138 1752
rect 5166 1748 5170 1752
rect 5190 1748 5194 1752
rect 2222 1738 2226 1742
rect 2390 1738 2394 1742
rect 2422 1738 2426 1742
rect 2478 1738 2482 1742
rect 2502 1738 2506 1742
rect 2510 1738 2514 1742
rect 2542 1738 2546 1742
rect 2702 1738 2706 1742
rect 2774 1738 2778 1742
rect 2838 1738 2842 1742
rect 2942 1738 2946 1742
rect 2966 1738 2970 1742
rect 2982 1738 2986 1742
rect 3062 1738 3066 1742
rect 3134 1738 3138 1742
rect 3246 1738 3250 1742
rect 3262 1738 3266 1742
rect 3358 1738 3362 1742
rect 3374 1738 3378 1742
rect 3390 1738 3394 1742
rect 3454 1738 3458 1742
rect 3510 1738 3514 1742
rect 3630 1738 3634 1742
rect 3718 1738 3722 1742
rect 3750 1738 3754 1742
rect 3806 1738 3810 1742
rect 3838 1738 3842 1742
rect 3910 1738 3914 1742
rect 3990 1738 3994 1742
rect 4054 1738 4058 1742
rect 4118 1738 4122 1742
rect 4246 1738 4250 1742
rect 4406 1738 4410 1742
rect 4414 1738 4418 1742
rect 4470 1738 4474 1742
rect 4558 1738 4562 1742
rect 4574 1738 4578 1742
rect 4606 1738 4610 1742
rect 4726 1738 4730 1742
rect 4782 1738 4786 1742
rect 4814 1738 4818 1742
rect 4846 1738 4850 1742
rect 4958 1738 4962 1742
rect 5014 1738 5018 1742
rect 5062 1738 5066 1742
rect 5118 1738 5122 1742
rect 5158 1738 5162 1742
rect 174 1728 178 1732
rect 206 1728 210 1732
rect 222 1728 226 1732
rect 254 1728 258 1732
rect 542 1728 546 1732
rect 686 1728 690 1732
rect 774 1728 778 1732
rect 1270 1728 1274 1732
rect 1294 1728 1298 1732
rect 1446 1728 1450 1732
rect 1454 1728 1458 1732
rect 2086 1728 2090 1732
rect 2118 1728 2122 1732
rect 2670 1728 2674 1732
rect 3030 1728 3034 1732
rect 3126 1728 3130 1732
rect 3166 1728 3170 1732
rect 3222 1728 3226 1732
rect 3374 1728 3378 1732
rect 3406 1728 3410 1732
rect 3606 1728 3610 1732
rect 3830 1728 3834 1732
rect 4014 1728 4018 1732
rect 4030 1728 4034 1732
rect 4254 1728 4258 1732
rect 4830 1728 4834 1732
rect 5118 1728 5122 1732
rect 5174 1728 5178 1732
rect 166 1718 170 1722
rect 182 1718 186 1722
rect 566 1718 570 1722
rect 670 1718 674 1722
rect 1070 1718 1074 1722
rect 1134 1718 1138 1722
rect 1262 1718 1266 1722
rect 1302 1718 1306 1722
rect 1462 1718 1466 1722
rect 1486 1718 1490 1722
rect 2190 1718 2194 1722
rect 2206 1718 2210 1722
rect 2278 1718 2282 1722
rect 2374 1718 2378 1722
rect 2534 1718 2538 1722
rect 2718 1718 2722 1722
rect 2998 1718 3002 1722
rect 3526 1718 3530 1722
rect 3646 1718 3650 1722
rect 3998 1718 4002 1722
rect 4214 1718 4218 1722
rect 4822 1718 4826 1722
rect 4966 1718 4970 1722
rect 5150 1718 5154 1722
rect 1050 1703 1054 1707
rect 1057 1703 1061 1707
rect 2074 1703 2078 1707
rect 2081 1703 2085 1707
rect 3098 1703 3102 1707
rect 3105 1703 3109 1707
rect 4114 1703 4118 1707
rect 4121 1703 4125 1707
rect 94 1688 98 1692
rect 222 1688 226 1692
rect 574 1688 578 1692
rect 702 1688 706 1692
rect 750 1688 754 1692
rect 766 1688 770 1692
rect 926 1688 930 1692
rect 958 1688 962 1692
rect 966 1688 970 1692
rect 990 1688 994 1692
rect 1030 1688 1034 1692
rect 1222 1688 1226 1692
rect 1270 1688 1274 1692
rect 1318 1688 1322 1692
rect 1430 1688 1434 1692
rect 1526 1688 1530 1692
rect 1830 1688 1834 1692
rect 1918 1688 1922 1692
rect 1950 1688 1954 1692
rect 2014 1688 2018 1692
rect 2158 1688 2162 1692
rect 2214 1688 2218 1692
rect 2398 1688 2402 1692
rect 2422 1688 2426 1692
rect 2430 1688 2434 1692
rect 2462 1688 2466 1692
rect 2470 1688 2474 1692
rect 2726 1688 2730 1692
rect 2774 1688 2778 1692
rect 2838 1688 2842 1692
rect 2862 1688 2866 1692
rect 3038 1688 3042 1692
rect 3182 1688 3186 1692
rect 3190 1688 3194 1692
rect 3398 1688 3402 1692
rect 3454 1688 3458 1692
rect 3462 1688 3466 1692
rect 3478 1688 3482 1692
rect 3686 1688 3690 1692
rect 3982 1688 3986 1692
rect 4014 1688 4018 1692
rect 4070 1688 4074 1692
rect 4102 1688 4106 1692
rect 4390 1688 4394 1692
rect 4470 1688 4474 1692
rect 4526 1688 4530 1692
rect 4566 1688 4570 1692
rect 4606 1688 4610 1692
rect 4686 1688 4690 1692
rect 4894 1688 4898 1692
rect 4910 1688 4914 1692
rect 4958 1688 4962 1692
rect 5078 1688 5082 1692
rect 126 1678 130 1682
rect 158 1678 162 1682
rect 254 1678 258 1682
rect 366 1678 370 1682
rect 502 1678 506 1682
rect 510 1678 514 1682
rect 518 1678 522 1682
rect 830 1678 834 1682
rect 1062 1678 1066 1682
rect 1102 1678 1106 1682
rect 1174 1678 1178 1682
rect 1302 1678 1306 1682
rect 1366 1678 1370 1682
rect 1902 1678 1906 1682
rect 6 1668 10 1672
rect 86 1668 90 1672
rect 326 1668 330 1672
rect 438 1668 442 1672
rect 494 1668 498 1672
rect 582 1668 586 1672
rect 622 1668 626 1672
rect 638 1668 642 1672
rect 646 1668 650 1672
rect 726 1668 730 1672
rect 782 1668 786 1672
rect 790 1668 794 1672
rect 806 1668 810 1672
rect 830 1668 834 1672
rect 894 1668 898 1672
rect 934 1668 938 1672
rect 982 1668 986 1672
rect 1014 1668 1018 1672
rect 1038 1668 1042 1672
rect 1054 1668 1058 1672
rect 1190 1668 1194 1672
rect 1230 1668 1234 1672
rect 1262 1668 1266 1672
rect 1462 1668 1466 1672
rect 1574 1668 1578 1672
rect 1678 1668 1682 1672
rect 1702 1668 1706 1672
rect 1726 1668 1730 1672
rect 1806 1668 1810 1672
rect 1862 1668 1866 1672
rect 2198 1678 2202 1682
rect 1926 1668 1930 1672
rect 1998 1668 2002 1672
rect 2086 1668 2090 1672
rect 2134 1668 2138 1672
rect 2174 1668 2178 1672
rect 2238 1678 2242 1682
rect 2438 1678 2442 1682
rect 2766 1678 2770 1682
rect 3158 1678 3162 1682
rect 3414 1678 3418 1682
rect 3470 1678 3474 1682
rect 3726 1678 3730 1682
rect 4646 1678 4650 1682
rect 4918 1678 4922 1682
rect 4974 1678 4978 1682
rect 2222 1668 2226 1672
rect 2310 1668 2314 1672
rect 2350 1668 2354 1672
rect 2382 1668 2386 1672
rect 2406 1668 2410 1672
rect 2446 1668 2450 1672
rect 2550 1668 2554 1672
rect 2614 1668 2618 1672
rect 2670 1668 2674 1672
rect 2734 1668 2738 1672
rect 2782 1668 2786 1672
rect 2870 1668 2874 1672
rect 2958 1668 2962 1672
rect 2974 1668 2978 1672
rect 3022 1668 3026 1672
rect 3046 1668 3050 1672
rect 3054 1668 3058 1672
rect 3118 1668 3122 1672
rect 3166 1668 3170 1672
rect 3310 1668 3314 1672
rect 3318 1668 3322 1672
rect 3390 1668 3394 1672
rect 3406 1668 3410 1672
rect 3574 1668 3578 1672
rect 3646 1668 3650 1672
rect 3758 1668 3762 1672
rect 3814 1668 3818 1672
rect 3870 1668 3874 1672
rect 3910 1668 3914 1672
rect 3990 1668 3994 1672
rect 4022 1668 4026 1672
rect 4062 1668 4066 1672
rect 4214 1668 4218 1672
rect 4222 1668 4226 1672
rect 4278 1668 4282 1672
rect 4286 1668 4290 1672
rect 4366 1668 4370 1672
rect 4398 1668 4402 1672
rect 4550 1668 4554 1672
rect 4598 1668 4602 1672
rect 4630 1668 4634 1672
rect 4678 1668 4682 1672
rect 4710 1668 4714 1672
rect 4718 1668 4722 1672
rect 4870 1668 4874 1672
rect 4886 1668 4890 1672
rect 4950 1668 4954 1672
rect 5014 1668 5018 1672
rect 5054 1668 5058 1672
rect 5158 1668 5162 1672
rect 78 1658 82 1662
rect 110 1658 114 1662
rect 182 1658 186 1662
rect 262 1658 266 1662
rect 374 1658 378 1662
rect 446 1658 450 1662
rect 486 1658 490 1662
rect 558 1658 562 1662
rect 590 1658 594 1662
rect 606 1658 610 1662
rect 646 1658 650 1662
rect 654 1658 658 1662
rect 662 1658 666 1662
rect 678 1658 682 1662
rect 686 1658 690 1662
rect 710 1658 714 1662
rect 734 1658 738 1662
rect 782 1658 786 1662
rect 814 1658 818 1662
rect 862 1659 866 1663
rect 942 1658 946 1662
rect 1014 1658 1018 1662
rect 1110 1658 1114 1662
rect 1190 1658 1194 1662
rect 1206 1658 1210 1662
rect 1254 1658 1258 1662
rect 1286 1658 1290 1662
rect 1334 1658 1338 1662
rect 1374 1658 1378 1662
rect 1438 1658 1442 1662
rect 1454 1658 1458 1662
rect 1478 1658 1482 1662
rect 1494 1658 1498 1662
rect 1510 1658 1514 1662
rect 1534 1658 1538 1662
rect 1542 1658 1546 1662
rect 1598 1658 1602 1662
rect 1670 1658 1674 1662
rect 1718 1658 1722 1662
rect 1742 1658 1746 1662
rect 1750 1658 1754 1662
rect 1758 1658 1762 1662
rect 1774 1658 1778 1662
rect 1798 1658 1802 1662
rect 1814 1658 1818 1662
rect 1822 1658 1826 1662
rect 1846 1658 1850 1662
rect 1886 1658 1890 1662
rect 1934 1658 1938 1662
rect 1974 1658 1978 1662
rect 2030 1658 2034 1662
rect 2038 1658 2042 1662
rect 2046 1658 2050 1662
rect 2070 1658 2074 1662
rect 2078 1658 2082 1662
rect 2126 1658 2130 1662
rect 2174 1658 2178 1662
rect 2230 1658 2234 1662
rect 2318 1659 2322 1663
rect 2350 1658 2354 1662
rect 2534 1659 2538 1663
rect 2566 1658 2570 1662
rect 2678 1658 2682 1662
rect 2694 1658 2698 1662
rect 2750 1658 2754 1662
rect 2942 1659 2946 1663
rect 3014 1658 3018 1662
rect 3118 1658 3122 1662
rect 3166 1658 3170 1662
rect 3222 1658 3226 1662
rect 3246 1658 3250 1662
rect 3302 1658 3306 1662
rect 3438 1658 3442 1662
rect 3510 1658 3514 1662
rect 3542 1659 3546 1663
rect 3574 1658 3578 1662
rect 3638 1658 3642 1662
rect 3654 1658 3658 1662
rect 3702 1658 3706 1662
rect 3734 1658 3738 1662
rect 3750 1658 3754 1662
rect 3774 1658 3778 1662
rect 3798 1658 3802 1662
rect 3806 1658 3810 1662
rect 3822 1658 3826 1662
rect 3854 1658 3858 1662
rect 3862 1658 3866 1662
rect 3902 1659 3906 1663
rect 3998 1658 4002 1662
rect 4046 1658 4050 1662
rect 4086 1658 4090 1662
rect 4118 1658 4122 1662
rect 4142 1658 4146 1662
rect 4150 1658 4154 1662
rect 4206 1658 4210 1662
rect 4230 1658 4234 1662
rect 4286 1658 4290 1662
rect 4294 1658 4298 1662
rect 4302 1658 4306 1662
rect 4318 1658 4322 1662
rect 4350 1658 4354 1662
rect 4414 1658 4418 1662
rect 4438 1658 4442 1662
rect 4446 1658 4450 1662
rect 4454 1658 4458 1662
rect 4462 1658 4466 1662
rect 4486 1658 4490 1662
rect 4502 1658 4506 1662
rect 4510 1658 4514 1662
rect 4534 1658 4538 1662
rect 4574 1658 4578 1662
rect 4590 1658 4594 1662
rect 4646 1658 4650 1662
rect 4654 1658 4658 1662
rect 4670 1658 4674 1662
rect 4702 1658 4706 1662
rect 4758 1658 4762 1662
rect 4766 1658 4770 1662
rect 4846 1658 4850 1662
rect 4942 1658 4946 1662
rect 5022 1659 5026 1663
rect 5150 1658 5154 1662
rect 446 1648 450 1652
rect 470 1648 474 1652
rect 574 1648 578 1652
rect 606 1648 610 1652
rect 614 1648 618 1652
rect 670 1648 674 1652
rect 750 1648 754 1652
rect 758 1648 762 1652
rect 958 1648 962 1652
rect 966 1648 970 1652
rect 990 1648 994 1652
rect 1022 1648 1026 1652
rect 1182 1648 1186 1652
rect 1246 1648 1250 1652
rect 1438 1648 1442 1652
rect 1494 1648 1498 1652
rect 1694 1648 1698 1652
rect 1758 1648 1762 1652
rect 1878 1648 1882 1652
rect 2150 1648 2154 1652
rect 2158 1648 2162 1652
rect 2374 1648 2378 1652
rect 2398 1648 2402 1652
rect 2422 1648 2426 1652
rect 2462 1648 2466 1652
rect 2630 1648 2634 1652
rect 2734 1648 2738 1652
rect 2990 1648 2994 1652
rect 3030 1648 3034 1652
rect 3286 1648 3290 1652
rect 3390 1648 3394 1652
rect 3454 1648 3458 1652
rect 3582 1648 3586 1652
rect 3606 1648 3610 1652
rect 3670 1648 3674 1652
rect 3686 1648 3690 1652
rect 4030 1648 4034 1652
rect 4190 1648 4194 1652
rect 4246 1648 4250 1652
rect 4566 1648 4570 1652
rect 4574 1648 4578 1652
rect 4606 1648 4610 1652
rect 4686 1648 4690 1652
rect 4734 1648 4738 1652
rect 4758 1648 4762 1652
rect 4902 1648 4906 1652
rect 4926 1648 4930 1652
rect 5070 1648 5074 1652
rect 430 1638 434 1642
rect 1150 1638 1154 1642
rect 1166 1638 1170 1642
rect 2358 1638 2362 1642
rect 2854 1638 2858 1642
rect 2878 1638 2882 1642
rect 3302 1638 3306 1642
rect 3726 1638 3730 1642
rect 3838 1638 3842 1642
rect 3966 1638 3970 1642
rect 4158 1638 4162 1642
rect 4310 1638 4314 1642
rect 4654 1638 4658 1642
rect 4942 1638 4946 1642
rect 4422 1628 4426 1632
rect 62 1618 66 1622
rect 318 1618 322 1622
rect 1318 1618 1322 1622
rect 1870 1618 1874 1622
rect 1950 1618 1954 1622
rect 2014 1618 2018 1622
rect 2118 1618 2122 1622
rect 2142 1618 2146 1622
rect 2582 1618 2586 1622
rect 2622 1618 2626 1622
rect 2838 1618 2842 1622
rect 3014 1618 3018 1622
rect 3790 1618 3794 1622
rect 4070 1618 4074 1622
rect 4270 1618 4274 1622
rect 4390 1618 4394 1622
rect 5062 1618 5066 1622
rect 538 1603 542 1607
rect 545 1603 549 1607
rect 1562 1603 1566 1607
rect 1569 1603 1573 1607
rect 2586 1603 2590 1607
rect 2593 1603 2597 1607
rect 3610 1603 3614 1607
rect 3617 1603 3621 1607
rect 4634 1603 4638 1607
rect 4641 1603 4645 1607
rect 246 1588 250 1592
rect 286 1588 290 1592
rect 366 1588 370 1592
rect 598 1588 602 1592
rect 622 1588 626 1592
rect 646 1588 650 1592
rect 662 1588 666 1592
rect 934 1588 938 1592
rect 1006 1588 1010 1592
rect 1046 1588 1050 1592
rect 1102 1588 1106 1592
rect 1174 1588 1178 1592
rect 1326 1588 1330 1592
rect 1462 1588 1466 1592
rect 1614 1588 1618 1592
rect 1726 1588 1730 1592
rect 1774 1588 1778 1592
rect 1854 1588 1858 1592
rect 1918 1588 1922 1592
rect 2022 1588 2026 1592
rect 2070 1588 2074 1592
rect 2182 1588 2186 1592
rect 2318 1588 2322 1592
rect 2406 1588 2410 1592
rect 2942 1588 2946 1592
rect 2990 1588 2994 1592
rect 3110 1588 3114 1592
rect 3206 1588 3210 1592
rect 3310 1588 3314 1592
rect 3414 1588 3418 1592
rect 3726 1588 3730 1592
rect 3838 1588 3842 1592
rect 3910 1588 3914 1592
rect 4022 1588 4026 1592
rect 4110 1588 4114 1592
rect 4182 1588 4186 1592
rect 4374 1588 4378 1592
rect 4838 1588 4842 1592
rect 4878 1588 4882 1592
rect 766 1578 770 1582
rect 1310 1578 1314 1582
rect 1430 1578 1434 1582
rect 2286 1578 2290 1582
rect 2918 1578 2922 1582
rect 3158 1578 3162 1582
rect 3334 1578 3338 1582
rect 3574 1578 3578 1582
rect 3870 1578 3874 1582
rect 94 1568 98 1572
rect 310 1568 314 1572
rect 550 1568 554 1572
rect 774 1568 778 1572
rect 1214 1568 1218 1572
rect 1334 1568 1338 1572
rect 3382 1568 3386 1572
rect 3430 1568 3434 1572
rect 4406 1568 4410 1572
rect 4894 1568 4898 1572
rect 38 1548 42 1552
rect 62 1548 66 1552
rect 102 1548 106 1552
rect 118 1548 122 1552
rect 134 1548 138 1552
rect 182 1547 186 1551
rect 270 1548 274 1552
rect 278 1548 282 1552
rect 382 1558 386 1562
rect 614 1558 618 1562
rect 654 1558 658 1562
rect 926 1558 930 1562
rect 998 1558 1002 1562
rect 1358 1558 1362 1562
rect 1374 1558 1378 1562
rect 1446 1558 1450 1562
rect 1454 1558 1458 1562
rect 1478 1558 1482 1562
rect 1494 1558 1498 1562
rect 1670 1558 1674 1562
rect 1878 1558 1882 1562
rect 1934 1558 1938 1562
rect 1990 1558 1994 1562
rect 2270 1558 2274 1562
rect 2302 1558 2306 1562
rect 2622 1558 2626 1562
rect 2806 1558 2810 1562
rect 2862 1558 2866 1562
rect 2910 1558 2914 1562
rect 3030 1558 3034 1562
rect 3190 1558 3194 1562
rect 3318 1558 3322 1562
rect 3358 1558 3362 1562
rect 326 1548 330 1552
rect 366 1548 370 1552
rect 414 1548 418 1552
rect 422 1548 426 1552
rect 446 1548 450 1552
rect 454 1548 458 1552
rect 502 1547 506 1551
rect 702 1547 706 1551
rect 838 1547 842 1551
rect 870 1548 874 1552
rect 902 1548 906 1552
rect 958 1548 962 1552
rect 982 1548 986 1552
rect 990 1548 994 1552
rect 1022 1548 1026 1552
rect 1030 1548 1034 1552
rect 1054 1548 1058 1552
rect 1086 1548 1090 1552
rect 1142 1548 1146 1552
rect 1158 1548 1162 1552
rect 1182 1548 1186 1552
rect 1190 1548 1194 1552
rect 1262 1548 1266 1552
rect 1358 1548 1362 1552
rect 1374 1548 1378 1552
rect 1398 1548 1402 1552
rect 1422 1548 1426 1552
rect 1502 1548 1506 1552
rect 1534 1548 1538 1552
rect 1558 1548 1562 1552
rect 1566 1548 1570 1552
rect 1590 1548 1594 1552
rect 1598 1548 1602 1552
rect 1622 1548 1626 1552
rect 1662 1548 1666 1552
rect 1678 1548 1682 1552
rect 1694 1548 1698 1552
rect 1702 1548 1706 1552
rect 1710 1548 1714 1552
rect 1734 1548 1738 1552
rect 1758 1548 1762 1552
rect 1782 1548 1786 1552
rect 1790 1548 1794 1552
rect 1806 1548 1810 1552
rect 1830 1548 1834 1552
rect 1838 1548 1842 1552
rect 1894 1548 1898 1552
rect 1902 1548 1906 1552
rect 1918 1548 1922 1552
rect 1950 1548 1954 1552
rect 1966 1548 1970 1552
rect 2006 1548 2010 1552
rect 2030 1548 2034 1552
rect 2038 1548 2042 1552
rect 2054 1548 2058 1552
rect 2078 1548 2082 1552
rect 2086 1548 2090 1552
rect 2110 1548 2114 1552
rect 2142 1548 2146 1552
rect 2150 1548 2154 1552
rect 2158 1548 2162 1552
rect 2190 1548 2194 1552
rect 2198 1548 2202 1552
rect 2206 1548 2210 1552
rect 2238 1548 2242 1552
rect 2246 1548 2250 1552
rect 2286 1548 2290 1552
rect 2334 1548 2338 1552
rect 2342 1548 2346 1552
rect 2398 1548 2402 1552
rect 2406 1548 2410 1552
rect 2454 1548 2458 1552
rect 2486 1548 2490 1552
rect 2526 1548 2530 1552
rect 2550 1548 2554 1552
rect 2630 1548 2634 1552
rect 2646 1548 2650 1552
rect 2654 1548 2658 1552
rect 2686 1548 2690 1552
rect 2718 1548 2722 1552
rect 2750 1548 2754 1552
rect 2790 1548 2794 1552
rect 2846 1548 2850 1552
rect 2862 1548 2866 1552
rect 2934 1548 2938 1552
rect 2966 1548 2970 1552
rect 2982 1548 2986 1552
rect 3070 1548 3074 1552
rect 3086 1548 3090 1552
rect 3126 1548 3130 1552
rect 3134 1548 3138 1552
rect 3150 1548 3154 1552
rect 3174 1548 3178 1552
rect 3182 1548 3186 1552
rect 3206 1548 3210 1552
rect 3254 1548 3258 1552
rect 3342 1548 3346 1552
rect 3358 1548 3362 1552
rect 3542 1558 3546 1562
rect 3558 1558 3562 1562
rect 3734 1558 3738 1562
rect 3790 1558 3794 1562
rect 3806 1558 3810 1562
rect 3974 1558 3978 1562
rect 4054 1558 4058 1562
rect 4150 1558 4154 1562
rect 4302 1558 4306 1562
rect 4350 1558 4354 1562
rect 4630 1558 4634 1562
rect 3398 1548 3402 1552
rect 110 1538 114 1542
rect 166 1538 170 1542
rect 278 1538 282 1542
rect 334 1538 338 1542
rect 390 1538 394 1542
rect 422 1538 426 1542
rect 486 1538 490 1542
rect 606 1538 610 1542
rect 630 1538 634 1542
rect 670 1538 674 1542
rect 686 1538 690 1542
rect 830 1538 834 1542
rect 878 1538 882 1542
rect 894 1538 898 1542
rect 926 1538 930 1542
rect 942 1538 946 1542
rect 1014 1538 1018 1542
rect 1118 1538 1122 1542
rect 1198 1538 1202 1542
rect 1230 1538 1234 1542
rect 1318 1538 1322 1542
rect 1366 1538 1370 1542
rect 1398 1538 1402 1542
rect 1470 1538 1474 1542
rect 1638 1538 1642 1542
rect 1694 1538 1698 1542
rect 1798 1538 1802 1542
rect 1870 1538 1874 1542
rect 3494 1547 3498 1551
rect 3526 1548 3530 1552
rect 3542 1548 3546 1552
rect 3582 1548 3586 1552
rect 3590 1548 3594 1552
rect 3614 1548 3618 1552
rect 3670 1548 3674 1552
rect 3750 1548 3754 1552
rect 3782 1548 3786 1552
rect 3822 1548 3826 1552
rect 3846 1548 3850 1552
rect 3854 1548 3858 1552
rect 3862 1548 3866 1552
rect 3918 1548 3922 1552
rect 3934 1548 3938 1552
rect 3958 1548 3962 1552
rect 3966 1548 3970 1552
rect 3990 1548 3994 1552
rect 4014 1548 4018 1552
rect 4038 1548 4042 1552
rect 4046 1548 4050 1552
rect 4078 1548 4082 1552
rect 4094 1548 4098 1552
rect 4118 1548 4122 1552
rect 4134 1548 4138 1552
rect 4166 1548 4170 1552
rect 1942 1538 1946 1542
rect 1974 1538 1978 1542
rect 2214 1538 2218 1542
rect 2254 1538 2258 1542
rect 2278 1538 2282 1542
rect 2358 1538 2362 1542
rect 2374 1538 2378 1542
rect 2614 1538 2618 1542
rect 2646 1538 2650 1542
rect 2758 1538 2762 1542
rect 2782 1538 2786 1542
rect 2822 1538 2826 1542
rect 2878 1538 2882 1542
rect 2926 1538 2930 1542
rect 3046 1538 3050 1542
rect 3214 1538 3218 1542
rect 3230 1538 3234 1542
rect 3342 1538 3346 1542
rect 3350 1538 3354 1542
rect 3406 1538 3410 1542
rect 3510 1538 3514 1542
rect 3550 1538 3554 1542
rect 3582 1538 3586 1542
rect 3662 1538 3666 1542
rect 3758 1538 3762 1542
rect 4246 1547 4250 1551
rect 4286 1548 4290 1552
rect 4310 1548 4314 1552
rect 4334 1548 4338 1552
rect 4350 1548 4354 1552
rect 4358 1548 4362 1552
rect 4366 1548 4370 1552
rect 4390 1548 4394 1552
rect 4462 1548 4466 1552
rect 4574 1548 4578 1552
rect 4670 1558 4674 1562
rect 4822 1558 4826 1562
rect 4846 1558 4850 1562
rect 4670 1548 4674 1552
rect 4710 1547 4714 1551
rect 4790 1548 4794 1552
rect 4806 1548 4810 1552
rect 4854 1548 4858 1552
rect 4934 1548 4938 1552
rect 4974 1548 4978 1552
rect 5006 1548 5010 1552
rect 5022 1548 5026 1552
rect 5078 1558 5082 1562
rect 5054 1548 5058 1552
rect 5078 1548 5082 1552
rect 5150 1548 5154 1552
rect 3926 1538 3930 1542
rect 3998 1538 4002 1542
rect 4078 1538 4082 1542
rect 4142 1538 4146 1542
rect 4174 1538 4178 1542
rect 4262 1538 4266 1542
rect 4278 1538 4282 1542
rect 4486 1538 4490 1542
rect 4574 1538 4578 1542
rect 4614 1538 4618 1542
rect 4678 1538 4682 1542
rect 4694 1538 4698 1542
rect 4718 1538 4722 1542
rect 4814 1538 4818 1542
rect 4830 1538 4834 1542
rect 4958 1538 4962 1542
rect 4982 1538 4986 1542
rect 5046 1538 5050 1542
rect 5054 1538 5058 1542
rect 5094 1538 5098 1542
rect 5158 1538 5162 1542
rect 150 1528 154 1532
rect 342 1528 346 1532
rect 470 1528 474 1532
rect 638 1528 642 1532
rect 974 1528 978 1532
rect 1406 1528 1410 1532
rect 1518 1528 1522 1532
rect 1550 1528 1554 1532
rect 1846 1528 1850 1532
rect 1862 1528 1866 1532
rect 2134 1528 2138 1532
rect 2422 1528 2426 1532
rect 2518 1528 2522 1532
rect 2670 1528 2674 1532
rect 2774 1528 2778 1532
rect 2902 1528 2906 1532
rect 2950 1528 2954 1532
rect 2958 1528 2962 1532
rect 2998 1528 3002 1532
rect 3006 1528 3010 1532
rect 3014 1528 3018 1532
rect 3038 1528 3042 1532
rect 3054 1528 3058 1532
rect 3422 1528 3426 1532
rect 3766 1528 3770 1532
rect 3886 1528 3890 1532
rect 4310 1528 4314 1532
rect 5022 1528 5026 1532
rect 262 1518 266 1522
rect 566 1518 570 1522
rect 766 1518 770 1522
rect 1214 1518 1218 1522
rect 1878 1518 1882 1522
rect 2270 1518 2274 1522
rect 2318 1518 2322 1522
rect 2438 1518 2442 1522
rect 2470 1518 2474 1522
rect 2702 1518 2706 1522
rect 2734 1518 2738 1522
rect 2766 1518 2770 1522
rect 2870 1518 2874 1522
rect 2894 1518 2898 1522
rect 2910 1518 2914 1522
rect 3062 1518 3066 1522
rect 3726 1518 3730 1522
rect 3734 1518 3738 1522
rect 3910 1518 3914 1522
rect 3974 1518 3978 1522
rect 4054 1518 4058 1522
rect 4502 1518 4506 1522
rect 4862 1518 4866 1522
rect 4990 1518 4994 1522
rect 5030 1518 5034 1522
rect 1050 1503 1054 1507
rect 1057 1503 1061 1507
rect 2074 1503 2078 1507
rect 2081 1503 2085 1507
rect 3098 1503 3102 1507
rect 3105 1503 3109 1507
rect 4114 1503 4118 1507
rect 4121 1503 4125 1507
rect 94 1488 98 1492
rect 182 1488 186 1492
rect 254 1488 258 1492
rect 382 1488 386 1492
rect 446 1488 450 1492
rect 622 1488 626 1492
rect 670 1488 674 1492
rect 702 1488 706 1492
rect 750 1488 754 1492
rect 774 1488 778 1492
rect 966 1488 970 1492
rect 1174 1488 1178 1492
rect 1222 1488 1226 1492
rect 1414 1488 1418 1492
rect 1438 1488 1442 1492
rect 1494 1488 1498 1492
rect 1670 1488 1674 1492
rect 1686 1488 1690 1492
rect 1806 1488 1810 1492
rect 1918 1488 1922 1492
rect 1934 1488 1938 1492
rect 1974 1488 1978 1492
rect 1982 1488 1986 1492
rect 2118 1488 2122 1492
rect 2158 1488 2162 1492
rect 2214 1488 2218 1492
rect 2430 1488 2434 1492
rect 2454 1488 2458 1492
rect 2566 1488 2570 1492
rect 2638 1488 2642 1492
rect 2670 1488 2674 1492
rect 2806 1488 2810 1492
rect 2822 1488 2826 1492
rect 2926 1488 2930 1492
rect 2966 1488 2970 1492
rect 3030 1488 3034 1492
rect 3190 1488 3194 1492
rect 3246 1488 3250 1492
rect 3366 1488 3370 1492
rect 3446 1488 3450 1492
rect 3534 1488 3538 1492
rect 3646 1488 3650 1492
rect 3670 1488 3674 1492
rect 3694 1488 3698 1492
rect 3846 1488 3850 1492
rect 3966 1488 3970 1492
rect 3982 1488 3986 1492
rect 4102 1488 4106 1492
rect 4238 1488 4242 1492
rect 4286 1488 4290 1492
rect 4382 1488 4386 1492
rect 4406 1488 4410 1492
rect 4526 1488 4530 1492
rect 4558 1488 4562 1492
rect 4766 1488 4770 1492
rect 4886 1488 4890 1492
rect 4910 1488 4914 1492
rect 5054 1488 5058 1492
rect 5094 1488 5098 1492
rect 190 1478 194 1482
rect 214 1478 218 1482
rect 102 1468 106 1472
rect 158 1468 162 1472
rect 174 1468 178 1472
rect 406 1478 410 1482
rect 574 1478 578 1482
rect 734 1478 738 1482
rect 1910 1478 1914 1482
rect 2278 1478 2282 1482
rect 2422 1478 2426 1482
rect 2518 1478 2522 1482
rect 2814 1478 2818 1482
rect 2934 1478 2938 1482
rect 3046 1478 3050 1482
rect 3102 1478 3106 1482
rect 3110 1478 3114 1482
rect 3158 1478 3162 1482
rect 3182 1478 3186 1482
rect 3222 1478 3226 1482
rect 3542 1478 3546 1482
rect 4254 1478 4258 1482
rect 4366 1478 4370 1482
rect 238 1468 242 1472
rect 278 1468 282 1472
rect 294 1468 298 1472
rect 398 1468 402 1472
rect 454 1468 458 1472
rect 494 1468 498 1472
rect 598 1468 602 1472
rect 654 1468 658 1472
rect 678 1468 682 1472
rect 694 1468 698 1472
rect 758 1468 762 1472
rect 766 1468 770 1472
rect 790 1468 794 1472
rect 830 1468 834 1472
rect 934 1468 938 1472
rect 942 1468 946 1472
rect 982 1468 986 1472
rect 1086 1468 1090 1472
rect 1118 1468 1122 1472
rect 1150 1468 1154 1472
rect 1166 1468 1170 1472
rect 1198 1468 1202 1472
rect 1254 1468 1258 1472
rect 1302 1468 1306 1472
rect 1390 1468 1394 1472
rect 1422 1468 1426 1472
rect 1470 1468 1474 1472
rect 1478 1468 1482 1472
rect 1502 1468 1506 1472
rect 1590 1468 1594 1472
rect 1678 1468 1682 1472
rect 1710 1468 1714 1472
rect 1766 1468 1770 1472
rect 1782 1468 1786 1472
rect 1870 1468 1874 1472
rect 1926 1468 1930 1472
rect 1950 1468 1954 1472
rect 2086 1468 2090 1472
rect 2094 1468 2098 1472
rect 2150 1468 2154 1472
rect 2182 1468 2186 1472
rect 2190 1468 2194 1472
rect 2246 1468 2250 1472
rect 2358 1468 2362 1472
rect 2438 1468 2442 1472
rect 2630 1468 2634 1472
rect 2846 1468 2850 1472
rect 2974 1468 2978 1472
rect 3038 1468 3042 1472
rect 3070 1468 3074 1472
rect 3094 1468 3098 1472
rect 3110 1468 3114 1472
rect 3134 1468 3138 1472
rect 3150 1468 3154 1472
rect 3230 1468 3234 1472
rect 3334 1468 3338 1472
rect 3350 1468 3354 1472
rect 3398 1468 3402 1472
rect 38 1458 42 1462
rect 62 1458 66 1462
rect 110 1458 114 1462
rect 118 1458 122 1462
rect 150 1458 154 1462
rect 166 1458 170 1462
rect 198 1458 202 1462
rect 246 1458 250 1462
rect 270 1458 274 1462
rect 310 1459 314 1463
rect 430 1458 434 1462
rect 462 1458 466 1462
rect 518 1458 522 1462
rect 606 1458 610 1462
rect 646 1458 650 1462
rect 686 1458 690 1462
rect 718 1458 722 1462
rect 798 1458 802 1462
rect 814 1458 818 1462
rect 846 1459 850 1463
rect 878 1458 882 1462
rect 950 1458 954 1462
rect 1006 1458 1010 1462
rect 1094 1458 1098 1462
rect 1134 1458 1138 1462
rect 1198 1458 1202 1462
rect 1206 1458 1210 1462
rect 1286 1458 1290 1462
rect 1334 1458 1338 1462
rect 1398 1458 1402 1462
rect 1446 1458 1450 1462
rect 1462 1458 1466 1462
rect 1510 1458 1514 1462
rect 1534 1458 1538 1462
rect 1630 1458 1634 1462
rect 1702 1458 1706 1462
rect 1734 1458 1738 1462
rect 1742 1458 1746 1462
rect 1750 1458 1754 1462
rect 1790 1458 1794 1462
rect 1878 1459 1882 1463
rect 1958 1458 1962 1462
rect 2014 1458 2018 1462
rect 2038 1458 2042 1462
rect 2102 1458 2106 1462
rect 2150 1458 2154 1462
rect 2190 1458 2194 1462
rect 2246 1458 2250 1462
rect 2254 1458 2258 1462
rect 2262 1458 2266 1462
rect 2334 1458 2338 1462
rect 2414 1458 2418 1462
rect 2446 1458 2450 1462
rect 2486 1458 2490 1462
rect 2510 1458 2514 1462
rect 2550 1458 2554 1462
rect 2622 1458 2626 1462
rect 2654 1458 2658 1462
rect 2686 1458 2690 1462
rect 2766 1458 2770 1462
rect 2774 1458 2778 1462
rect 2830 1458 2834 1462
rect 2870 1458 2874 1462
rect 2950 1458 2954 1462
rect 2982 1458 2986 1462
rect 3022 1458 3026 1462
rect 3158 1458 3162 1462
rect 3174 1458 3178 1462
rect 3198 1458 3202 1462
rect 3206 1458 3210 1462
rect 3318 1459 3322 1463
rect 3430 1468 3434 1472
rect 3438 1468 3442 1472
rect 3462 1468 3466 1472
rect 3518 1468 3522 1472
rect 3574 1468 3578 1472
rect 3606 1468 3610 1472
rect 3662 1468 3666 1472
rect 3686 1468 3690 1472
rect 3710 1468 3714 1472
rect 3822 1468 3826 1472
rect 3838 1468 3842 1472
rect 3862 1468 3866 1472
rect 3894 1468 3898 1472
rect 3950 1468 3954 1472
rect 3958 1468 3962 1472
rect 4094 1468 4098 1472
rect 4142 1468 4146 1472
rect 4246 1468 4250 1472
rect 4318 1468 4322 1472
rect 4694 1478 4698 1482
rect 4726 1478 4730 1482
rect 4878 1478 4882 1482
rect 5158 1478 5162 1482
rect 4390 1468 4394 1472
rect 4486 1468 4490 1472
rect 4502 1468 4506 1472
rect 4550 1468 4554 1472
rect 4622 1468 4626 1472
rect 4670 1468 4674 1472
rect 4734 1468 4738 1472
rect 4798 1468 4802 1472
rect 4846 1468 4850 1472
rect 4854 1468 4858 1472
rect 4894 1468 4898 1472
rect 4934 1468 4938 1472
rect 4942 1468 4946 1472
rect 4958 1468 4962 1472
rect 5014 1468 5018 1472
rect 5062 1468 5066 1472
rect 5086 1468 5090 1472
rect 3390 1458 3394 1462
rect 3406 1458 3410 1462
rect 3422 1458 3426 1462
rect 3470 1458 3474 1462
rect 3510 1458 3514 1462
rect 3526 1458 3530 1462
rect 3566 1458 3570 1462
rect 3622 1458 3626 1462
rect 3630 1458 3634 1462
rect 3718 1458 3722 1462
rect 3734 1458 3738 1462
rect 3806 1459 3810 1463
rect 3870 1458 3874 1462
rect 3878 1458 3882 1462
rect 3894 1458 3898 1462
rect 3918 1458 3922 1462
rect 3942 1458 3946 1462
rect 4030 1458 4034 1462
rect 4054 1458 4058 1462
rect 4158 1459 4162 1463
rect 4278 1458 4282 1462
rect 4302 1458 4306 1462
rect 4310 1458 4314 1462
rect 4326 1458 4330 1462
rect 4350 1458 4354 1462
rect 4398 1458 4402 1462
rect 4438 1458 4442 1462
rect 4462 1458 4466 1462
rect 4510 1458 4514 1462
rect 4614 1458 4618 1462
rect 4710 1458 4714 1462
rect 4742 1458 4746 1462
rect 4750 1458 4754 1462
rect 4758 1458 4762 1462
rect 4782 1458 4786 1462
rect 4806 1458 4810 1462
rect 4902 1458 4906 1462
rect 4926 1458 4930 1462
rect 4990 1459 4994 1463
rect 5022 1458 5026 1462
rect 5070 1458 5074 1462
rect 5126 1458 5130 1462
rect 5142 1458 5146 1462
rect 134 1448 138 1452
rect 254 1448 258 1452
rect 382 1448 386 1452
rect 446 1448 450 1452
rect 630 1448 634 1452
rect 662 1448 666 1452
rect 742 1448 746 1452
rect 782 1448 786 1452
rect 814 1448 818 1452
rect 934 1448 938 1452
rect 966 1448 970 1452
rect 1110 1448 1114 1452
rect 1150 1448 1154 1452
rect 1414 1448 1418 1452
rect 1494 1448 1498 1452
rect 1694 1448 1698 1452
rect 1806 1448 1810 1452
rect 1942 1448 1946 1452
rect 1974 1448 1978 1452
rect 2118 1448 2122 1452
rect 2126 1448 2130 1452
rect 2142 1448 2146 1452
rect 2158 1448 2162 1452
rect 2206 1448 2210 1452
rect 2214 1448 2218 1452
rect 2270 1448 2274 1452
rect 2646 1448 2650 1452
rect 3022 1448 3026 1452
rect 3054 1448 3058 1452
rect 3094 1448 3098 1452
rect 3150 1448 3154 1452
rect 3374 1448 3378 1452
rect 3390 1448 3394 1452
rect 3406 1448 3410 1452
rect 3454 1448 3458 1452
rect 3566 1448 3570 1452
rect 3582 1448 3586 1452
rect 3678 1448 3682 1452
rect 3702 1448 3706 1452
rect 3854 1448 3858 1452
rect 3926 1448 3930 1452
rect 3974 1448 3978 1452
rect 4118 1448 4122 1452
rect 4262 1448 4266 1452
rect 4326 1448 4330 1452
rect 4342 1448 4346 1452
rect 4534 1448 4538 1452
rect 4686 1448 4690 1452
rect 4806 1448 4810 1452
rect 4822 1448 4826 1452
rect 4830 1448 4834 1452
rect 4854 1448 4858 1452
rect 4910 1448 4914 1452
rect 4950 1448 4954 1452
rect 4958 1448 4962 1452
rect 5086 1448 5090 1452
rect 478 1438 482 1442
rect 1062 1438 1066 1442
rect 1238 1438 1242 1442
rect 1382 1438 1386 1442
rect 1438 1438 1442 1442
rect 1526 1438 1530 1442
rect 1814 1438 1818 1442
rect 2310 1438 2314 1442
rect 3254 1438 3258 1442
rect 3366 1438 3370 1442
rect 3494 1438 3498 1442
rect 3550 1438 3554 1442
rect 3886 1438 3890 1442
rect 3902 1438 3906 1442
rect 4574 1438 4578 1442
rect 4870 1438 4874 1442
rect 374 1428 378 1432
rect 222 1418 226 1422
rect 462 1418 466 1422
rect 910 1418 914 1422
rect 1246 1418 1250 1422
rect 1270 1418 1274 1422
rect 1510 1418 1514 1422
rect 1550 1418 1554 1422
rect 1670 1418 1674 1422
rect 2198 1418 2202 1422
rect 2398 1418 2402 1422
rect 2566 1418 2570 1422
rect 2606 1418 2610 1422
rect 2670 1418 2674 1422
rect 2702 1418 2706 1422
rect 2998 1418 3002 1422
rect 3126 1418 3130 1422
rect 3214 1418 3218 1422
rect 3470 1418 3474 1422
rect 3598 1418 3602 1422
rect 3718 1418 3722 1422
rect 3942 1418 3946 1422
rect 4678 1418 4682 1422
rect 4838 1418 4842 1422
rect 538 1403 542 1407
rect 545 1403 549 1407
rect 1562 1403 1566 1407
rect 1569 1403 1573 1407
rect 2586 1403 2590 1407
rect 2593 1403 2597 1407
rect 3610 1403 3614 1407
rect 3617 1403 3621 1407
rect 4634 1403 4638 1407
rect 4641 1403 4645 1407
rect 174 1388 178 1392
rect 270 1388 274 1392
rect 526 1388 530 1392
rect 566 1388 570 1392
rect 806 1388 810 1392
rect 966 1388 970 1392
rect 1014 1388 1018 1392
rect 1366 1388 1370 1392
rect 1534 1388 1538 1392
rect 1606 1388 1610 1392
rect 1638 1388 1642 1392
rect 1678 1388 1682 1392
rect 1958 1388 1962 1392
rect 1990 1388 1994 1392
rect 2038 1388 2042 1392
rect 2654 1388 2658 1392
rect 2966 1388 2970 1392
rect 3070 1388 3074 1392
rect 3198 1388 3202 1392
rect 3534 1388 3538 1392
rect 3542 1388 3546 1392
rect 3814 1388 3818 1392
rect 3854 1388 3858 1392
rect 3910 1388 3914 1392
rect 4022 1388 4026 1392
rect 4102 1388 4106 1392
rect 5086 1388 5090 1392
rect 94 1378 98 1382
rect 2926 1378 2930 1382
rect 134 1368 138 1372
rect 286 1368 290 1372
rect 310 1368 314 1372
rect 830 1368 834 1372
rect 870 1368 874 1372
rect 1094 1368 1098 1372
rect 1110 1368 1114 1372
rect 1206 1368 1210 1372
rect 1710 1368 1714 1372
rect 2486 1368 2490 1372
rect 2742 1368 2746 1372
rect 2958 1368 2962 1372
rect 3062 1368 3066 1372
rect 3414 1368 3418 1372
rect 3926 1368 3930 1372
rect 4622 1368 4626 1372
rect 102 1358 106 1362
rect 46 1348 50 1352
rect 62 1348 66 1352
rect 102 1348 106 1352
rect 118 1348 122 1352
rect 134 1348 138 1352
rect 150 1348 154 1352
rect 222 1348 226 1352
rect 286 1348 290 1352
rect 326 1348 330 1352
rect 350 1348 354 1352
rect 374 1358 378 1362
rect 430 1358 434 1362
rect 550 1358 554 1362
rect 582 1358 586 1362
rect 598 1358 602 1362
rect 622 1358 626 1362
rect 390 1348 394 1352
rect 414 1348 418 1352
rect 430 1348 434 1352
rect 462 1347 466 1351
rect 566 1348 570 1352
rect 598 1348 602 1352
rect 670 1348 674 1352
rect 694 1347 698 1351
rect 734 1348 738 1352
rect 758 1358 762 1362
rect 846 1358 850 1362
rect 854 1358 858 1362
rect 910 1358 914 1362
rect 1078 1358 1082 1362
rect 1230 1358 1234 1362
rect 1270 1358 1274 1362
rect 1350 1358 1354 1362
rect 1438 1358 1442 1362
rect 1654 1358 1658 1362
rect 1822 1358 1826 1362
rect 1838 1358 1842 1362
rect 1854 1358 1858 1362
rect 2086 1358 2090 1362
rect 2214 1358 2218 1362
rect 2286 1358 2290 1362
rect 2294 1358 2298 1362
rect 2310 1358 2314 1362
rect 2326 1358 2330 1362
rect 2470 1358 2474 1362
rect 2614 1358 2618 1362
rect 2862 1358 2866 1362
rect 2942 1358 2946 1362
rect 3190 1358 3194 1362
rect 3278 1358 3282 1362
rect 3654 1358 3658 1362
rect 3670 1358 3674 1362
rect 3798 1358 3802 1362
rect 3878 1358 3882 1362
rect 3894 1358 3898 1362
rect 4054 1358 4058 1362
rect 4166 1358 4170 1362
rect 806 1348 810 1352
rect 902 1348 906 1352
rect 918 1348 922 1352
rect 926 1348 930 1352
rect 942 1348 946 1352
rect 950 1348 954 1352
rect 974 1348 978 1352
rect 998 1348 1002 1352
rect 1022 1348 1026 1352
rect 1030 1348 1034 1352
rect 1054 1348 1058 1352
rect 1078 1348 1082 1352
rect 1094 1348 1098 1352
rect 126 1338 130 1342
rect 166 1338 170 1342
rect 190 1338 194 1342
rect 278 1338 282 1342
rect 334 1338 338 1342
rect 342 1338 346 1342
rect 358 1338 362 1342
rect 398 1338 402 1342
rect 406 1338 410 1342
rect 574 1338 578 1342
rect 726 1338 730 1342
rect 742 1338 746 1342
rect 774 1338 778 1342
rect 798 1338 802 1342
rect 830 1338 834 1342
rect 870 1338 874 1342
rect 878 1338 882 1342
rect 934 1338 938 1342
rect 1054 1338 1058 1342
rect 1142 1347 1146 1351
rect 1238 1348 1242 1352
rect 1286 1348 1290 1352
rect 1310 1348 1314 1352
rect 1334 1348 1338 1352
rect 1342 1348 1346 1352
rect 1366 1348 1370 1352
rect 1406 1348 1410 1352
rect 1422 1348 1426 1352
rect 1438 1348 1442 1352
rect 1470 1347 1474 1351
rect 1494 1348 1498 1352
rect 1582 1348 1586 1352
rect 1590 1348 1594 1352
rect 1614 1348 1618 1352
rect 1638 1348 1642 1352
rect 1654 1348 1658 1352
rect 1694 1348 1698 1352
rect 1702 1348 1706 1352
rect 1710 1348 1714 1352
rect 1726 1348 1730 1352
rect 1742 1348 1746 1352
rect 1758 1348 1762 1352
rect 1766 1348 1770 1352
rect 1798 1348 1802 1352
rect 1806 1348 1810 1352
rect 1838 1348 1842 1352
rect 1894 1348 1898 1352
rect 1982 1348 1986 1352
rect 2006 1348 2010 1352
rect 2014 1348 2018 1352
rect 2030 1348 2034 1352
rect 2054 1348 2058 1352
rect 2062 1348 2066 1352
rect 2070 1348 2074 1352
rect 2110 1348 2114 1352
rect 2158 1348 2162 1352
rect 2214 1348 2218 1352
rect 2238 1348 2242 1352
rect 2270 1348 2274 1352
rect 2318 1348 2322 1352
rect 2342 1348 2346 1352
rect 2350 1348 2354 1352
rect 2430 1348 2434 1352
rect 2510 1348 2514 1352
rect 2542 1348 2546 1352
rect 2550 1348 2554 1352
rect 2558 1348 2562 1352
rect 2590 1348 2594 1352
rect 2638 1348 2642 1352
rect 2646 1348 2650 1352
rect 2670 1348 2674 1352
rect 2702 1348 2706 1352
rect 2718 1348 2722 1352
rect 2734 1348 2738 1352
rect 2774 1348 2778 1352
rect 2782 1348 2786 1352
rect 2846 1348 2850 1352
rect 2862 1348 2866 1352
rect 2870 1348 2874 1352
rect 2886 1348 2890 1352
rect 2902 1348 2906 1352
rect 2934 1348 2938 1352
rect 2950 1348 2954 1352
rect 3006 1348 3010 1352
rect 3126 1348 3130 1352
rect 1086 1338 1090 1342
rect 1214 1338 1218 1342
rect 1294 1338 1298 1342
rect 1374 1338 1378 1342
rect 1390 1338 1394 1342
rect 1414 1338 1418 1342
rect 1558 1338 1562 1342
rect 1630 1338 1634 1342
rect 1734 1338 1738 1342
rect 1790 1338 1794 1342
rect 1814 1338 1818 1342
rect 1830 1338 1834 1342
rect 1870 1338 1874 1342
rect 1942 1338 1946 1342
rect 2110 1338 2114 1342
rect 2126 1338 2130 1342
rect 2174 1338 2178 1342
rect 2318 1338 2322 1342
rect 3350 1347 3354 1351
rect 3382 1348 3386 1352
rect 3438 1348 3442 1352
rect 3470 1347 3474 1351
rect 3502 1348 3506 1352
rect 3574 1348 3578 1352
rect 3598 1348 3602 1352
rect 3670 1348 3674 1352
rect 3734 1348 3738 1352
rect 3758 1348 3762 1352
rect 3822 1348 3826 1352
rect 3830 1348 3834 1352
rect 3838 1348 3842 1352
rect 3862 1348 3866 1352
rect 3902 1348 3906 1352
rect 3966 1348 3970 1352
rect 4014 1348 4018 1352
rect 4038 1348 4042 1352
rect 4046 1348 4050 1352
rect 4070 1348 4074 1352
rect 4094 1348 4098 1352
rect 4118 1348 4122 1352
rect 4126 1348 4130 1352
rect 4190 1358 4194 1362
rect 4190 1348 4194 1352
rect 4206 1348 4210 1352
rect 4230 1348 4234 1352
rect 4254 1358 4258 1362
rect 4542 1358 4546 1362
rect 4670 1358 4674 1362
rect 4686 1358 4690 1362
rect 4830 1358 4834 1362
rect 5038 1358 5042 1362
rect 5054 1358 5058 1362
rect 4334 1348 4338 1352
rect 4430 1348 4434 1352
rect 4486 1348 4490 1352
rect 4518 1348 4522 1352
rect 4582 1348 4586 1352
rect 4670 1348 4674 1352
rect 2454 1338 2458 1342
rect 2486 1338 2490 1342
rect 2534 1338 2538 1342
rect 2606 1338 2610 1342
rect 2630 1338 2634 1342
rect 2726 1338 2730 1342
rect 2838 1338 2842 1342
rect 2878 1338 2882 1342
rect 2910 1338 2914 1342
rect 2926 1338 2930 1342
rect 3006 1338 3010 1342
rect 3134 1338 3138 1342
rect 3206 1338 3210 1342
rect 3214 1338 3218 1342
rect 3262 1338 3266 1342
rect 3318 1338 3322 1342
rect 3422 1338 3426 1342
rect 3438 1338 3442 1342
rect 3646 1338 3650 1342
rect 3822 1338 3826 1342
rect 3902 1338 3906 1342
rect 3974 1338 3978 1342
rect 4054 1338 4058 1342
rect 4078 1338 4082 1342
rect 4150 1338 4154 1342
rect 4198 1338 4202 1342
rect 4734 1347 4738 1351
rect 4806 1348 4810 1352
rect 4814 1348 4818 1352
rect 4830 1348 4834 1352
rect 4894 1348 4898 1352
rect 4950 1348 4954 1352
rect 4998 1348 5002 1352
rect 5006 1348 5010 1352
rect 5054 1348 5058 1352
rect 5126 1348 5130 1352
rect 5142 1348 5146 1352
rect 4270 1338 4274 1342
rect 4326 1338 4330 1342
rect 4438 1338 4442 1342
rect 4510 1338 4514 1342
rect 4526 1338 4530 1342
rect 4654 1338 4658 1342
rect 4694 1338 4698 1342
rect 4718 1338 4722 1342
rect 4838 1338 4842 1342
rect 4934 1338 4938 1342
rect 4950 1338 4954 1342
rect 5014 1338 5018 1342
rect 5030 1338 5034 1342
rect 5062 1338 5066 1342
rect 5166 1338 5170 1342
rect 166 1328 170 1332
rect 462 1328 466 1332
rect 782 1328 786 1332
rect 1142 1328 1146 1332
rect 1270 1328 1274 1332
rect 1550 1328 1554 1332
rect 1742 1328 1746 1332
rect 1886 1328 1890 1332
rect 1966 1328 1970 1332
rect 2246 1328 2250 1332
rect 2494 1328 2498 1332
rect 2686 1328 2690 1332
rect 2894 1328 2898 1332
rect 3078 1328 3082 1332
rect 3134 1328 3138 1332
rect 3166 1328 3170 1332
rect 3182 1328 3186 1332
rect 3222 1328 3226 1332
rect 4206 1328 4210 1332
rect 4470 1328 4474 1332
rect 4574 1328 4578 1332
rect 4702 1328 4706 1332
rect 4982 1328 4986 1332
rect 5030 1328 5034 1332
rect 790 1318 794 1322
rect 846 1318 850 1322
rect 1230 1318 1234 1322
rect 1254 1318 1258 1322
rect 1326 1318 1330 1322
rect 1750 1318 1754 1322
rect 1950 1318 1954 1322
rect 2206 1318 2210 1322
rect 2286 1318 2290 1322
rect 2326 1318 2330 1322
rect 2526 1318 2530 1322
rect 2622 1318 2626 1322
rect 3110 1318 3114 1322
rect 3174 1318 3178 1322
rect 3190 1318 3194 1322
rect 3246 1318 3250 1322
rect 3278 1318 3282 1322
rect 3294 1318 3298 1322
rect 3686 1318 3690 1322
rect 4246 1318 4250 1322
rect 4278 1318 4282 1322
rect 4374 1318 4378 1322
rect 4502 1318 4506 1322
rect 4542 1318 4546 1322
rect 4638 1318 4642 1322
rect 4798 1318 4802 1322
rect 4966 1318 4970 1322
rect 5046 1318 5050 1322
rect 1050 1303 1054 1307
rect 1057 1303 1061 1307
rect 2074 1303 2078 1307
rect 2081 1303 2085 1307
rect 3098 1303 3102 1307
rect 3105 1303 3109 1307
rect 4114 1303 4118 1307
rect 4121 1303 4125 1307
rect 94 1288 98 1292
rect 190 1288 194 1292
rect 238 1288 242 1292
rect 334 1288 338 1292
rect 350 1288 354 1292
rect 438 1288 442 1292
rect 566 1288 570 1292
rect 614 1288 618 1292
rect 662 1288 666 1292
rect 710 1288 714 1292
rect 726 1288 730 1292
rect 878 1288 882 1292
rect 1046 1288 1050 1292
rect 1190 1288 1194 1292
rect 1326 1288 1330 1292
rect 1334 1288 1338 1292
rect 1430 1288 1434 1292
rect 1478 1288 1482 1292
rect 1734 1288 1738 1292
rect 1918 1288 1922 1292
rect 1942 1288 1946 1292
rect 1990 1288 1994 1292
rect 2030 1288 2034 1292
rect 2102 1288 2106 1292
rect 2126 1288 2130 1292
rect 2142 1288 2146 1292
rect 2166 1288 2170 1292
rect 2198 1288 2202 1292
rect 2214 1288 2218 1292
rect 2310 1288 2314 1292
rect 2414 1288 2418 1292
rect 2478 1288 2482 1292
rect 2694 1288 2698 1292
rect 2838 1288 2842 1292
rect 2926 1288 2930 1292
rect 3150 1288 3154 1292
rect 3222 1288 3226 1292
rect 3246 1288 3250 1292
rect 3310 1288 3314 1292
rect 3342 1288 3346 1292
rect 3414 1288 3418 1292
rect 3662 1288 3666 1292
rect 3766 1288 3770 1292
rect 3790 1288 3794 1292
rect 3830 1288 3834 1292
rect 3870 1288 3874 1292
rect 3990 1288 3994 1292
rect 4158 1288 4162 1292
rect 4270 1288 4274 1292
rect 4334 1288 4338 1292
rect 4358 1288 4362 1292
rect 4430 1288 4434 1292
rect 4478 1288 4482 1292
rect 4486 1288 4490 1292
rect 4606 1288 4610 1292
rect 4710 1288 4714 1292
rect 4734 1288 4738 1292
rect 4758 1288 4762 1292
rect 4782 1288 4786 1292
rect 4894 1288 4898 1292
rect 5014 1288 5018 1292
rect 5182 1288 5186 1292
rect 358 1278 362 1282
rect 454 1278 458 1282
rect 102 1268 106 1272
rect 158 1268 162 1272
rect 182 1268 186 1272
rect 214 1268 218 1272
rect 222 1268 226 1272
rect 254 1268 258 1272
rect 270 1268 274 1272
rect 366 1268 370 1272
rect 398 1268 402 1272
rect 446 1268 450 1272
rect 470 1268 474 1272
rect 590 1268 594 1272
rect 638 1268 642 1272
rect 654 1268 658 1272
rect 678 1278 682 1282
rect 702 1278 706 1282
rect 894 1278 898 1282
rect 982 1278 986 1282
rect 1166 1278 1170 1282
rect 1342 1278 1346 1282
rect 1462 1278 1466 1282
rect 1574 1278 1578 1282
rect 38 1258 42 1262
rect 62 1258 66 1262
rect 110 1258 114 1262
rect 150 1258 154 1262
rect 278 1258 282 1262
rect 342 1258 346 1262
rect 374 1258 378 1262
rect 390 1258 394 1262
rect 510 1258 514 1262
rect 534 1258 538 1262
rect 598 1258 602 1262
rect 646 1258 650 1262
rect 694 1258 698 1262
rect 718 1258 722 1262
rect 758 1258 762 1262
rect 790 1259 794 1263
rect 854 1268 858 1272
rect 950 1268 954 1272
rect 966 1268 970 1272
rect 1070 1268 1074 1272
rect 1102 1268 1106 1272
rect 1158 1268 1162 1272
rect 1182 1268 1186 1272
rect 1198 1268 1202 1272
rect 1206 1268 1210 1272
rect 1350 1268 1354 1272
rect 1382 1268 1386 1272
rect 1470 1268 1474 1272
rect 1526 1268 1530 1272
rect 1614 1268 1618 1272
rect 1630 1268 1634 1272
rect 1654 1268 1658 1272
rect 1670 1268 1674 1272
rect 1686 1268 1690 1272
rect 1710 1278 1714 1282
rect 1886 1268 1890 1272
rect 1926 1268 1930 1272
rect 1958 1278 1962 1282
rect 2422 1278 2426 1282
rect 2590 1278 2594 1282
rect 1982 1268 1986 1272
rect 2022 1268 2026 1272
rect 2054 1268 2058 1272
rect 2078 1268 2082 1272
rect 2158 1268 2162 1272
rect 2182 1268 2186 1272
rect 2190 1268 2194 1272
rect 2238 1268 2242 1272
rect 2246 1268 2250 1272
rect 2270 1268 2274 1272
rect 2302 1268 2306 1272
rect 2350 1268 2354 1272
rect 2390 1268 2394 1272
rect 3214 1278 3218 1282
rect 3270 1278 3274 1282
rect 3318 1278 3322 1282
rect 3374 1278 3378 1282
rect 3838 1278 3842 1282
rect 3974 1278 3978 1282
rect 4302 1278 4306 1282
rect 4390 1278 4394 1282
rect 4638 1278 4642 1282
rect 5086 1278 5090 1282
rect 2630 1268 2634 1272
rect 2678 1268 2682 1272
rect 2774 1268 2778 1272
rect 2806 1268 2810 1272
rect 2822 1268 2826 1272
rect 2942 1268 2946 1272
rect 2990 1268 2994 1272
rect 3006 1268 3010 1272
rect 3102 1268 3106 1272
rect 3126 1268 3130 1272
rect 3158 1268 3162 1272
rect 3190 1268 3194 1272
rect 3246 1268 3250 1272
rect 3262 1268 3266 1272
rect 3302 1268 3306 1272
rect 3334 1268 3338 1272
rect 3438 1268 3442 1272
rect 3446 1268 3450 1272
rect 3470 1268 3474 1272
rect 3574 1268 3578 1272
rect 3614 1268 3618 1272
rect 3702 1268 3706 1272
rect 3734 1268 3738 1272
rect 3814 1268 3818 1272
rect 3894 1268 3898 1272
rect 4030 1268 4034 1272
rect 4070 1268 4074 1272
rect 4086 1268 4090 1272
rect 4102 1268 4106 1272
rect 4134 1268 4138 1272
rect 4238 1268 4242 1272
rect 4342 1268 4346 1272
rect 4438 1268 4442 1272
rect 4462 1268 4466 1272
rect 4566 1268 4570 1272
rect 4582 1268 4586 1272
rect 4702 1268 4706 1272
rect 4726 1268 4730 1272
rect 4750 1268 4754 1272
rect 4766 1268 4770 1272
rect 4878 1268 4882 1272
rect 4934 1268 4938 1272
rect 4974 1268 4978 1272
rect 4990 1268 4994 1272
rect 5038 1268 5042 1272
rect 5102 1268 5106 1272
rect 822 1258 826 1262
rect 830 1258 834 1262
rect 862 1258 866 1262
rect 990 1258 994 1262
rect 1094 1258 1098 1262
rect 1110 1258 1114 1262
rect 1134 1258 1138 1262
rect 1166 1258 1170 1262
rect 1214 1258 1218 1262
rect 1222 1258 1226 1262
rect 1262 1259 1266 1263
rect 1286 1258 1290 1262
rect 1358 1258 1362 1262
rect 1382 1258 1386 1262
rect 1406 1258 1410 1262
rect 1414 1258 1418 1262
rect 1438 1258 1442 1262
rect 1542 1259 1546 1263
rect 1606 1258 1610 1262
rect 1638 1258 1642 1262
rect 1662 1258 1666 1262
rect 1678 1258 1682 1262
rect 1710 1258 1714 1262
rect 1726 1258 1730 1262
rect 1766 1258 1770 1262
rect 1790 1258 1794 1262
rect 1854 1259 1858 1263
rect 1926 1258 1930 1262
rect 1974 1258 1978 1262
rect 2046 1258 2050 1262
rect 2086 1258 2090 1262
rect 2110 1258 2114 1262
rect 2230 1258 2234 1262
rect 2254 1258 2258 1262
rect 2294 1258 2298 1262
rect 2366 1258 2370 1262
rect 2406 1258 2410 1262
rect 2438 1258 2442 1262
rect 2462 1258 2466 1262
rect 2470 1258 2474 1262
rect 2510 1258 2514 1262
rect 2526 1258 2530 1262
rect 2574 1258 2578 1262
rect 2638 1258 2642 1262
rect 2646 1258 2650 1262
rect 2654 1258 2658 1262
rect 2678 1258 2682 1262
rect 2750 1258 2754 1262
rect 2790 1258 2794 1262
rect 2846 1258 2850 1262
rect 2878 1258 2882 1262
rect 2902 1258 2906 1262
rect 2974 1258 2978 1262
rect 2990 1258 2994 1262
rect 3022 1259 3026 1263
rect 3166 1258 3170 1262
rect 3182 1258 3186 1262
rect 3190 1258 3194 1262
rect 3286 1258 3290 1262
rect 3294 1258 3298 1262
rect 3326 1258 3330 1262
rect 3358 1258 3362 1262
rect 3382 1258 3386 1262
rect 3406 1258 3410 1262
rect 3430 1258 3434 1262
rect 3534 1258 3538 1262
rect 3558 1259 3562 1263
rect 3606 1258 3610 1262
rect 3638 1258 3642 1262
rect 3646 1258 3650 1262
rect 3670 1258 3674 1262
rect 3726 1258 3730 1262
rect 3742 1258 3746 1262
rect 3750 1258 3754 1262
rect 3774 1258 3778 1262
rect 3806 1258 3810 1262
rect 3822 1258 3826 1262
rect 3846 1258 3850 1262
rect 3854 1258 3858 1262
rect 3878 1258 3882 1262
rect 3886 1258 3890 1262
rect 3910 1258 3914 1262
rect 3950 1258 3954 1262
rect 4046 1258 4050 1262
rect 4094 1258 4098 1262
rect 4222 1259 4226 1263
rect 4254 1258 4258 1262
rect 4262 1258 4266 1262
rect 4294 1258 4298 1262
rect 4318 1258 4322 1262
rect 4350 1258 4354 1262
rect 4374 1258 4378 1262
rect 4414 1258 4418 1262
rect 4542 1258 4546 1262
rect 4622 1258 4626 1262
rect 4678 1258 4682 1262
rect 4862 1259 4866 1263
rect 4958 1259 4962 1263
rect 5030 1258 5034 1262
rect 5062 1258 5066 1262
rect 5070 1258 5074 1262
rect 5118 1259 5122 1263
rect 110 1248 114 1252
rect 134 1248 138 1252
rect 166 1248 170 1252
rect 238 1248 242 1252
rect 390 1248 394 1252
rect 454 1248 458 1252
rect 622 1248 626 1252
rect 830 1248 834 1252
rect 846 1248 850 1252
rect 878 1248 882 1252
rect 1110 1248 1114 1252
rect 1126 1248 1130 1252
rect 1134 1248 1138 1252
rect 1182 1248 1186 1252
rect 1230 1248 1234 1252
rect 1398 1248 1402 1252
rect 1646 1248 1650 1252
rect 1998 1248 2002 1252
rect 2006 1248 2010 1252
rect 2102 1248 2106 1252
rect 2142 1248 2146 1252
rect 2158 1248 2162 1252
rect 2206 1248 2210 1252
rect 2214 1248 2218 1252
rect 2278 1248 2282 1252
rect 2606 1248 2610 1252
rect 2838 1248 2842 1252
rect 2958 1248 2962 1252
rect 3150 1248 3154 1252
rect 3222 1248 3226 1252
rect 3238 1248 3242 1252
rect 3414 1248 3418 1252
rect 3446 1248 3450 1252
rect 3470 1248 3474 1252
rect 3590 1248 3594 1252
rect 3606 1248 3610 1252
rect 3790 1248 3794 1252
rect 4110 1248 4114 1252
rect 4150 1248 4154 1252
rect 4358 1248 4362 1252
rect 4454 1248 4458 1252
rect 4598 1248 4602 1252
rect 4694 1248 4698 1252
rect 4742 1248 4746 1252
rect 5006 1248 5010 1252
rect 5014 1248 5018 1252
rect 5046 1248 5050 1252
rect 5062 1248 5066 1252
rect 406 1238 410 1242
rect 430 1238 434 1242
rect 1454 1238 1458 1242
rect 2454 1238 2458 1242
rect 3182 1238 3186 1242
rect 3206 1238 3210 1242
rect 3462 1238 3466 1242
rect 3686 1238 3690 1242
rect 3726 1238 3730 1242
rect 3918 1238 3922 1242
rect 4006 1238 4010 1242
rect 4478 1238 4482 1242
rect 4726 1238 4730 1242
rect 4774 1238 4778 1242
rect 4790 1238 4794 1242
rect 4814 1238 4818 1242
rect 4798 1228 4802 1232
rect 374 1218 378 1222
rect 2126 1218 2130 1222
rect 2862 1218 2866 1222
rect 2894 1218 2898 1222
rect 3286 1218 3290 1222
rect 3494 1218 3498 1222
rect 3934 1218 3938 1222
rect 4142 1218 4146 1222
rect 4678 1218 4682 1222
rect 4998 1218 5002 1222
rect 538 1203 542 1207
rect 545 1203 549 1207
rect 1562 1203 1566 1207
rect 1569 1203 1573 1207
rect 2586 1203 2590 1207
rect 2593 1203 2597 1207
rect 3610 1203 3614 1207
rect 3617 1203 3621 1207
rect 4634 1203 4638 1207
rect 4641 1203 4645 1207
rect 62 1188 66 1192
rect 166 1188 170 1192
rect 238 1188 242 1192
rect 446 1188 450 1192
rect 462 1188 466 1192
rect 526 1188 530 1192
rect 878 1188 882 1192
rect 974 1188 978 1192
rect 1006 1188 1010 1192
rect 1118 1188 1122 1192
rect 1214 1188 1218 1192
rect 1238 1188 1242 1192
rect 1366 1188 1370 1192
rect 1422 1188 1426 1192
rect 1694 1188 1698 1192
rect 1758 1188 1762 1192
rect 2238 1188 2242 1192
rect 2270 1188 2274 1192
rect 2574 1188 2578 1192
rect 2670 1188 2674 1192
rect 2710 1188 2714 1192
rect 2910 1188 2914 1192
rect 3158 1188 3162 1192
rect 3198 1188 3202 1192
rect 3286 1188 3290 1192
rect 3374 1188 3378 1192
rect 3398 1188 3402 1192
rect 3582 1188 3586 1192
rect 3646 1188 3650 1192
rect 3686 1188 3690 1192
rect 3718 1188 3722 1192
rect 3854 1188 3858 1192
rect 3942 1188 3946 1192
rect 4078 1188 4082 1192
rect 4382 1188 4386 1192
rect 4662 1188 4666 1192
rect 4862 1188 4866 1192
rect 5182 1188 5186 1192
rect 614 1168 618 1172
rect 726 1168 730 1172
rect 742 1168 746 1172
rect 782 1168 786 1172
rect 1534 1168 1538 1172
rect 1590 1168 1594 1172
rect 1806 1168 1810 1172
rect 1870 1168 1874 1172
rect 1934 1168 1938 1172
rect 2446 1168 2450 1172
rect 2734 1168 2738 1172
rect 190 1158 194 1162
rect 206 1158 210 1162
rect 574 1158 578 1162
rect 590 1158 594 1162
rect 630 1158 634 1162
rect 758 1158 762 1162
rect 798 1158 802 1162
rect 1022 1158 1026 1162
rect 1030 1158 1034 1162
rect 1254 1158 1258 1162
rect 1438 1158 1442 1162
rect 1446 1158 1450 1162
rect 1462 1158 1466 1162
rect 1478 1158 1482 1162
rect 110 1148 114 1152
rect 190 1148 194 1152
rect 214 1148 218 1152
rect 222 1148 226 1152
rect 278 1148 282 1152
rect 390 1148 394 1152
rect 470 1148 474 1152
rect 558 1148 562 1152
rect 574 1148 578 1152
rect 606 1148 610 1152
rect 678 1148 682 1152
rect 686 1148 690 1152
rect 742 1148 746 1152
rect 766 1148 770 1152
rect 798 1148 802 1152
rect 846 1148 850 1152
rect 854 1148 858 1152
rect 886 1148 890 1152
rect 894 1148 898 1152
rect 934 1148 938 1152
rect 950 1148 954 1152
rect 958 1148 962 1152
rect 982 1148 986 1152
rect 1006 1148 1010 1152
rect 1038 1148 1042 1152
rect 1046 1148 1050 1152
rect 1078 1148 1082 1152
rect 1150 1148 1154 1152
rect 1238 1148 1242 1152
rect 1294 1148 1298 1152
rect 1390 1148 1394 1152
rect 1422 1148 1426 1152
rect 1462 1148 1466 1152
rect 1478 1148 1482 1152
rect 1494 1148 1498 1152
rect 1518 1148 1522 1152
rect 1558 1158 1562 1162
rect 1734 1158 1738 1162
rect 1790 1158 1794 1162
rect 1558 1148 1562 1152
rect 1646 1148 1650 1152
rect 1694 1148 1698 1152
rect 1750 1148 1754 1152
rect 1774 1148 1778 1152
rect 1782 1148 1786 1152
rect 1806 1148 1810 1152
rect 1846 1148 1850 1152
rect 2102 1158 2106 1162
rect 2118 1158 2122 1162
rect 2158 1158 2162 1162
rect 2406 1158 2410 1162
rect 2422 1158 2426 1162
rect 3742 1168 3746 1172
rect 2462 1158 2466 1162
rect 2622 1158 2626 1162
rect 2726 1158 2730 1162
rect 3502 1158 3506 1162
rect 1902 1148 1906 1152
rect 1926 1148 1930 1152
rect 1966 1148 1970 1152
rect 1990 1148 1994 1152
rect 2054 1148 2058 1152
rect 2086 1148 2090 1152
rect 2102 1148 2106 1152
rect 2118 1148 2122 1152
rect 2174 1148 2178 1152
rect 2190 1148 2194 1152
rect 2254 1148 2258 1152
rect 2278 1148 2282 1152
rect 2342 1148 2346 1152
rect 2390 1148 2394 1152
rect 2422 1148 2426 1152
rect 2510 1148 2514 1152
rect 2526 1148 2530 1152
rect 2638 1148 2642 1152
rect 2662 1148 2666 1152
rect 2686 1148 2690 1152
rect 2694 1148 2698 1152
rect 2710 1148 2714 1152
rect 2766 1148 2770 1152
rect 2782 1148 2786 1152
rect 2798 1148 2802 1152
rect 2838 1148 2842 1152
rect 2846 1148 2850 1152
rect 2926 1148 2930 1152
rect 2934 1148 2938 1152
rect 2950 1148 2954 1152
rect 2966 1148 2970 1152
rect 6 1138 10 1142
rect 86 1138 90 1142
rect 198 1138 202 1142
rect 230 1138 234 1142
rect 246 1138 250 1142
rect 286 1138 290 1142
rect 366 1138 370 1142
rect 550 1138 554 1142
rect 582 1138 586 1142
rect 734 1138 738 1142
rect 790 1138 794 1142
rect 814 1138 818 1142
rect 822 1138 826 1142
rect 998 1138 1002 1142
rect 1054 1138 1058 1142
rect 1158 1138 1162 1142
rect 1230 1138 1234 1142
rect 1470 1138 1474 1142
rect 1502 1138 1506 1142
rect 1510 1138 1514 1142
rect 1566 1138 1570 1142
rect 1686 1138 1690 1142
rect 1718 1138 1722 1142
rect 1838 1138 1842 1142
rect 1894 1138 1898 1142
rect 2078 1138 2082 1142
rect 2110 1138 2114 1142
rect 3014 1147 3018 1151
rect 3150 1148 3154 1152
rect 3174 1148 3178 1152
rect 3206 1148 3210 1152
rect 3214 1148 3218 1152
rect 3222 1148 3226 1152
rect 3254 1148 3258 1152
rect 3262 1148 3266 1152
rect 3278 1148 3282 1152
rect 3302 1148 3306 1152
rect 3310 1148 3314 1152
rect 3342 1148 3346 1152
rect 3350 1148 3354 1152
rect 3358 1148 3362 1152
rect 3382 1148 3386 1152
rect 3462 1147 3466 1151
rect 3502 1148 3506 1152
rect 3526 1158 3530 1162
rect 3726 1158 3730 1162
rect 3774 1158 3778 1162
rect 3878 1158 3882 1162
rect 3910 1158 3914 1162
rect 4054 1158 4058 1162
rect 4110 1158 4114 1162
rect 4198 1158 4202 1162
rect 4214 1158 4218 1162
rect 4342 1158 4346 1162
rect 4470 1158 4474 1162
rect 4494 1158 4498 1162
rect 4574 1158 4578 1162
rect 4622 1158 4626 1162
rect 4694 1158 4698 1162
rect 5006 1158 5010 1162
rect 3542 1148 3546 1152
rect 3574 1148 3578 1152
rect 3606 1148 3610 1152
rect 3630 1148 3634 1152
rect 3670 1148 3674 1152
rect 3694 1148 3698 1152
rect 3710 1148 3714 1152
rect 3758 1148 3762 1152
rect 3774 1148 3778 1152
rect 3790 1148 3794 1152
rect 3814 1148 3818 1152
rect 3822 1148 3826 1152
rect 3838 1148 3842 1152
rect 3862 1148 3866 1152
rect 3870 1148 3874 1152
rect 3886 1148 3890 1152
rect 3902 1148 3906 1152
rect 3918 1148 3922 1152
rect 3926 1148 3930 1152
rect 3982 1148 3986 1152
rect 4054 1148 4058 1152
rect 4070 1148 4074 1152
rect 4094 1148 4098 1152
rect 4142 1148 4146 1152
rect 4158 1148 4162 1152
rect 4190 1148 4194 1152
rect 4214 1148 4218 1152
rect 4302 1148 4306 1152
rect 4366 1148 4370 1152
rect 4374 1148 4378 1152
rect 4398 1148 4402 1152
rect 4406 1148 4410 1152
rect 4446 1148 4450 1152
rect 4494 1148 4498 1152
rect 4510 1148 4514 1152
rect 4518 1148 4522 1152
rect 4534 1148 4538 1152
rect 4590 1148 4594 1152
rect 4598 1148 4602 1152
rect 4638 1148 4642 1152
rect 4646 1148 4650 1152
rect 4654 1148 4658 1152
rect 4678 1148 4682 1152
rect 4710 1148 4714 1152
rect 4798 1148 4802 1152
rect 4854 1148 4858 1152
rect 4886 1148 4890 1152
rect 2350 1138 2354 1142
rect 2382 1138 2386 1142
rect 2414 1138 2418 1142
rect 2446 1138 2450 1142
rect 2550 1138 2554 1142
rect 2606 1138 2610 1142
rect 2654 1138 2658 1142
rect 2702 1138 2706 1142
rect 2790 1138 2794 1142
rect 2902 1138 2906 1142
rect 2942 1138 2946 1142
rect 2998 1138 3002 1142
rect 3102 1138 3106 1142
rect 3150 1138 3154 1142
rect 3230 1138 3234 1142
rect 3478 1138 3482 1142
rect 3494 1138 3498 1142
rect 3550 1138 3554 1142
rect 3598 1138 3602 1142
rect 3662 1138 3666 1142
rect 3742 1138 3746 1142
rect 3750 1138 3754 1142
rect 3782 1138 3786 1142
rect 3902 1138 3906 1142
rect 3934 1138 3938 1142
rect 4006 1138 4010 1142
rect 4038 1138 4042 1142
rect 4102 1138 4106 1142
rect 4126 1138 4130 1142
rect 4222 1138 4226 1142
rect 4326 1138 4330 1142
rect 4358 1138 4362 1142
rect 4422 1138 4426 1142
rect 4486 1138 4490 1142
rect 4518 1138 4522 1142
rect 4926 1148 4930 1152
rect 4974 1148 4978 1152
rect 4982 1148 4986 1152
rect 4990 1148 4994 1152
rect 5006 1148 5010 1152
rect 5086 1148 5090 1152
rect 4606 1138 4610 1142
rect 4702 1138 4706 1142
rect 4822 1138 4826 1142
rect 4878 1138 4882 1142
rect 4910 1138 4914 1142
rect 4918 1138 4922 1142
rect 4934 1138 4938 1142
rect 5014 1138 5018 1142
rect 5078 1138 5082 1142
rect 5110 1138 5114 1142
rect 5126 1138 5130 1142
rect 246 1128 250 1132
rect 454 1128 458 1132
rect 502 1128 506 1132
rect 510 1128 514 1132
rect 518 1128 522 1132
rect 934 1128 938 1132
rect 942 1128 946 1132
rect 1110 1128 1114 1132
rect 1286 1128 1290 1132
rect 1358 1128 1362 1132
rect 1374 1128 1378 1132
rect 1398 1128 1402 1132
rect 1654 1128 1658 1132
rect 1830 1128 1834 1132
rect 1862 1128 1866 1132
rect 2038 1128 2042 1132
rect 2246 1128 2250 1132
rect 2406 1128 2410 1132
rect 2742 1128 2746 1132
rect 2750 1128 2754 1132
rect 2982 1128 2986 1132
rect 3046 1128 3050 1132
rect 3166 1128 3170 1132
rect 3326 1128 3330 1132
rect 3558 1128 3562 1132
rect 3710 1128 3714 1132
rect 4166 1128 4170 1132
rect 4310 1128 4314 1132
rect 4462 1128 4466 1132
rect 4542 1128 4546 1132
rect 4838 1128 4842 1132
rect 4894 1128 4898 1132
rect 4958 1128 4962 1132
rect 62 1118 66 1122
rect 342 1118 346 1122
rect 486 1118 490 1122
rect 574 1118 578 1122
rect 630 1118 634 1122
rect 806 1118 810 1122
rect 910 1118 914 1122
rect 1094 1118 1098 1122
rect 1134 1118 1138 1122
rect 1350 1118 1354 1122
rect 1382 1118 1386 1122
rect 1910 1118 1914 1122
rect 2286 1118 2290 1122
rect 2462 1118 2466 1122
rect 2574 1118 2578 1122
rect 2622 1118 2626 1122
rect 2806 1118 2810 1122
rect 3126 1118 3130 1122
rect 4054 1118 4058 1122
rect 4350 1118 4354 1122
rect 4430 1118 4434 1122
rect 4478 1118 4482 1122
rect 4726 1118 4730 1122
rect 4902 1118 4906 1122
rect 4942 1118 4946 1122
rect 1050 1103 1054 1107
rect 1057 1103 1061 1107
rect 2074 1103 2078 1107
rect 2081 1103 2085 1107
rect 3098 1103 3102 1107
rect 3105 1103 3109 1107
rect 4114 1103 4118 1107
rect 4121 1103 4125 1107
rect 94 1088 98 1092
rect 670 1088 674 1092
rect 854 1088 858 1092
rect 870 1088 874 1092
rect 902 1088 906 1092
rect 998 1088 1002 1092
rect 1014 1088 1018 1092
rect 1030 1088 1034 1092
rect 1294 1088 1298 1092
rect 1406 1088 1410 1092
rect 1454 1088 1458 1092
rect 1470 1088 1474 1092
rect 1862 1088 1866 1092
rect 1998 1088 2002 1092
rect 2062 1088 2066 1092
rect 2214 1088 2218 1092
rect 2222 1088 2226 1092
rect 2398 1088 2402 1092
rect 2430 1088 2434 1092
rect 2606 1088 2610 1092
rect 2718 1088 2722 1092
rect 2734 1088 2738 1092
rect 2990 1088 2994 1092
rect 3254 1088 3258 1092
rect 3462 1088 3466 1092
rect 3622 1088 3626 1092
rect 3726 1088 3730 1092
rect 3838 1088 3842 1092
rect 3862 1088 3866 1092
rect 3886 1088 3890 1092
rect 3998 1088 4002 1092
rect 4190 1088 4194 1092
rect 4246 1088 4250 1092
rect 4310 1088 4314 1092
rect 4470 1088 4474 1092
rect 4574 1088 4578 1092
rect 4662 1088 4666 1092
rect 4830 1088 4834 1092
rect 4870 1088 4874 1092
rect 4886 1088 4890 1092
rect 5014 1088 5018 1092
rect 166 1078 170 1082
rect 214 1078 218 1082
rect 270 1078 274 1082
rect 462 1078 466 1082
rect 774 1078 778 1082
rect 806 1078 810 1082
rect 862 1078 866 1082
rect 1342 1078 1346 1082
rect 1414 1078 1418 1082
rect 1830 1078 1834 1082
rect 2470 1078 2474 1082
rect 2542 1078 2546 1082
rect 2878 1078 2882 1082
rect 3302 1078 3306 1082
rect 3622 1078 3626 1082
rect 3710 1078 3714 1082
rect 126 1068 130 1072
rect 158 1068 162 1072
rect 174 1068 178 1072
rect 206 1068 210 1072
rect 238 1068 242 1072
rect 342 1068 346 1072
rect 374 1068 378 1072
rect 406 1068 410 1072
rect 430 1068 434 1072
rect 574 1068 578 1072
rect 590 1068 594 1072
rect 606 1068 610 1072
rect 686 1068 690 1072
rect 814 1068 818 1072
rect 830 1068 834 1072
rect 878 1068 882 1072
rect 918 1068 922 1072
rect 1022 1068 1026 1072
rect 1046 1068 1050 1072
rect 1070 1068 1074 1072
rect 1094 1068 1098 1072
rect 1134 1068 1138 1072
rect 1190 1068 1194 1072
rect 1310 1068 1314 1072
rect 1326 1068 1330 1072
rect 1430 1068 1434 1072
rect 1446 1068 1450 1072
rect 1526 1068 1530 1072
rect 1606 1068 1610 1072
rect 38 1058 42 1062
rect 62 1058 66 1062
rect 102 1058 106 1062
rect 118 1058 122 1062
rect 134 1058 138 1062
rect 150 1058 154 1062
rect 182 1058 186 1062
rect 198 1058 202 1062
rect 238 1058 242 1062
rect 278 1058 282 1062
rect 350 1058 354 1062
rect 374 1058 378 1062
rect 414 1058 418 1062
rect 462 1059 466 1063
rect 534 1058 538 1062
rect 566 1058 570 1062
rect 614 1058 618 1062
rect 710 1058 714 1062
rect 726 1058 730 1062
rect 790 1058 794 1062
rect 822 1058 826 1062
rect 838 1058 842 1062
rect 886 1058 890 1062
rect 942 1058 946 1062
rect 1070 1058 1074 1062
rect 1118 1058 1122 1062
rect 1158 1058 1162 1062
rect 1190 1058 1194 1062
rect 1222 1059 1226 1063
rect 1254 1058 1258 1062
rect 1350 1058 1354 1062
rect 1438 1058 1442 1062
rect 1502 1058 1506 1062
rect 1534 1059 1538 1063
rect 1638 1068 1642 1072
rect 1646 1068 1650 1072
rect 1662 1068 1666 1072
rect 1678 1068 1682 1072
rect 1822 1068 1826 1072
rect 1862 1068 1866 1072
rect 1878 1068 1882 1072
rect 1902 1068 1906 1072
rect 1910 1068 1914 1072
rect 1950 1068 1954 1072
rect 2022 1068 2026 1072
rect 2070 1068 2074 1072
rect 2118 1068 2122 1072
rect 2158 1068 2162 1072
rect 2238 1068 2242 1072
rect 2246 1068 2250 1072
rect 2302 1068 2306 1072
rect 2318 1068 2322 1072
rect 2406 1068 2410 1072
rect 2438 1068 2442 1072
rect 2630 1068 2634 1072
rect 2702 1068 2706 1072
rect 2726 1068 2730 1072
rect 2774 1068 2778 1072
rect 2830 1068 2834 1072
rect 2854 1068 2858 1072
rect 3110 1068 3114 1072
rect 3190 1068 3194 1072
rect 3222 1068 3226 1072
rect 3262 1068 3266 1072
rect 3366 1068 3370 1072
rect 3382 1068 3386 1072
rect 3406 1068 3410 1072
rect 3422 1068 3426 1072
rect 3438 1068 3442 1072
rect 3486 1068 3490 1072
rect 3502 1068 3506 1072
rect 3534 1068 3538 1072
rect 3590 1068 3594 1072
rect 3670 1068 3674 1072
rect 3734 1068 3738 1072
rect 3758 1068 3762 1072
rect 3846 1068 3850 1072
rect 3934 1068 3938 1072
rect 3990 1068 3994 1072
rect 4030 1068 4034 1072
rect 4070 1068 4074 1072
rect 4174 1068 4178 1072
rect 4214 1068 4218 1072
rect 1598 1058 1602 1062
rect 1614 1058 1618 1062
rect 1646 1058 1650 1062
rect 1654 1058 1658 1062
rect 1734 1058 1738 1062
rect 1766 1059 1770 1063
rect 1830 1058 1834 1062
rect 1854 1058 1858 1062
rect 1918 1058 1922 1062
rect 1974 1058 1978 1062
rect 1982 1058 1986 1062
rect 2014 1058 2018 1062
rect 2030 1058 2034 1062
rect 2118 1058 2122 1062
rect 2150 1059 2154 1063
rect 2254 1058 2258 1062
rect 2278 1058 2282 1062
rect 2294 1058 2298 1062
rect 2334 1059 2338 1063
rect 2406 1058 2410 1062
rect 2430 1058 2434 1062
rect 2494 1058 2498 1062
rect 2550 1058 2554 1062
rect 2566 1058 2570 1062
rect 2590 1058 2594 1062
rect 2614 1058 2618 1062
rect 2622 1058 2626 1062
rect 2630 1058 2634 1062
rect 2662 1058 2666 1062
rect 2670 1058 2674 1062
rect 2678 1058 2682 1062
rect 2694 1058 2698 1062
rect 2766 1058 2770 1062
rect 2790 1058 2794 1062
rect 2830 1058 2834 1062
rect 2862 1058 2866 1062
rect 2926 1058 2930 1062
rect 2942 1058 2946 1062
rect 3006 1058 3010 1062
rect 3038 1058 3042 1062
rect 3070 1058 3074 1062
rect 3078 1058 3082 1062
rect 3150 1058 3154 1062
rect 3238 1058 3242 1062
rect 3350 1059 3354 1063
rect 3398 1058 3402 1062
rect 3430 1058 3434 1062
rect 3438 1058 3442 1062
rect 3526 1058 3530 1062
rect 3542 1058 3546 1062
rect 3598 1058 3602 1062
rect 3638 1058 3642 1062
rect 3694 1058 3698 1062
rect 3742 1058 3746 1062
rect 3774 1059 3778 1063
rect 4254 1068 4258 1072
rect 4326 1068 4330 1072
rect 4366 1068 4370 1072
rect 4454 1068 4458 1072
rect 4526 1068 4530 1072
rect 4566 1068 4570 1072
rect 4598 1068 4602 1072
rect 4622 1078 4626 1082
rect 4862 1078 4866 1082
rect 5046 1078 5050 1082
rect 5078 1078 5082 1082
rect 4790 1068 4794 1072
rect 4966 1068 4970 1072
rect 5006 1068 5010 1072
rect 5110 1068 5114 1072
rect 5174 1068 5178 1072
rect 3862 1058 3866 1062
rect 3878 1058 3882 1062
rect 3902 1058 3906 1062
rect 3966 1058 3970 1062
rect 4014 1058 4018 1062
rect 4022 1058 4026 1062
rect 4054 1058 4058 1062
rect 4142 1058 4146 1062
rect 4206 1058 4210 1062
rect 4222 1058 4226 1062
rect 4230 1058 4234 1062
rect 4334 1058 4338 1062
rect 4342 1058 4346 1062
rect 4422 1058 4426 1062
rect 4518 1058 4522 1062
rect 4582 1058 4586 1062
rect 4638 1058 4642 1062
rect 4694 1058 4698 1062
rect 4718 1058 4722 1062
rect 4758 1058 4762 1062
rect 4814 1058 4818 1062
rect 4822 1058 4826 1062
rect 4846 1058 4850 1062
rect 4878 1058 4882 1062
rect 4942 1058 4946 1062
rect 4982 1058 4986 1062
rect 4998 1058 5002 1062
rect 5054 1058 5058 1062
rect 102 1048 106 1052
rect 214 1048 218 1052
rect 366 1048 370 1052
rect 398 1048 402 1052
rect 430 1048 434 1052
rect 542 1048 546 1052
rect 854 1048 858 1052
rect 902 1048 906 1052
rect 1006 1048 1010 1052
rect 1022 1048 1026 1052
rect 1102 1048 1106 1052
rect 1166 1048 1170 1052
rect 1294 1048 1298 1052
rect 1414 1048 1418 1052
rect 1462 1048 1466 1052
rect 1566 1048 1570 1052
rect 1598 1048 1602 1052
rect 1614 1048 1618 1052
rect 1814 1048 1818 1052
rect 1830 1048 1834 1052
rect 1862 1048 1866 1052
rect 1878 1048 1882 1052
rect 1934 1048 1938 1052
rect 2030 1048 2034 1052
rect 2046 1048 2050 1052
rect 2054 1048 2058 1052
rect 2094 1048 2098 1052
rect 2110 1048 2114 1052
rect 2222 1048 2226 1052
rect 2254 1048 2258 1052
rect 2270 1048 2274 1052
rect 2278 1048 2282 1052
rect 2430 1048 2434 1052
rect 2446 1048 2450 1052
rect 2470 1048 2474 1052
rect 2510 1048 2514 1052
rect 2678 1048 2682 1052
rect 2710 1048 2714 1052
rect 3614 1048 3618 1052
rect 3646 1048 3650 1052
rect 3662 1048 3666 1052
rect 3918 1048 3922 1052
rect 4054 1048 4058 1052
rect 4190 1048 4194 1052
rect 4246 1048 4250 1052
rect 4350 1048 4354 1052
rect 4582 1048 4586 1052
rect 4614 1048 4618 1052
rect 4806 1048 4810 1052
rect 4982 1048 4986 1052
rect 134 1038 138 1042
rect 198 1038 202 1042
rect 334 1038 338 1042
rect 350 1038 354 1042
rect 382 1038 386 1042
rect 1142 1038 1146 1042
rect 1182 1038 1186 1042
rect 1286 1038 1290 1042
rect 1702 1038 1706 1042
rect 1798 1038 1802 1042
rect 1902 1038 1906 1042
rect 3198 1038 3202 1042
rect 3470 1038 3474 1042
rect 3582 1038 3586 1042
rect 3686 1038 3690 1042
rect 3862 1038 3866 1042
rect 3974 1038 3978 1042
rect 3022 1018 3026 1022
rect 3054 1018 3058 1022
rect 3094 1018 3098 1022
rect 3174 1018 3178 1022
rect 3678 1018 3682 1022
rect 3926 1018 3930 1022
rect 3950 1018 3954 1022
rect 4774 1018 4778 1022
rect 4798 1018 4802 1022
rect 5118 1018 5122 1022
rect 538 1003 542 1007
rect 545 1003 549 1007
rect 1562 1003 1566 1007
rect 1569 1003 1573 1007
rect 2586 1003 2590 1007
rect 2593 1003 2597 1007
rect 3610 1003 3614 1007
rect 3617 1003 3621 1007
rect 4634 1003 4638 1007
rect 4641 1003 4645 1007
rect 94 988 98 992
rect 190 988 194 992
rect 262 988 266 992
rect 366 988 370 992
rect 782 988 786 992
rect 806 988 810 992
rect 966 988 970 992
rect 1110 988 1114 992
rect 1206 988 1210 992
rect 1222 988 1226 992
rect 1358 988 1362 992
rect 1406 988 1410 992
rect 1510 988 1514 992
rect 1614 988 1618 992
rect 1718 988 1722 992
rect 1774 988 1778 992
rect 1862 988 1866 992
rect 2038 988 2042 992
rect 2222 988 2226 992
rect 2246 988 2250 992
rect 2342 988 2346 992
rect 2518 988 2522 992
rect 2542 988 2546 992
rect 2638 988 2642 992
rect 2750 988 2754 992
rect 2942 988 2946 992
rect 2982 988 2986 992
rect 3150 988 3154 992
rect 3398 988 3402 992
rect 3606 988 3610 992
rect 3718 988 3722 992
rect 3734 988 3738 992
rect 3814 988 3818 992
rect 3998 988 4002 992
rect 4414 988 4418 992
rect 4630 988 4634 992
rect 4678 988 4682 992
rect 4982 988 4986 992
rect 2054 978 2058 982
rect 230 968 234 972
rect 390 968 394 972
rect 502 968 506 972
rect 838 968 842 972
rect 1126 968 1130 972
rect 1150 968 1154 972
rect 1558 968 1562 972
rect 1622 968 1626 972
rect 1982 968 1986 972
rect 2838 968 2842 972
rect 3254 968 3258 972
rect 3830 968 3834 972
rect 4094 968 4098 972
rect 4878 968 4882 972
rect 206 958 210 962
rect 46 948 50 952
rect 134 948 138 952
rect 206 948 210 952
rect 246 948 250 952
rect 318 948 322 952
rect 366 948 370 952
rect 470 958 474 962
rect 510 958 514 962
rect 646 958 650 962
rect 406 948 410 952
rect 438 948 442 952
rect 454 948 458 952
rect 486 948 490 952
rect 502 948 506 952
rect 614 947 618 951
rect 662 948 666 952
rect 694 948 698 952
rect 718 948 722 952
rect 822 948 826 952
rect 974 958 978 962
rect 854 948 858 952
rect 862 948 866 952
rect 14 938 18 942
rect 110 938 114 942
rect 198 938 202 942
rect 254 938 258 942
rect 326 938 330 942
rect 358 938 362 942
rect 414 938 418 942
rect 446 938 450 942
rect 478 938 482 942
rect 526 938 530 942
rect 606 938 610 942
rect 646 938 650 942
rect 670 938 674 942
rect 902 947 906 951
rect 982 948 986 952
rect 1006 948 1010 952
rect 1062 948 1066 952
rect 1126 948 1130 952
rect 1262 958 1266 962
rect 1398 958 1402 962
rect 1438 958 1442 962
rect 1502 958 1506 962
rect 1518 958 1522 962
rect 1166 948 1170 952
rect 1246 948 1250 952
rect 1262 948 1266 952
rect 1294 947 1298 951
rect 1366 948 1370 952
rect 1382 948 1386 952
rect 1446 948 1450 952
rect 1534 948 1538 952
rect 1590 958 1594 962
rect 1790 958 1794 962
rect 1822 958 1826 962
rect 1838 958 1842 962
rect 1590 948 1594 952
rect 1678 948 1682 952
rect 1758 948 1762 952
rect 1774 948 1778 952
rect 1806 948 1810 952
rect 1822 948 1826 952
rect 1838 948 1842 952
rect 1918 948 1922 952
rect 1966 948 1970 952
rect 2006 958 2010 962
rect 2150 958 2154 962
rect 2166 958 2170 962
rect 2182 958 2186 962
rect 2238 958 2242 962
rect 2510 958 2514 962
rect 3014 958 3018 962
rect 2022 948 2026 952
rect 2110 948 2114 952
rect 2166 948 2170 952
rect 2198 948 2202 952
rect 2222 948 2226 952
rect 2294 948 2298 952
rect 2350 948 2354 952
rect 702 938 706 942
rect 726 938 730 942
rect 814 938 818 942
rect 870 938 874 942
rect 918 938 922 942
rect 998 938 1002 942
rect 1030 938 1034 942
rect 1118 938 1122 942
rect 1174 938 1178 942
rect 1214 938 1218 942
rect 1238 938 1242 942
rect 1278 938 1282 942
rect 1390 938 1394 942
rect 1422 938 1426 942
rect 1478 938 1482 942
rect 1494 938 1498 942
rect 1502 938 1506 942
rect 1526 938 1530 942
rect 1598 938 1602 942
rect 1702 938 1706 942
rect 1766 938 1770 942
rect 1798 938 1802 942
rect 1830 938 1834 942
rect 1918 938 1922 942
rect 1942 938 1946 942
rect 1958 938 1962 942
rect 2014 938 2018 942
rect 2134 938 2138 942
rect 2174 938 2178 942
rect 2206 938 2210 942
rect 2214 938 2218 942
rect 2278 938 2282 942
rect 2326 938 2330 942
rect 2382 947 2386 951
rect 2454 948 2458 952
rect 2486 948 2490 952
rect 2558 948 2562 952
rect 2566 948 2570 952
rect 2614 948 2618 952
rect 2622 948 2626 952
rect 2646 948 2650 952
rect 2662 948 2666 952
rect 2798 948 2802 952
rect 2862 948 2866 952
rect 2918 948 2922 952
rect 2926 948 2930 952
rect 2950 948 2954 952
rect 2958 948 2962 952
rect 2966 948 2970 952
rect 2974 948 2978 952
rect 2998 948 3002 952
rect 3070 948 3074 952
rect 3198 948 3202 952
rect 3262 948 3266 952
rect 3278 948 3282 952
rect 3294 958 3298 962
rect 3366 958 3370 962
rect 3478 958 3482 962
rect 3310 948 3314 952
rect 3350 948 3354 952
rect 3406 948 3410 952
rect 3414 948 3418 952
rect 3422 948 3426 952
rect 3462 948 3466 952
rect 3750 958 3754 962
rect 3798 958 3802 962
rect 3942 958 3946 962
rect 3982 958 3986 962
rect 4014 958 4018 962
rect 3494 948 3498 952
rect 3502 948 3506 952
rect 3550 948 3554 952
rect 3662 948 3666 952
rect 3726 948 3730 952
rect 3782 948 3786 952
rect 3798 948 3802 952
rect 3822 948 3826 952
rect 3886 948 3890 952
rect 3974 948 3978 952
rect 4006 948 4010 952
rect 4054 948 4058 952
rect 4070 948 4074 952
rect 4086 948 4090 952
rect 4166 948 4170 952
rect 4214 948 4218 952
rect 2462 938 2466 942
rect 2534 938 2538 942
rect 2686 938 2690 942
rect 2806 938 2810 942
rect 2870 938 2874 942
rect 3030 938 3034 942
rect 62 928 66 932
rect 422 928 426 932
rect 678 928 682 932
rect 798 928 802 932
rect 1230 928 1234 932
rect 1294 928 1298 932
rect 1606 928 1610 932
rect 1726 928 1730 932
rect 2022 928 2026 932
rect 2350 928 2354 932
rect 2382 928 2386 932
rect 2502 928 2506 932
rect 2878 928 2882 932
rect 3158 938 3162 942
rect 3174 938 3178 942
rect 3198 938 3202 942
rect 3262 938 3266 942
rect 3318 938 3322 942
rect 3454 938 3458 942
rect 3510 938 3514 942
rect 3550 938 3554 942
rect 3638 938 3642 942
rect 3686 938 3690 942
rect 3726 938 3730 942
rect 3774 938 3778 942
rect 3886 938 3890 942
rect 3926 938 3930 942
rect 4014 938 4018 942
rect 4030 938 4034 942
rect 4078 938 4082 942
rect 4190 938 4194 942
rect 4286 947 4290 951
rect 4326 948 4330 952
rect 4334 948 4338 952
rect 4350 958 4354 962
rect 4390 958 4394 962
rect 4398 958 4402 962
rect 4470 958 4474 962
rect 4734 958 4738 962
rect 4742 958 4746 962
rect 4758 958 4762 962
rect 4886 958 4890 962
rect 4998 958 5002 962
rect 5182 958 5186 962
rect 4414 948 4418 952
rect 4454 948 4458 952
rect 4470 948 4474 952
rect 4518 948 4522 952
rect 4670 948 4674 952
rect 4694 948 4698 952
rect 4702 948 4706 952
rect 4718 948 4722 952
rect 4734 948 4738 952
rect 4758 948 4762 952
rect 4814 947 4818 951
rect 4886 948 4890 952
rect 4902 948 4906 952
rect 4918 948 4922 952
rect 4950 948 4954 952
rect 4966 948 4970 952
rect 4974 948 4978 952
rect 4302 938 4306 942
rect 4318 938 4322 942
rect 4366 938 4370 942
rect 4374 938 4378 942
rect 4526 938 4530 942
rect 4558 938 4562 942
rect 4574 938 4578 942
rect 4710 938 4714 942
rect 4766 938 4770 942
rect 5102 947 5106 951
rect 5134 948 5138 952
rect 5142 948 5146 952
rect 5158 948 5162 952
rect 4910 938 4914 942
rect 4926 938 4930 942
rect 4990 938 4994 942
rect 5014 938 5018 942
rect 5030 938 5034 942
rect 5118 938 5122 942
rect 5166 938 5170 942
rect 2894 928 2898 932
rect 3062 928 3066 932
rect 3094 928 3098 932
rect 3326 928 3330 932
rect 3766 928 3770 932
rect 3806 928 3810 932
rect 4014 928 4018 932
rect 4038 928 4042 932
rect 4438 928 4442 932
rect 4782 928 4786 932
rect 4814 928 4818 932
rect 4966 928 4970 932
rect 430 918 434 922
rect 470 918 474 922
rect 518 918 522 922
rect 550 918 554 922
rect 1206 918 1210 922
rect 1430 918 1434 922
rect 1462 918 1466 922
rect 1742 918 1746 922
rect 2182 918 2186 922
rect 2246 918 2250 922
rect 2446 918 2450 922
rect 2470 918 2474 922
rect 2582 918 2586 922
rect 2854 918 2858 922
rect 3022 918 3026 922
rect 3134 918 3138 922
rect 3718 918 3722 922
rect 3942 918 3946 922
rect 3958 918 3962 922
rect 4390 918 4394 922
rect 4478 918 4482 922
rect 4934 918 4938 922
rect 5006 918 5010 922
rect 1050 903 1054 907
rect 1057 903 1061 907
rect 2074 903 2078 907
rect 2081 903 2085 907
rect 3098 903 3102 907
rect 3105 903 3109 907
rect 4114 903 4118 907
rect 4121 903 4125 907
rect 94 888 98 892
rect 254 888 258 892
rect 438 888 442 892
rect 534 888 538 892
rect 566 888 570 892
rect 758 888 762 892
rect 790 888 794 892
rect 878 888 882 892
rect 894 888 898 892
rect 918 888 922 892
rect 974 888 978 892
rect 990 888 994 892
rect 1126 888 1130 892
rect 1222 888 1226 892
rect 1254 888 1258 892
rect 1374 888 1378 892
rect 1534 888 1538 892
rect 1630 888 1634 892
rect 1654 888 1658 892
rect 1678 888 1682 892
rect 1806 888 1810 892
rect 1910 888 1914 892
rect 2110 888 2114 892
rect 2142 888 2146 892
rect 2238 888 2242 892
rect 2294 888 2298 892
rect 2334 888 2338 892
rect 2382 888 2386 892
rect 2534 888 2538 892
rect 2614 888 2618 892
rect 2702 888 2706 892
rect 2886 888 2890 892
rect 2998 888 3002 892
rect 3094 888 3098 892
rect 3206 888 3210 892
rect 3318 888 3322 892
rect 3750 888 3754 892
rect 3798 888 3802 892
rect 3814 888 3818 892
rect 3918 888 3922 892
rect 3998 888 4002 892
rect 4134 888 4138 892
rect 4238 888 4242 892
rect 4262 888 4266 892
rect 4278 888 4282 892
rect 4310 888 4314 892
rect 4478 888 4482 892
rect 4542 888 4546 892
rect 4766 888 4770 892
rect 4870 888 4874 892
rect 4974 888 4978 892
rect 5126 888 5130 892
rect 342 878 346 882
rect 550 878 554 882
rect 1422 878 1426 882
rect 2262 878 2266 882
rect 2366 878 2370 882
rect 2646 878 2650 882
rect 2958 878 2962 882
rect 3246 878 3250 882
rect 3406 878 3410 882
rect 3494 878 3498 882
rect 3670 878 3674 882
rect 3718 878 3722 882
rect 3974 878 3978 882
rect 4078 878 4082 882
rect 4374 878 4378 882
rect 4454 878 4458 882
rect 4574 878 4578 882
rect 4726 878 4730 882
rect 14 868 18 872
rect 102 868 106 872
rect 158 868 162 872
rect 174 868 178 872
rect 286 868 290 872
rect 302 868 306 872
rect 318 868 322 872
rect 374 868 378 872
rect 478 868 482 872
rect 598 868 602 872
rect 606 868 610 872
rect 662 868 666 872
rect 678 868 682 872
rect 766 868 770 872
rect 822 868 826 872
rect 830 868 834 872
rect 838 868 842 872
rect 870 868 874 872
rect 910 868 914 872
rect 934 868 938 872
rect 982 868 986 872
rect 1014 868 1018 872
rect 1030 868 1034 872
rect 1134 868 1138 872
rect 1150 868 1154 872
rect 1198 868 1202 872
rect 1214 868 1218 872
rect 1246 868 1250 872
rect 1294 868 1298 872
rect 1334 868 1338 872
rect 1350 868 1354 872
rect 1406 868 1410 872
rect 1454 868 1458 872
rect 1486 868 1490 872
rect 1542 868 1546 872
rect 1574 868 1578 872
rect 1614 868 1618 872
rect 1622 868 1626 872
rect 1646 868 1650 872
rect 1702 868 1706 872
rect 1758 868 1762 872
rect 1766 868 1770 872
rect 1782 868 1786 872
rect 1798 868 1802 872
rect 1822 868 1826 872
rect 1918 868 1922 872
rect 2022 868 2026 872
rect 2038 868 2042 872
rect 2078 868 2082 872
rect 2134 868 2138 872
rect 2222 868 2226 872
rect 2254 868 2258 872
rect 2302 868 2306 872
rect 2438 868 2442 872
rect 2454 868 2458 872
rect 2574 868 2578 872
rect 2638 868 2642 872
rect 2686 868 2690 872
rect 2806 868 2810 872
rect 2894 868 2898 872
rect 2910 868 2914 872
rect 2950 868 2954 872
rect 3014 868 3018 872
rect 3062 868 3066 872
rect 3118 868 3122 872
rect 3174 868 3178 872
rect 3182 868 3186 872
rect 3238 868 3242 872
rect 3286 868 3290 872
rect 3342 868 3346 872
rect 3374 868 3378 872
rect 3406 868 3410 872
rect 3470 868 3474 872
rect 3542 868 3546 872
rect 3582 868 3586 872
rect 3614 868 3618 872
rect 3686 868 3690 872
rect 3758 868 3762 872
rect 3774 868 3778 872
rect 3806 868 3810 872
rect 3838 868 3842 872
rect 3886 868 3890 872
rect 3934 868 3938 872
rect 3950 868 3954 872
rect 4030 868 4034 872
rect 4214 868 4218 872
rect 4230 868 4234 872
rect 4246 868 4250 872
rect 4302 868 4306 872
rect 4414 868 4418 872
rect 4462 868 4466 872
rect 4526 868 4530 872
rect 4606 868 4610 872
rect 4622 868 4626 872
rect 4638 868 4642 872
rect 4678 868 4682 872
rect 4702 868 4706 872
rect 4830 878 4834 882
rect 4750 868 4754 872
rect 4862 868 4866 872
rect 4894 868 4898 872
rect 4982 868 4986 872
rect 5022 868 5026 872
rect 5094 868 5098 872
rect 5158 868 5162 872
rect 38 858 42 862
rect 110 858 114 862
rect 118 858 122 862
rect 150 858 154 862
rect 206 858 210 862
rect 286 858 290 862
rect 294 858 298 862
rect 326 858 330 862
rect 382 858 386 862
rect 398 858 402 862
rect 470 859 474 863
rect 590 858 594 862
rect 614 858 618 862
rect 646 858 650 862
rect 654 858 658 862
rect 694 859 698 863
rect 774 858 778 862
rect 1006 858 1010 862
rect 1070 858 1074 862
rect 1142 858 1146 862
rect 1182 858 1186 862
rect 1238 858 1242 862
rect 1318 859 1322 863
rect 1358 858 1362 862
rect 1398 858 1402 862
rect 1438 858 1442 862
rect 1478 858 1482 862
rect 1550 858 1554 862
rect 1606 858 1610 862
rect 1694 858 1698 862
rect 1710 858 1714 862
rect 1750 858 1754 862
rect 1774 858 1778 862
rect 1894 858 1898 862
rect 1958 858 1962 862
rect 1974 858 1978 862
rect 2030 858 2034 862
rect 2070 858 2074 862
rect 2182 858 2186 862
rect 2278 858 2282 862
rect 2310 858 2314 862
rect 2318 858 2322 862
rect 2350 858 2354 862
rect 2470 859 2474 863
rect 2566 858 2570 862
rect 2630 858 2634 862
rect 2662 858 2666 862
rect 2694 858 2698 862
rect 2758 858 2762 862
rect 2830 858 2834 862
rect 2846 858 2850 862
rect 2902 858 2906 862
rect 2942 858 2946 862
rect 2982 858 2986 862
rect 3038 858 3042 862
rect 3126 858 3130 862
rect 3166 858 3170 862
rect 3190 858 3194 862
rect 3230 858 3234 862
rect 3270 858 3274 862
rect 3294 858 3298 862
rect 3302 858 3306 862
rect 3326 858 3330 862
rect 3382 858 3386 862
rect 3422 858 3426 862
rect 3462 858 3466 862
rect 3478 858 3482 862
rect 3558 858 3562 862
rect 3710 858 3714 862
rect 3734 858 3738 862
rect 3766 858 3770 862
rect 3782 858 3786 862
rect 3870 858 3874 862
rect 3926 858 3930 862
rect 3958 858 3962 862
rect 3982 858 3986 862
rect 4054 858 4058 862
rect 4086 858 4090 862
rect 4118 858 4122 862
rect 4190 858 4194 862
rect 4294 858 4298 862
rect 4374 859 4378 863
rect 4406 858 4410 862
rect 4422 858 4426 862
rect 4438 858 4442 862
rect 4486 858 4490 862
rect 4494 858 4498 862
rect 4526 858 4530 862
rect 4558 858 4562 862
rect 4566 858 4570 862
rect 4590 858 4594 862
rect 4614 858 4618 862
rect 4662 858 4666 862
rect 4710 858 4714 862
rect 4742 858 4746 862
rect 4758 858 4762 862
rect 4822 858 4826 862
rect 4934 858 4938 862
rect 4990 858 4994 862
rect 5078 858 5082 862
rect 5142 858 5146 862
rect 5166 858 5170 862
rect 5174 858 5178 862
rect 134 848 138 852
rect 574 848 578 852
rect 630 848 634 852
rect 790 848 794 852
rect 798 848 802 852
rect 886 848 890 852
rect 894 848 898 852
rect 918 848 922 852
rect 958 848 962 852
rect 966 848 970 852
rect 982 848 986 852
rect 1166 848 1170 852
rect 1198 848 1202 852
rect 1382 848 1386 852
rect 1566 848 1570 852
rect 1638 848 1642 852
rect 1662 848 1666 852
rect 1734 848 1738 852
rect 1798 848 1802 852
rect 1814 848 1818 852
rect 2238 848 2242 852
rect 2598 848 2602 852
rect 2926 848 2930 852
rect 2998 848 3002 852
rect 3126 848 3130 852
rect 3150 848 3154 852
rect 3214 848 3218 852
rect 3286 848 3290 852
rect 3446 848 3450 852
rect 3798 848 3802 852
rect 3822 848 3826 852
rect 4014 848 4018 852
rect 4110 848 4114 852
rect 4254 848 4258 852
rect 4270 848 4274 852
rect 4278 848 4282 852
rect 4478 848 4482 852
rect 4630 848 4634 852
rect 4686 848 4690 852
rect 4878 848 4882 852
rect 4990 848 4994 852
rect 5006 848 5010 852
rect 5126 848 5130 852
rect 5182 848 5186 852
rect 518 838 522 842
rect 870 838 874 842
rect 942 838 946 842
rect 2014 838 2018 842
rect 2054 838 2058 842
rect 2518 838 2522 842
rect 2670 838 2674 842
rect 3358 838 3362 842
rect 3422 838 3426 842
rect 3502 838 3506 842
rect 4550 838 4554 842
rect 278 818 282 822
rect 590 818 594 822
rect 806 818 810 822
rect 846 818 850 822
rect 1654 818 1658 822
rect 1710 818 1714 822
rect 1878 818 1882 822
rect 2550 818 2554 822
rect 3486 818 3490 822
rect 3998 818 4002 822
rect 4054 818 4058 822
rect 4502 818 4506 822
rect 538 803 542 807
rect 545 803 549 807
rect 1562 803 1566 807
rect 1569 803 1573 807
rect 2586 803 2590 807
rect 2593 803 2597 807
rect 3610 803 3614 807
rect 3617 803 3621 807
rect 4634 803 4638 807
rect 4641 803 4645 807
rect 182 788 186 792
rect 350 788 354 792
rect 694 788 698 792
rect 710 788 714 792
rect 742 788 746 792
rect 766 788 770 792
rect 942 788 946 792
rect 990 788 994 792
rect 1014 788 1018 792
rect 1078 788 1082 792
rect 1302 788 1306 792
rect 1390 788 1394 792
rect 1526 788 1530 792
rect 1622 788 1626 792
rect 1774 788 1778 792
rect 1782 788 1786 792
rect 1806 788 1810 792
rect 1822 788 1826 792
rect 2006 788 2010 792
rect 2022 788 2026 792
rect 2134 788 2138 792
rect 2286 788 2290 792
rect 2390 788 2394 792
rect 2414 788 2418 792
rect 2454 788 2458 792
rect 2486 788 2490 792
rect 2614 788 2618 792
rect 2694 788 2698 792
rect 2822 788 2826 792
rect 2854 788 2858 792
rect 2894 788 2898 792
rect 3086 788 3090 792
rect 3262 788 3266 792
rect 3438 788 3442 792
rect 3454 788 3458 792
rect 3678 788 3682 792
rect 3742 788 3746 792
rect 3758 788 3762 792
rect 3782 788 3786 792
rect 3822 788 3826 792
rect 3878 788 3882 792
rect 3990 788 3994 792
rect 4030 788 4034 792
rect 4286 788 4290 792
rect 4350 788 4354 792
rect 4526 788 4530 792
rect 4590 788 4594 792
rect 4606 788 4610 792
rect 5054 788 5058 792
rect 5182 788 5186 792
rect 1230 778 1234 782
rect 1710 778 1714 782
rect 238 768 242 772
rect 454 768 458 772
rect 494 768 498 772
rect 566 768 570 772
rect 678 768 682 772
rect 1246 768 1250 772
rect 1294 768 1298 772
rect 1518 768 1522 772
rect 1550 768 1554 772
rect 1614 768 1618 772
rect 1662 768 1666 772
rect 2238 768 2242 772
rect 2342 768 2346 772
rect 2366 768 2370 772
rect 3470 768 3474 772
rect 4278 768 4282 772
rect 4654 768 4658 772
rect 254 758 258 762
rect 470 758 474 762
rect 38 748 42 752
rect 102 748 106 752
rect 134 748 138 752
rect 166 748 170 752
rect 190 748 194 752
rect 198 748 202 752
rect 222 748 226 752
rect 238 748 242 752
rect 254 748 258 752
rect 398 748 402 752
rect 470 748 474 752
rect 526 748 530 752
rect 590 758 594 762
rect 726 758 730 762
rect 734 758 738 762
rect 798 758 802 762
rect 846 758 850 762
rect 950 758 954 762
rect 1022 758 1026 762
rect 590 748 594 752
rect 630 747 634 751
rect 710 748 714 752
rect 774 748 778 752
rect 782 748 786 752
rect 814 748 818 752
rect 830 748 834 752
rect 838 748 842 752
rect 878 747 882 751
rect 974 748 978 752
rect 990 748 994 752
rect 1062 748 1066 752
rect 1070 748 1074 752
rect 1094 748 1098 752
rect 1102 748 1106 752
rect 1262 758 1266 762
rect 1278 758 1282 762
rect 1406 758 1410 762
rect 1438 758 1442 762
rect 1462 758 1466 762
rect 1470 758 1474 762
rect 1590 758 1594 762
rect 1798 758 1802 762
rect 2118 758 2122 762
rect 2270 758 2274 762
rect 1126 748 1130 752
rect 1182 748 1186 752
rect 1246 748 1250 752
rect 1278 748 1282 752
rect 1350 748 1354 752
rect 1366 748 1370 752
rect 1390 748 1394 752
rect 1422 748 1426 752
rect 1430 748 1434 752
rect 1638 748 1642 752
rect 1646 748 1650 752
rect 1670 748 1674 752
rect 1686 748 1690 752
rect 1694 748 1698 752
rect 1718 748 1722 752
rect 1758 748 1762 752
rect 1862 748 1866 752
rect 1942 747 1946 751
rect 1974 748 1978 752
rect 2038 748 2042 752
rect 2070 748 2074 752
rect 2078 748 2082 752
rect 2118 748 2122 752
rect 2166 747 2170 751
rect 2238 748 2242 752
rect 2254 748 2258 752
rect 2286 748 2290 752
rect 2326 748 2330 752
rect 2430 758 2434 762
rect 2598 758 2602 762
rect 2654 758 2658 762
rect 2926 758 2930 762
rect 3014 758 3018 762
rect 2366 748 2370 752
rect 2406 748 2410 752
rect 2414 748 2418 752
rect 2438 748 2442 752
rect 2470 748 2474 752
rect 2478 748 2482 752
rect 2518 748 2522 752
rect 2542 748 2546 752
rect 2614 748 2618 752
rect 2622 748 2626 752
rect 2678 748 2682 752
rect 2726 747 2730 751
rect 2798 748 2802 752
rect 2806 748 2810 752
rect 2830 748 2834 752
rect 2862 748 2866 752
rect 2974 747 2978 751
rect 3014 748 3018 752
rect 3038 758 3042 762
rect 3134 758 3138 762
rect 3158 758 3162 762
rect 3182 758 3186 762
rect 3278 758 3282 762
rect 3310 758 3314 762
rect 3054 748 3058 752
rect 3078 748 3082 752
rect 3102 748 3106 752
rect 3110 748 3114 752
rect 3118 748 3122 752
rect 3206 748 3210 752
rect 3262 748 3266 752
rect 3294 748 3298 752
rect 3350 758 3354 762
rect 3334 748 3338 752
rect 3390 748 3394 752
rect 3406 758 3410 762
rect 3702 758 3706 762
rect 3814 758 3818 762
rect 3854 758 3858 762
rect 3422 748 3426 752
rect 3526 748 3530 752
rect 3654 748 3658 752
rect 3686 748 3690 752
rect 3694 748 3698 752
rect 3702 748 3706 752
rect 3718 748 3722 752
rect 3766 748 3770 752
rect 3774 748 3778 752
rect 3798 748 3802 752
rect 4062 758 4066 762
rect 3878 748 3882 752
rect 3910 748 3914 752
rect 3934 748 3938 752
rect 3950 748 3954 752
rect 3982 748 3986 752
rect 4014 748 4018 752
rect 4022 748 4026 752
rect 4054 748 4058 752
rect 4062 748 4066 752
rect 4086 748 4090 752
rect 4134 747 4138 751
rect 4230 748 4234 752
rect 4254 758 4258 762
rect 4326 758 4330 762
rect 4382 758 4386 762
rect 5062 758 5066 762
rect 4294 748 4298 752
rect 4310 748 4314 752
rect 4366 748 4370 752
rect 4374 748 4378 752
rect 4382 748 4386 752
rect 4398 748 4402 752
rect 14 738 18 742
rect 110 738 114 742
rect 206 738 210 742
rect 230 738 234 742
rect 286 738 290 742
rect 294 738 298 742
rect 398 738 402 742
rect 462 738 466 742
rect 518 738 522 742
rect 598 738 602 742
rect 614 738 618 742
rect 702 738 706 742
rect 750 738 754 742
rect 822 738 826 742
rect 862 738 866 742
rect 950 738 954 742
rect 966 738 970 742
rect 998 738 1002 742
rect 1038 738 1042 742
rect 1134 738 1138 742
rect 1150 738 1154 742
rect 1238 738 1242 742
rect 1270 738 1274 742
rect 1318 738 1322 742
rect 1350 738 1354 742
rect 1414 738 1418 742
rect 1446 738 1450 742
rect 1494 738 1498 742
rect 1534 738 1538 742
rect 1558 738 1562 742
rect 1590 738 1594 742
rect 1630 738 1634 742
rect 1814 738 1818 742
rect 1878 738 1882 742
rect 2094 738 2098 742
rect 2150 738 2154 742
rect 2262 738 2266 742
rect 2318 738 2322 742
rect 2374 738 2378 742
rect 2398 738 2402 742
rect 2590 738 2594 742
rect 2622 738 2626 742
rect 2670 738 2674 742
rect 2710 738 2714 742
rect 2958 738 2962 742
rect 3006 738 3010 742
rect 3070 738 3074 742
rect 3150 738 3154 742
rect 3174 738 3178 742
rect 3198 738 3202 742
rect 3286 738 3290 742
rect 3342 738 3346 742
rect 3366 738 3370 742
rect 3374 738 3378 742
rect 3430 738 3434 742
rect 3550 738 3554 742
rect 3566 738 3570 742
rect 3726 738 3730 742
rect 3830 738 3834 742
rect 3838 738 3842 742
rect 3926 738 3930 742
rect 4102 738 4106 742
rect 4222 738 4226 742
rect 4270 738 4274 742
rect 4294 738 4298 742
rect 4438 747 4442 751
rect 4510 748 4514 752
rect 4518 748 4522 752
rect 4558 748 4562 752
rect 4574 748 4578 752
rect 4582 748 4586 752
rect 4678 748 4682 752
rect 4734 748 4738 752
rect 4758 748 4762 752
rect 4806 748 4810 752
rect 4862 748 4866 752
rect 4926 748 4930 752
rect 4958 748 4962 752
rect 5006 748 5010 752
rect 5022 748 5026 752
rect 5118 748 5122 752
rect 5142 748 5146 752
rect 4406 738 4410 742
rect 4422 738 4426 742
rect 4686 738 4690 742
rect 4790 738 4794 742
rect 4798 738 4802 742
rect 4894 738 4898 742
rect 4950 738 4954 742
rect 4974 738 4978 742
rect 5078 738 5082 742
rect 5094 738 5098 742
rect 118 728 122 732
rect 150 728 154 732
rect 630 728 634 732
rect 758 728 762 732
rect 1006 728 1010 732
rect 1310 728 1314 732
rect 1366 728 1370 732
rect 1518 728 1522 732
rect 1766 728 1770 732
rect 1790 728 1794 732
rect 2126 728 2130 732
rect 2310 728 2314 732
rect 2382 728 2386 732
rect 2646 728 2650 732
rect 2686 728 2690 732
rect 2726 728 2730 732
rect 2846 728 2850 732
rect 3238 728 3242 732
rect 3446 728 3450 732
rect 3462 728 3466 732
rect 3734 728 3738 732
rect 3750 728 3754 732
rect 3910 728 3914 732
rect 3926 728 3930 732
rect 3950 728 3954 732
rect 3974 728 3978 732
rect 4006 728 4010 732
rect 4134 728 4138 732
rect 4214 728 4218 732
rect 4558 728 4562 732
rect 4598 728 4602 732
rect 4758 728 4762 732
rect 4774 728 4778 732
rect 4910 728 4914 732
rect 5038 728 5042 732
rect 5190 728 5194 732
rect 94 718 98 722
rect 214 718 218 722
rect 1022 718 1026 722
rect 1110 718 1114 722
rect 1454 718 1458 722
rect 1478 718 1482 722
rect 1502 718 1506 722
rect 1550 718 1554 722
rect 1590 718 1594 722
rect 1614 718 1618 722
rect 1742 718 1746 722
rect 2006 718 2010 722
rect 2022 718 2026 722
rect 2054 718 2058 722
rect 2790 718 2794 722
rect 2878 718 2882 722
rect 3166 718 3170 722
rect 3182 718 3186 722
rect 3222 718 3226 722
rect 3318 718 3322 722
rect 3358 718 3362 722
rect 3622 718 3626 722
rect 3942 718 3946 722
rect 4246 718 4250 722
rect 4502 718 4506 722
rect 4566 718 4570 722
rect 4742 718 4746 722
rect 4814 718 4818 722
rect 4942 718 4946 722
rect 5070 718 5074 722
rect 5174 718 5178 722
rect 1050 703 1054 707
rect 1057 703 1061 707
rect 2074 703 2078 707
rect 2081 703 2085 707
rect 3098 703 3102 707
rect 3105 703 3109 707
rect 4114 703 4118 707
rect 4121 703 4125 707
rect 14 688 18 692
rect 166 688 170 692
rect 230 688 234 692
rect 574 688 578 692
rect 598 688 602 692
rect 694 688 698 692
rect 902 688 906 692
rect 942 688 946 692
rect 982 688 986 692
rect 1102 688 1106 692
rect 1150 688 1154 692
rect 1406 688 1410 692
rect 1446 688 1450 692
rect 1654 688 1658 692
rect 1702 688 1706 692
rect 1926 688 1930 692
rect 2134 688 2138 692
rect 2190 688 2194 692
rect 2286 688 2290 692
rect 2334 688 2338 692
rect 2358 688 2362 692
rect 2390 688 2394 692
rect 2414 688 2418 692
rect 2574 688 2578 692
rect 2782 688 2786 692
rect 2966 688 2970 692
rect 2990 688 2994 692
rect 3270 688 3274 692
rect 3278 688 3282 692
rect 3390 688 3394 692
rect 3398 688 3402 692
rect 3430 688 3434 692
rect 3534 688 3538 692
rect 3822 688 3826 692
rect 3870 688 3874 692
rect 4046 688 4050 692
rect 4070 688 4074 692
rect 4078 688 4082 692
rect 4190 688 4194 692
rect 4374 688 4378 692
rect 4414 688 4418 692
rect 4470 688 4474 692
rect 4486 688 4490 692
rect 4622 688 4626 692
rect 4678 688 4682 692
rect 4710 688 4714 692
rect 4862 688 4866 692
rect 4886 688 4890 692
rect 4894 688 4898 692
rect 5006 688 5010 692
rect 198 678 202 682
rect 590 678 594 682
rect 630 678 634 682
rect 758 678 762 682
rect 1022 678 1026 682
rect 1310 678 1314 682
rect 1990 678 1994 682
rect 2222 678 2226 682
rect 2350 678 2354 682
rect 3902 678 3906 682
rect 4254 678 4258 682
rect 4478 678 4482 682
rect 4582 678 4586 682
rect 4742 678 4746 682
rect 5038 678 5042 682
rect 70 668 74 672
rect 86 668 90 672
rect 182 668 186 672
rect 206 668 210 672
rect 254 668 258 672
rect 262 668 266 672
rect 294 668 298 672
rect 326 668 330 672
rect 382 668 386 672
rect 398 668 402 672
rect 430 668 434 672
rect 486 668 490 672
rect 518 668 522 672
rect 558 668 562 672
rect 582 668 586 672
rect 702 668 706 672
rect 718 668 722 672
rect 830 668 834 672
rect 886 668 890 672
rect 910 668 914 672
rect 918 668 922 672
rect 966 668 970 672
rect 990 668 994 672
rect 1134 668 1138 672
rect 110 658 114 662
rect 174 658 178 662
rect 190 658 194 662
rect 214 658 218 662
rect 270 658 274 662
rect 294 658 298 662
rect 334 658 338 662
rect 342 658 346 662
rect 382 658 386 662
rect 422 658 426 662
rect 494 658 498 662
rect 566 658 570 662
rect 638 658 642 662
rect 710 658 714 662
rect 766 658 770 662
rect 838 658 842 662
rect 846 658 850 662
rect 886 658 890 662
rect 894 658 898 662
rect 926 658 930 662
rect 1030 658 1034 662
rect 1134 658 1138 662
rect 1166 668 1170 672
rect 1230 668 1234 672
rect 1246 668 1250 672
rect 1334 668 1338 672
rect 1350 668 1354 672
rect 1390 668 1394 672
rect 1414 668 1418 672
rect 1422 668 1426 672
rect 1462 668 1466 672
rect 1486 668 1490 672
rect 1566 668 1570 672
rect 1582 668 1586 672
rect 1598 668 1602 672
rect 1630 668 1634 672
rect 1678 668 1682 672
rect 1686 668 1690 672
rect 1710 668 1714 672
rect 1766 668 1770 672
rect 1902 668 1906 672
rect 1934 668 1938 672
rect 1966 668 1970 672
rect 1998 668 2002 672
rect 2054 668 2058 672
rect 2142 668 2146 672
rect 2174 668 2178 672
rect 1166 658 1170 662
rect 1270 658 1274 662
rect 1342 658 1346 662
rect 1382 658 1386 662
rect 1430 658 1434 662
rect 1494 658 1498 662
rect 1574 658 1578 662
rect 1606 658 1610 662
rect 1670 658 1674 662
rect 1718 658 1722 662
rect 1758 658 1762 662
rect 1806 658 1810 662
rect 1822 658 1826 662
rect 1894 658 1898 662
rect 1910 658 1914 662
rect 1942 658 1946 662
rect 1974 658 1978 662
rect 2006 658 2010 662
rect 2070 659 2074 663
rect 2150 658 2154 662
rect 2166 658 2170 662
rect 2222 659 2226 663
rect 2318 668 2322 672
rect 2342 668 2346 672
rect 2366 668 2370 672
rect 2398 668 2402 672
rect 2422 668 2426 672
rect 2454 668 2458 672
rect 2518 668 2522 672
rect 2606 668 2610 672
rect 2622 668 2626 672
rect 2654 668 2658 672
rect 2662 668 2666 672
rect 2726 668 2730 672
rect 2790 668 2794 672
rect 2814 668 2818 672
rect 2902 668 2906 672
rect 2934 668 2938 672
rect 3006 668 3010 672
rect 3014 668 3018 672
rect 3046 668 3050 672
rect 3062 668 3066 672
rect 3078 668 3082 672
rect 3118 668 3122 672
rect 3158 668 3162 672
rect 3174 668 3178 672
rect 3190 668 3194 672
rect 3294 668 3298 672
rect 3310 668 3314 672
rect 3414 668 3418 672
rect 3422 668 3426 672
rect 3470 668 3474 672
rect 3494 668 3498 672
rect 3526 668 3530 672
rect 3614 668 3618 672
rect 3726 668 3730 672
rect 3742 668 3746 672
rect 3798 668 3802 672
rect 3942 668 3946 672
rect 3966 668 3970 672
rect 4054 668 4058 672
rect 4214 668 4218 672
rect 4326 668 4330 672
rect 4366 668 4370 672
rect 4438 668 4442 672
rect 4454 668 4458 672
rect 4542 668 4546 672
rect 4606 668 4610 672
rect 4614 668 4618 672
rect 4654 668 4658 672
rect 4702 668 4706 672
rect 4734 668 4738 672
rect 4766 668 4770 672
rect 4782 668 4786 672
rect 4870 668 4874 672
rect 4974 668 4978 672
rect 4998 668 5002 672
rect 5038 668 5042 672
rect 5078 668 5082 672
rect 5142 668 5146 672
rect 2294 658 2298 662
rect 2310 658 2314 662
rect 2374 658 2378 662
rect 2430 658 2434 662
rect 2446 658 2450 662
rect 2462 658 2466 662
rect 2510 659 2514 663
rect 2614 658 2618 662
rect 2638 658 2642 662
rect 2646 658 2650 662
rect 2662 658 2666 662
rect 2718 659 2722 663
rect 2806 658 2810 662
rect 2822 658 2826 662
rect 2854 658 2858 662
rect 2886 658 2890 662
rect 2926 658 2930 662
rect 2942 658 2946 662
rect 2950 658 2954 662
rect 2974 658 2978 662
rect 3022 658 3026 662
rect 3094 658 3098 662
rect 3126 658 3130 662
rect 3166 658 3170 662
rect 3206 659 3210 663
rect 3326 659 3330 663
rect 3438 658 3442 662
rect 3478 658 3482 662
rect 3518 658 3522 662
rect 3590 658 3594 662
rect 3678 658 3682 662
rect 3702 658 3706 662
rect 3742 658 3746 662
rect 3790 658 3794 662
rect 3814 658 3818 662
rect 3838 658 3842 662
rect 3846 658 3850 662
rect 3854 658 3858 662
rect 3886 658 3890 662
rect 3894 658 3898 662
rect 3918 658 3922 662
rect 3934 658 3938 662
rect 3950 658 3954 662
rect 3982 659 3986 663
rect 4134 658 4138 662
rect 4158 659 4162 663
rect 4206 658 4210 662
rect 4222 658 4226 662
rect 4318 658 4322 662
rect 4390 658 4394 662
rect 4398 658 4402 662
rect 4422 658 4426 662
rect 4446 658 4450 662
rect 4534 658 4538 662
rect 4582 658 4586 662
rect 4606 658 4610 662
rect 4694 658 4698 662
rect 4726 658 4730 662
rect 4750 658 4754 662
rect 4766 658 4770 662
rect 4798 659 4802 663
rect 4942 658 4946 662
rect 4990 658 4994 662
rect 5022 658 5026 662
rect 5054 658 5058 662
rect 5062 658 5066 662
rect 5126 658 5130 662
rect 5150 658 5154 662
rect 238 648 242 652
rect 286 648 290 652
rect 302 648 306 652
rect 318 648 322 652
rect 350 648 354 652
rect 510 648 514 652
rect 726 648 730 652
rect 862 648 866 652
rect 950 648 954 652
rect 974 648 978 652
rect 1110 648 1114 652
rect 1142 648 1146 652
rect 1446 648 1450 652
rect 1590 648 1594 652
rect 1622 648 1626 652
rect 1646 648 1650 652
rect 1702 648 1706 652
rect 1758 648 1762 652
rect 1926 648 1930 652
rect 1942 648 1946 652
rect 1958 648 1962 652
rect 1990 648 1994 652
rect 2006 648 2010 652
rect 2030 648 2034 652
rect 2174 648 2178 652
rect 2190 648 2194 652
rect 2326 648 2330 652
rect 2390 648 2394 652
rect 2446 648 2450 652
rect 2462 648 2466 652
rect 2478 648 2482 652
rect 2598 648 2602 652
rect 2686 648 2690 652
rect 2926 648 2930 652
rect 3142 648 3146 652
rect 3502 648 3506 652
rect 3750 648 3754 652
rect 3774 648 3778 652
rect 4070 648 4074 652
rect 4190 648 4194 652
rect 4382 648 4386 652
rect 4462 648 4466 652
rect 4646 648 4650 652
rect 4670 648 4674 652
rect 4710 648 4714 652
rect 4886 648 4890 652
rect 5070 648 5074 652
rect 358 638 362 642
rect 374 638 378 642
rect 462 638 466 642
rect 478 638 482 642
rect 550 638 554 642
rect 822 638 826 642
rect 1326 638 1330 642
rect 1366 638 1370 642
rect 1398 638 1402 642
rect 1542 638 1546 642
rect 1606 638 1610 642
rect 1734 638 1738 642
rect 1774 638 1778 642
rect 2118 638 2122 642
rect 2414 638 2418 642
rect 2630 638 2634 642
rect 2990 638 2994 642
rect 3046 638 3050 642
rect 3278 638 3282 642
rect 3398 638 3402 642
rect 3550 638 3554 642
rect 2670 628 2674 632
rect 14 618 18 622
rect 270 618 274 622
rect 1878 618 1882 622
rect 2838 618 2842 622
rect 2870 618 2874 622
rect 3430 618 3434 622
rect 3454 618 3458 622
rect 4094 618 4098 622
rect 4238 618 4242 622
rect 538 603 542 607
rect 545 603 549 607
rect 1562 603 1566 607
rect 1569 603 1573 607
rect 2586 603 2590 607
rect 2593 603 2597 607
rect 3610 603 3614 607
rect 3617 603 3621 607
rect 4634 603 4638 607
rect 4641 603 4645 607
rect 174 588 178 592
rect 446 588 450 592
rect 542 588 546 592
rect 750 588 754 592
rect 814 588 818 592
rect 846 588 850 592
rect 870 588 874 592
rect 902 588 906 592
rect 966 588 970 592
rect 1038 588 1042 592
rect 1094 588 1098 592
rect 1126 588 1130 592
rect 1190 588 1194 592
rect 1270 588 1274 592
rect 1494 588 1498 592
rect 1646 588 1650 592
rect 1662 588 1666 592
rect 1982 588 1986 592
rect 2238 588 2242 592
rect 2350 588 2354 592
rect 2446 588 2450 592
rect 2574 588 2578 592
rect 2598 588 2602 592
rect 2614 588 2618 592
rect 2886 588 2890 592
rect 2998 588 3002 592
rect 3006 588 3010 592
rect 3182 588 3186 592
rect 3310 588 3314 592
rect 3398 588 3402 592
rect 3494 588 3498 592
rect 3534 588 3538 592
rect 3574 588 3578 592
rect 3734 588 3738 592
rect 3742 588 3746 592
rect 3862 588 3866 592
rect 3886 588 3890 592
rect 4014 588 4018 592
rect 4150 588 4154 592
rect 4182 588 4186 592
rect 4206 588 4210 592
rect 4278 588 4282 592
rect 4414 588 4418 592
rect 4686 588 4690 592
rect 4750 588 4754 592
rect 262 578 266 582
rect 1470 578 1474 582
rect 3910 578 3914 582
rect 94 568 98 572
rect 134 568 138 572
rect 230 568 234 572
rect 430 568 434 572
rect 590 568 594 572
rect 926 568 930 572
rect 1318 568 1322 572
rect 1358 568 1362 572
rect 1702 568 1706 572
rect 1806 568 1810 572
rect 1822 568 1826 572
rect 1854 568 1858 572
rect 1966 568 1970 572
rect 2006 568 2010 572
rect 2086 568 2090 572
rect 2222 568 2226 572
rect 3774 568 3778 572
rect 3830 568 3834 572
rect 4070 568 4074 572
rect 4094 568 4098 572
rect 4670 568 4674 572
rect 4934 568 4938 572
rect 5086 568 5090 572
rect 110 558 114 562
rect 38 548 42 552
rect 110 548 114 552
rect 150 548 154 552
rect 198 548 202 552
rect 206 548 210 552
rect 254 548 258 552
rect 310 548 314 552
rect 382 547 386 551
rect 478 547 482 551
rect 574 548 578 552
rect 614 558 618 562
rect 630 558 634 562
rect 758 558 762 562
rect 774 558 778 562
rect 798 558 802 562
rect 830 558 834 562
rect 886 558 890 562
rect 910 558 914 562
rect 990 558 994 562
rect 1022 558 1026 562
rect 1206 558 1210 562
rect 614 548 618 552
rect 646 548 650 552
rect 686 547 690 551
rect 830 548 834 552
rect 846 548 850 552
rect 870 548 874 552
rect 926 548 930 552
rect 942 548 946 552
rect 950 548 954 552
rect 974 548 978 552
rect 998 548 1002 552
rect 1014 548 1018 552
rect 1038 548 1042 552
rect 1070 548 1074 552
rect 1078 548 1082 552
rect 1102 548 1106 552
rect 1150 548 1154 552
rect 1174 548 1178 552
rect 1190 548 1194 552
rect 1238 548 1242 552
rect 1246 548 1250 552
rect 1254 548 1258 552
rect 1278 548 1282 552
rect 1294 548 1298 552
rect 1454 558 1458 562
rect 1486 558 1490 562
rect 1670 558 1674 562
rect 1334 548 1338 552
rect 1342 548 1346 552
rect 1414 548 1418 552
rect 1478 548 1482 552
rect 1534 548 1538 552
rect 1598 548 1602 552
rect 1670 548 1674 552
rect 1686 548 1690 552
rect 1694 548 1698 552
rect 1718 548 1722 552
rect 1766 548 1770 552
rect 1838 548 1842 552
rect 2022 558 2026 562
rect 1878 548 1882 552
rect 1926 548 1930 552
rect 2014 548 2018 552
rect 2022 548 2026 552
rect 2038 548 2042 552
rect 2054 548 2058 552
rect 2302 558 2306 562
rect 2334 558 2338 562
rect 2478 558 2482 562
rect 2822 558 2826 562
rect 2990 558 2994 562
rect 3214 558 3218 562
rect 3326 558 3330 562
rect 3342 558 3346 562
rect 3350 558 3354 562
rect 3366 558 3370 562
rect 3382 558 3386 562
rect 3438 558 3442 562
rect 3470 558 3474 562
rect 3526 558 3530 562
rect 3542 558 3546 562
rect 3638 558 3642 562
rect 3758 558 3762 562
rect 3790 558 3794 562
rect 3846 558 3850 562
rect 3878 558 3882 562
rect 4030 558 4034 562
rect 4110 558 4114 562
rect 2110 548 2114 552
rect 2118 548 2122 552
rect 2166 548 2170 552
rect 2246 548 2250 552
rect 2270 548 2274 552
rect 2310 548 2314 552
rect 2334 548 2338 552
rect 2398 548 2402 552
rect 2462 548 2466 552
rect 2478 548 2482 552
rect 14 538 18 542
rect 46 538 50 542
rect 102 538 106 542
rect 158 538 162 542
rect 198 538 202 542
rect 222 538 226 542
rect 254 538 258 542
rect 342 538 346 542
rect 462 538 466 542
rect 502 538 506 542
rect 566 538 570 542
rect 622 538 626 542
rect 638 538 642 542
rect 654 538 658 542
rect 670 538 674 542
rect 774 538 778 542
rect 782 538 786 542
rect 822 538 826 542
rect 854 538 858 542
rect 862 538 866 542
rect 934 538 938 542
rect 1014 538 1018 542
rect 1046 538 1050 542
rect 1150 538 1154 542
rect 1182 538 1186 542
rect 1214 538 1218 542
rect 1294 538 1298 542
rect 1350 538 1354 542
rect 1414 538 1418 542
rect 1478 538 1482 542
rect 1502 538 1506 542
rect 1566 538 1570 542
rect 2510 547 2514 551
rect 2694 547 2698 551
rect 2742 548 2746 552
rect 2782 548 2786 552
rect 2806 548 2810 552
rect 2830 548 2834 552
rect 2918 548 2922 552
rect 2950 548 2954 552
rect 2966 548 2970 552
rect 2974 548 2978 552
rect 3038 548 3042 552
rect 3070 547 3074 551
rect 3134 548 3138 552
rect 3166 548 3170 552
rect 3198 548 3202 552
rect 3254 548 3258 552
rect 3270 548 3274 552
rect 3326 548 3330 552
rect 3374 548 3378 552
rect 3398 548 3402 552
rect 3422 548 3426 552
rect 3438 548 3442 552
rect 3454 548 3458 552
rect 3486 548 3490 552
rect 3510 548 3514 552
rect 3518 548 3522 552
rect 3574 548 3578 552
rect 3622 548 3626 552
rect 3678 548 3682 552
rect 3702 548 3706 552
rect 3782 548 3786 552
rect 3790 548 3794 552
rect 3806 548 3810 552
rect 3822 548 3826 552
rect 3862 548 3866 552
rect 3886 548 3890 552
rect 3958 548 3962 552
rect 4014 548 4018 552
rect 4038 548 4042 552
rect 4054 548 4058 552
rect 4166 558 4170 562
rect 4198 558 4202 562
rect 4390 558 4394 562
rect 4398 558 4402 562
rect 4446 558 4450 562
rect 4622 558 4626 562
rect 4654 558 4658 562
rect 4150 548 4154 552
rect 4182 548 4186 552
rect 4238 548 4242 552
rect 4270 548 4274 552
rect 4318 548 4322 552
rect 4414 548 4418 552
rect 4446 548 4450 552
rect 4494 548 4498 552
rect 1694 538 1698 542
rect 1726 538 1730 542
rect 1742 538 1746 542
rect 1830 538 1834 542
rect 1862 538 1866 542
rect 1886 538 1890 542
rect 1902 538 1906 542
rect 1950 538 1954 542
rect 2014 538 2018 542
rect 2046 538 2050 542
rect 2054 538 2058 542
rect 2126 538 2130 542
rect 2158 538 2162 542
rect 2270 538 2274 542
rect 2278 538 2282 542
rect 2310 538 2314 542
rect 2454 538 2458 542
rect 2494 538 2498 542
rect 2750 538 2754 542
rect 2766 538 2770 542
rect 2830 538 2834 542
rect 2942 538 2946 542
rect 2958 538 2962 542
rect 3142 538 3146 542
rect 3174 538 3178 542
rect 3190 538 3194 542
rect 3318 538 3322 542
rect 3374 538 3378 542
rect 3406 538 3410 542
rect 3414 538 3418 542
rect 3446 538 3450 542
rect 3550 538 3554 542
rect 3566 538 3570 542
rect 3606 538 3610 542
rect 3630 538 3634 542
rect 3782 538 3786 542
rect 3814 538 3818 542
rect 3822 538 3826 542
rect 3854 538 3858 542
rect 3966 538 3970 542
rect 4006 538 4010 542
rect 4062 538 4066 542
rect 4094 538 4098 542
rect 4158 538 4162 542
rect 4190 538 4194 542
rect 4214 538 4218 542
rect 4262 538 4266 542
rect 4326 538 4330 542
rect 4334 538 4338 542
rect 4374 538 4378 542
rect 4422 538 4426 542
rect 4430 538 4434 542
rect 4526 547 4530 551
rect 4558 548 4562 552
rect 4606 548 4610 552
rect 4654 548 4658 552
rect 4782 548 4786 552
rect 4814 548 4818 552
rect 4838 548 4842 552
rect 4870 548 4874 552
rect 4894 548 4898 552
rect 4910 548 4914 552
rect 4926 548 4930 552
rect 4966 548 4970 552
rect 4974 548 4978 552
rect 5030 548 5034 552
rect 5054 548 5058 552
rect 5078 548 5082 552
rect 5126 548 5130 552
rect 5142 548 5146 552
rect 4478 538 4482 542
rect 4542 538 4546 542
rect 4598 538 4602 542
rect 4646 538 4650 542
rect 4742 538 4746 542
rect 4806 538 4810 542
rect 4862 538 4866 542
rect 4918 538 4922 542
rect 5038 538 5042 542
rect 166 528 170 532
rect 182 528 186 532
rect 782 528 786 532
rect 894 528 898 532
rect 1654 528 1658 532
rect 2230 528 2234 532
rect 2302 528 2306 532
rect 2342 528 2346 532
rect 2382 528 2386 532
rect 2606 528 2610 532
rect 2622 528 2626 532
rect 2694 528 2698 532
rect 2726 528 2730 532
rect 2782 528 2786 532
rect 2902 528 2906 532
rect 2990 528 2994 532
rect 3118 528 3122 532
rect 3174 528 3178 532
rect 3590 528 3594 532
rect 3750 528 3754 532
rect 3902 528 3906 532
rect 4054 528 4058 532
rect 4222 528 4226 532
rect 4758 528 4762 532
rect 4766 528 4770 532
rect 4822 528 4826 532
rect 4878 528 4882 532
rect 4998 528 5002 532
rect 5062 528 5066 532
rect 1518 518 1522 522
rect 2630 518 2634 522
rect 2934 518 2938 522
rect 3214 518 3218 522
rect 3470 518 3474 522
rect 3526 518 3530 522
rect 3550 518 3554 522
rect 3582 518 3586 522
rect 4046 518 4050 522
rect 4254 518 4258 522
rect 4278 518 4282 522
rect 4382 518 4386 522
rect 4590 518 4594 522
rect 4622 518 4626 522
rect 4798 518 4802 522
rect 4854 518 4858 522
rect 1050 503 1054 507
rect 1057 503 1061 507
rect 2074 503 2078 507
rect 2081 503 2085 507
rect 3098 503 3102 507
rect 3105 503 3109 507
rect 4114 503 4118 507
rect 4121 503 4125 507
rect 302 488 306 492
rect 478 488 482 492
rect 598 488 602 492
rect 646 488 650 492
rect 750 488 754 492
rect 886 488 890 492
rect 918 488 922 492
rect 974 488 978 492
rect 1006 488 1010 492
rect 1022 488 1026 492
rect 1062 488 1066 492
rect 1198 488 1202 492
rect 1454 488 1458 492
rect 1590 488 1594 492
rect 1798 488 1802 492
rect 1886 488 1890 492
rect 1990 488 1994 492
rect 2182 488 2186 492
rect 2206 488 2210 492
rect 2310 488 2314 492
rect 2390 488 2394 492
rect 2502 488 2506 492
rect 2622 488 2626 492
rect 2822 488 2826 492
rect 2870 488 2874 492
rect 2998 488 3002 492
rect 3254 488 3258 492
rect 3366 488 3370 492
rect 3382 488 3386 492
rect 3422 488 3426 492
rect 3510 488 3514 492
rect 3638 488 3642 492
rect 3678 488 3682 492
rect 3926 488 3930 492
rect 3990 488 3994 492
rect 4094 488 4098 492
rect 4214 488 4218 492
rect 4254 488 4258 492
rect 4366 488 4370 492
rect 4406 488 4410 492
rect 4486 488 4490 492
rect 4518 488 4522 492
rect 4662 488 4666 492
rect 4726 488 4730 492
rect 4750 488 4754 492
rect 4846 488 4850 492
rect 4942 488 4946 492
rect 5102 488 5106 492
rect 5126 488 5130 492
rect 14 478 18 482
rect 62 468 66 472
rect 94 468 98 472
rect 126 468 130 472
rect 166 468 170 472
rect 206 468 210 472
rect 318 468 322 472
rect 342 468 346 472
rect 406 468 410 472
rect 422 468 426 472
rect 462 468 466 472
rect 486 468 490 472
rect 502 468 506 472
rect 606 468 610 472
rect 654 468 658 472
rect 758 468 762 472
rect 814 468 818 472
rect 846 468 850 472
rect 902 468 906 472
rect 926 468 930 472
rect 30 458 34 462
rect 54 458 58 462
rect 70 458 74 462
rect 86 458 90 462
rect 102 458 106 462
rect 142 458 146 462
rect 150 458 154 462
rect 158 458 162 462
rect 222 459 226 463
rect 350 458 354 462
rect 414 458 418 462
rect 454 458 458 462
rect 542 458 546 462
rect 614 458 618 462
rect 638 458 642 462
rect 694 458 698 462
rect 710 458 714 462
rect 766 458 770 462
rect 806 458 810 462
rect 830 458 834 462
rect 838 458 842 462
rect 854 458 858 462
rect 878 458 882 462
rect 926 458 930 462
rect 942 478 946 482
rect 1014 478 1018 482
rect 1414 478 1418 482
rect 1630 478 1634 482
rect 1742 478 1746 482
rect 1950 478 1954 482
rect 3358 478 3362 482
rect 3470 478 3474 482
rect 950 468 954 472
rect 998 468 1002 472
rect 1038 468 1042 472
rect 1086 468 1090 472
rect 1102 468 1106 472
rect 1206 468 1210 472
rect 1214 468 1218 472
rect 1254 468 1258 472
rect 1270 468 1274 472
rect 1278 468 1282 472
rect 1342 468 1346 472
rect 1462 468 1466 472
rect 1494 468 1498 472
rect 958 458 962 462
rect 1078 458 1082 462
rect 1118 459 1122 463
rect 1222 458 1226 462
rect 1262 458 1266 462
rect 1382 458 1386 462
rect 1414 459 1418 463
rect 1526 468 1530 472
rect 1734 468 1738 472
rect 1766 468 1770 472
rect 1822 468 1826 472
rect 1862 468 1866 472
rect 1878 468 1882 472
rect 2014 468 2018 472
rect 2070 468 2074 472
rect 2262 468 2266 472
rect 2318 468 2322 472
rect 2334 468 2338 472
rect 2350 468 2354 472
rect 2374 468 2378 472
rect 2398 468 2402 472
rect 2422 468 2426 472
rect 1494 458 1498 462
rect 1502 458 1506 462
rect 1518 458 1522 462
rect 1558 458 1562 462
rect 1606 458 1610 462
rect 1646 458 1650 462
rect 1678 459 1682 463
rect 1726 458 1730 462
rect 1758 458 1762 462
rect 1774 458 1778 462
rect 1782 458 1786 462
rect 1822 458 1826 462
rect 1830 458 1834 462
rect 1878 458 1882 462
rect 1934 458 1938 462
rect 2006 458 2010 462
rect 2022 458 2026 462
rect 2054 458 2058 462
rect 2062 458 2066 462
rect 2118 459 2122 463
rect 2150 458 2154 462
rect 2190 458 2194 462
rect 2254 458 2258 462
rect 2326 458 2330 462
rect 2350 458 2354 462
rect 2366 458 2370 462
rect 2422 458 2426 462
rect 2446 468 2450 472
rect 2462 468 2466 472
rect 2510 468 2514 472
rect 2550 468 2554 472
rect 2654 468 2658 472
rect 2662 468 2666 472
rect 2694 468 2698 472
rect 2782 468 2786 472
rect 2830 468 2834 472
rect 2862 468 2866 472
rect 2918 468 2922 472
rect 2966 468 2970 472
rect 3014 468 3018 472
rect 3038 468 3042 472
rect 3086 468 3090 472
rect 3102 468 3106 472
rect 3142 468 3146 472
rect 3158 468 3162 472
rect 3174 468 3178 472
rect 3270 468 3274 472
rect 3390 468 3394 472
rect 3398 468 3402 472
rect 3430 468 3434 472
rect 3934 478 3938 482
rect 4198 478 4202 482
rect 4238 478 4242 482
rect 3494 468 3498 472
rect 3590 468 3594 472
rect 3622 468 3626 472
rect 3646 468 3650 472
rect 3742 468 3746 472
rect 3774 468 3778 472
rect 3798 468 3802 472
rect 3806 468 3810 472
rect 3846 468 3850 472
rect 3958 468 3962 472
rect 3974 468 3978 472
rect 4070 468 4074 472
rect 4086 468 4090 472
rect 4134 468 4138 472
rect 4470 478 4474 482
rect 4550 478 4554 482
rect 4654 478 4658 482
rect 4878 478 4882 482
rect 5038 478 5042 482
rect 4262 468 4266 472
rect 4390 468 4394 472
rect 4398 468 4402 472
rect 4430 468 4434 472
rect 4446 468 4450 472
rect 4478 468 4482 472
rect 4510 468 4514 472
rect 4582 468 4586 472
rect 4710 468 4714 472
rect 4742 468 4746 472
rect 4830 468 4834 472
rect 4926 468 4930 472
rect 4998 468 5002 472
rect 5062 468 5066 472
rect 5078 468 5082 472
rect 5094 468 5098 472
rect 5182 468 5186 472
rect 2438 458 2442 462
rect 2470 458 2474 462
rect 2494 458 2498 462
rect 2542 459 2546 463
rect 2622 458 2626 462
rect 2646 458 2650 462
rect 2718 458 2722 462
rect 2790 458 2794 462
rect 2798 458 2802 462
rect 2814 458 2818 462
rect 2838 458 2842 462
rect 2854 458 2858 462
rect 2934 459 2938 463
rect 2974 458 2978 462
rect 3022 458 3026 462
rect 3054 458 3058 462
rect 3110 458 3114 462
rect 3150 458 3154 462
rect 3190 459 3194 463
rect 3294 458 3298 462
rect 3406 458 3410 462
rect 3454 458 3458 462
rect 3502 458 3506 462
rect 3566 458 3570 462
rect 3654 458 3658 462
rect 3670 458 3674 462
rect 3734 458 3738 462
rect 3790 458 3794 462
rect 3814 458 3818 462
rect 3830 458 3834 462
rect 3862 459 3866 463
rect 3950 458 3954 462
rect 3982 458 3986 462
rect 4038 458 4042 462
rect 4158 458 4162 462
rect 4182 458 4186 462
rect 4222 458 4226 462
rect 4270 458 4274 462
rect 4310 458 4314 462
rect 4334 458 4338 462
rect 4374 458 4378 462
rect 4422 458 4426 462
rect 4454 458 4458 462
rect 4502 458 4506 462
rect 4534 458 4538 462
rect 4598 458 4602 462
rect 4686 458 4690 462
rect 4718 458 4722 462
rect 4798 458 4802 462
rect 4902 458 4906 462
rect 5006 459 5010 463
rect 5054 458 5058 462
rect 5086 458 5090 462
rect 38 448 42 452
rect 158 448 162 452
rect 190 448 194 452
rect 470 448 474 452
rect 614 448 618 452
rect 638 448 642 452
rect 766 448 770 452
rect 782 448 786 452
rect 790 448 794 452
rect 806 448 810 452
rect 886 448 890 452
rect 910 448 914 452
rect 982 448 986 452
rect 1054 448 1058 452
rect 1246 448 1250 452
rect 1446 448 1450 452
rect 1470 448 1474 452
rect 1486 448 1490 452
rect 1502 448 1506 452
rect 1726 448 1730 452
rect 1742 448 1746 452
rect 1846 448 1850 452
rect 2038 448 2042 452
rect 2342 448 2346 452
rect 2382 448 2386 452
rect 2406 448 2410 452
rect 2414 448 2418 452
rect 2454 448 2458 452
rect 2486 448 2490 452
rect 2494 448 2498 452
rect 2678 448 2682 452
rect 2806 448 2810 452
rect 2838 448 2842 452
rect 2990 448 2994 452
rect 3126 448 3130 452
rect 3446 448 3450 452
rect 3638 448 3642 452
rect 3774 448 3778 452
rect 3830 448 3834 452
rect 4102 448 4106 452
rect 4374 448 4378 452
rect 4414 448 4418 452
rect 4494 448 4498 452
rect 4726 448 4730 452
rect 5110 448 5114 452
rect 70 438 74 442
rect 174 438 178 442
rect 270 438 274 442
rect 286 438 290 442
rect 398 438 402 442
rect 438 438 442 442
rect 822 438 826 442
rect 1022 438 1026 442
rect 1238 438 1242 442
rect 1350 438 1354 442
rect 1614 438 1618 442
rect 1710 438 1714 442
rect 2774 438 2778 442
rect 2998 438 3002 442
rect 3374 438 3378 442
rect 4942 438 4946 442
rect 3478 428 3482 432
rect 54 418 58 422
rect 118 418 122 422
rect 1182 418 1186 422
rect 1222 418 1226 422
rect 1542 418 1546 422
rect 1990 418 1994 422
rect 2670 418 2674 422
rect 2974 418 2978 422
rect 4694 418 4698 422
rect 538 403 542 407
rect 545 403 549 407
rect 1562 403 1566 407
rect 1569 403 1573 407
rect 2586 403 2590 407
rect 2593 403 2597 407
rect 3610 403 3614 407
rect 3617 403 3621 407
rect 4634 403 4638 407
rect 4641 403 4645 407
rect 94 388 98 392
rect 158 388 162 392
rect 614 388 618 392
rect 630 388 634 392
rect 662 388 666 392
rect 790 388 794 392
rect 838 388 842 392
rect 854 388 858 392
rect 934 388 938 392
rect 1030 388 1034 392
rect 1062 388 1066 392
rect 1078 388 1082 392
rect 1222 388 1226 392
rect 1398 388 1402 392
rect 1422 388 1426 392
rect 1694 388 1698 392
rect 1718 388 1722 392
rect 1790 388 1794 392
rect 1910 388 1914 392
rect 2110 388 2114 392
rect 2358 388 2362 392
rect 2422 388 2426 392
rect 2614 388 2618 392
rect 2662 388 2666 392
rect 2758 388 2762 392
rect 2838 388 2842 392
rect 2934 388 2938 392
rect 2950 388 2954 392
rect 3158 388 3162 392
rect 3174 388 3178 392
rect 3342 388 3346 392
rect 3446 388 3450 392
rect 3574 388 3578 392
rect 3606 388 3610 392
rect 3638 388 3642 392
rect 3694 388 3698 392
rect 3862 388 3866 392
rect 4030 388 4034 392
rect 4406 388 4410 392
rect 4646 388 4650 392
rect 4814 388 4818 392
rect 4846 388 4850 392
rect 342 378 346 382
rect 598 378 602 382
rect 2022 378 2026 382
rect 2278 378 2282 382
rect 326 368 330 372
rect 390 368 394 372
rect 502 368 506 372
rect 1014 368 1018 372
rect 1110 368 1114 372
rect 1382 368 1386 372
rect 1406 368 1410 372
rect 1454 368 1458 372
rect 1542 368 1546 372
rect 1566 368 1570 372
rect 1670 368 1674 372
rect 2054 368 2058 372
rect 2094 368 2098 372
rect 2150 368 2154 372
rect 2262 368 2266 372
rect 2326 368 2330 372
rect 2342 368 2346 372
rect 2518 368 2522 372
rect 2918 368 2922 372
rect 3270 368 3274 372
rect 3502 368 3506 372
rect 3830 368 3834 372
rect 4070 368 4074 372
rect 4174 368 4178 372
rect 4414 368 4418 372
rect 4430 368 4434 372
rect 4510 368 4514 372
rect 4926 368 4930 372
rect 198 358 202 362
rect 54 348 58 352
rect 182 348 186 352
rect 358 358 362 362
rect 374 358 378 362
rect 398 358 402 362
rect 454 358 458 362
rect 470 358 474 362
rect 646 358 650 362
rect 694 358 698 362
rect 830 358 834 362
rect 886 358 890 362
rect 222 348 226 352
rect 278 348 282 352
rect 342 348 346 352
rect 374 348 378 352
rect 390 348 394 352
rect 414 348 418 352
rect 454 348 458 352
rect 470 348 474 352
rect 534 347 538 351
rect 622 348 626 352
rect 678 348 682 352
rect 686 348 690 352
rect 734 348 738 352
rect 806 348 810 352
rect 870 348 874 352
rect 1094 358 1098 362
rect 1126 358 1130 362
rect 1230 358 1234 362
rect 1438 358 1442 362
rect 1526 358 1530 362
rect 1678 358 1682 362
rect 1750 358 1754 362
rect 1766 358 1770 362
rect 1926 358 1930 362
rect 910 348 914 352
rect 974 348 978 352
rect 1078 348 1082 352
rect 1110 348 1114 352
rect 1166 348 1170 352
rect 1230 348 1234 352
rect 1246 348 1250 352
rect 1286 348 1290 352
rect 1326 348 1330 352
rect 1422 348 1426 352
rect 1454 348 1458 352
rect 1470 348 1474 352
rect 1502 348 1506 352
rect 1542 348 1546 352
rect 1606 347 1610 351
rect 1694 348 1698 352
rect 1734 348 1738 352
rect 1750 348 1754 352
rect 1766 348 1770 352
rect 1838 348 1842 352
rect 1910 348 1914 352
rect 1974 348 1978 352
rect 2038 348 2042 352
rect 2094 348 2098 352
rect 2134 348 2138 352
rect 2286 358 2290 362
rect 2374 358 2378 362
rect 2390 358 2394 362
rect 2414 358 2418 362
rect 2678 358 2682 362
rect 2694 358 2698 362
rect 2174 348 2178 352
rect 46 338 50 342
rect 102 338 106 342
rect 174 338 178 342
rect 230 338 234 342
rect 270 338 274 342
rect 334 338 338 342
rect 366 338 370 342
rect 422 338 426 342
rect 430 338 434 342
rect 462 338 466 342
rect 542 338 546 342
rect 622 338 626 342
rect 670 338 674 342
rect 710 338 714 342
rect 798 338 802 342
rect 814 338 818 342
rect 862 338 866 342
rect 918 338 922 342
rect 950 338 954 342
rect 1070 338 1074 342
rect 1102 338 1106 342
rect 1174 338 1178 342
rect 1254 338 1258 342
rect 1302 338 1306 342
rect 1430 338 1434 342
rect 1462 338 1466 342
rect 1494 338 1498 342
rect 1502 338 1506 342
rect 1534 338 1538 342
rect 1622 338 1626 342
rect 1702 338 1706 342
rect 1726 338 1730 342
rect 2214 347 2218 351
rect 2302 348 2306 352
rect 2318 348 2322 352
rect 2326 348 2330 352
rect 2342 348 2346 352
rect 2374 348 2378 352
rect 1758 338 1762 342
rect 1846 338 1850 342
rect 1942 338 1946 342
rect 2030 338 2034 342
rect 2102 338 2106 342
rect 2126 338 2130 342
rect 2182 338 2186 342
rect 2198 338 2202 342
rect 2454 347 2458 351
rect 2486 348 2490 352
rect 2558 348 2562 352
rect 2654 348 2658 352
rect 2694 348 2698 352
rect 2718 358 2722 362
rect 2790 358 2794 362
rect 2806 358 2810 362
rect 2830 358 2834 362
rect 2958 358 2962 362
rect 3014 358 3018 362
rect 2734 348 2738 352
rect 2774 348 2778 352
rect 2806 348 2810 352
rect 2878 348 2882 352
rect 2958 348 2962 352
rect 2974 348 2978 352
rect 2998 348 3002 352
rect 3286 358 3290 362
rect 3030 348 3034 352
rect 3038 348 3042 352
rect 3094 347 3098 351
rect 3214 348 3218 352
rect 3286 348 3290 352
rect 3310 358 3314 362
rect 3454 358 3458 362
rect 3486 358 3490 362
rect 3518 358 3522 362
rect 3590 358 3594 362
rect 3654 358 3658 362
rect 3686 358 3690 362
rect 3814 358 3818 362
rect 3846 358 3850 362
rect 3878 358 3882 362
rect 4198 358 4202 362
rect 4214 358 4218 362
rect 4526 358 4530 362
rect 4542 358 4546 362
rect 3326 348 3330 352
rect 3398 348 3402 352
rect 3454 348 3458 352
rect 3470 348 3474 352
rect 3502 348 3506 352
rect 3542 348 3546 352
rect 3574 348 3578 352
rect 3638 348 3642 352
rect 3670 348 3674 352
rect 3686 348 3690 352
rect 3734 348 3738 352
rect 3798 348 3802 352
rect 3814 348 3818 352
rect 3830 348 3834 352
rect 3862 348 3866 352
rect 3878 348 3882 352
rect 3934 348 3938 352
rect 2318 338 2322 342
rect 2350 338 2354 342
rect 2382 338 2386 342
rect 2686 338 2690 342
rect 2742 338 2746 342
rect 2766 338 2770 342
rect 2798 338 2802 342
rect 2854 338 2858 342
rect 2982 338 2986 342
rect 2990 338 2994 342
rect 3046 338 3050 342
rect 3062 338 3066 342
rect 3078 338 3082 342
rect 606 328 610 332
rect 654 328 658 332
rect 830 328 834 332
rect 846 328 850 332
rect 926 328 930 332
rect 1014 328 1018 332
rect 1038 328 1042 332
rect 3190 338 3194 342
rect 3238 338 3242 342
rect 3278 338 3282 342
rect 3334 338 3338 342
rect 3366 338 3370 342
rect 3478 338 3482 342
rect 3510 338 3514 342
rect 3550 338 3554 342
rect 3630 338 3634 342
rect 3662 338 3666 342
rect 3742 338 3746 342
rect 3790 338 3794 342
rect 3966 347 3970 351
rect 4038 348 4042 352
rect 4062 348 4066 352
rect 3822 338 3826 342
rect 3854 338 3858 342
rect 3910 338 3914 342
rect 3950 338 3954 342
rect 4134 347 4138 351
rect 4198 348 4202 352
rect 4206 348 4210 352
rect 4238 348 4242 352
rect 4286 348 4290 352
rect 4342 348 4346 352
rect 4398 348 4402 352
rect 4478 347 4482 351
rect 4526 348 4530 352
rect 4534 348 4538 352
rect 4558 348 4562 352
rect 4590 348 4594 352
rect 4622 348 4626 352
rect 4678 348 4682 352
rect 4694 348 4698 352
rect 4742 348 4746 352
rect 4774 348 4778 352
rect 4790 348 4794 352
rect 4798 348 4802 352
rect 4806 348 4810 352
rect 4830 348 4834 352
rect 4862 348 4866 352
rect 4870 348 4874 352
rect 4894 348 4898 352
rect 4966 348 4970 352
rect 5006 348 5010 352
rect 5054 348 5058 352
rect 5062 348 5066 352
rect 5094 348 5098 352
rect 4150 338 4154 342
rect 4206 338 4210 342
rect 4238 338 4242 342
rect 4294 338 4298 342
rect 4350 338 4354 342
rect 4494 338 4498 342
rect 4534 338 4538 342
rect 4566 338 4570 342
rect 4614 338 4618 342
rect 4758 338 4762 342
rect 4782 338 4786 342
rect 5014 338 5018 342
rect 5070 338 5074 342
rect 5182 338 5186 342
rect 1526 328 1530 332
rect 1710 328 1714 332
rect 1886 328 1890 332
rect 2118 328 2122 332
rect 2414 328 2418 332
rect 2550 328 2554 332
rect 2638 328 2642 332
rect 2750 328 2754 332
rect 2830 328 2834 332
rect 2942 328 2946 332
rect 3126 328 3130 332
rect 3166 328 3170 332
rect 3350 328 3354 332
rect 3550 328 3554 332
rect 3598 328 3602 332
rect 3918 328 3922 332
rect 4374 328 4378 332
rect 4390 328 4394 332
rect 4574 328 4578 332
rect 4766 328 4770 332
rect 4854 328 4858 332
rect 4974 328 4978 332
rect 5038 328 5042 332
rect 5110 328 5114 332
rect 206 318 210 322
rect 894 318 898 322
rect 1270 318 1274 322
rect 2158 318 2162 322
rect 2286 318 2290 322
rect 2790 318 2794 322
rect 3518 318 3522 322
rect 3902 318 3906 322
rect 4246 318 4250 322
rect 4358 318 4362 322
rect 4606 318 4610 322
rect 4750 318 4754 322
rect 4878 318 4882 322
rect 4910 318 4914 322
rect 5022 318 5026 322
rect 5078 318 5082 322
rect 5126 318 5130 322
rect 1050 303 1054 307
rect 1057 303 1061 307
rect 2074 303 2078 307
rect 2081 303 2085 307
rect 3098 303 3102 307
rect 3105 303 3109 307
rect 4114 303 4118 307
rect 4121 303 4125 307
rect 286 288 290 292
rect 422 288 426 292
rect 462 288 466 292
rect 646 288 650 292
rect 702 288 706 292
rect 878 288 882 292
rect 974 288 978 292
rect 1006 288 1010 292
rect 1070 288 1074 292
rect 1206 288 1210 292
rect 1246 288 1250 292
rect 1342 288 1346 292
rect 1518 288 1522 292
rect 1566 288 1570 292
rect 1734 288 1738 292
rect 1918 288 1922 292
rect 2382 288 2386 292
rect 2454 288 2458 292
rect 2654 288 2658 292
rect 2870 288 2874 292
rect 3126 288 3130 292
rect 3302 288 3306 292
rect 3326 288 3330 292
rect 3438 288 3442 292
rect 3454 288 3458 292
rect 3598 288 3602 292
rect 3790 288 3794 292
rect 3918 288 3922 292
rect 4070 288 4074 292
rect 4238 288 4242 292
rect 4358 288 4362 292
rect 4366 288 4370 292
rect 4462 288 4466 292
rect 4646 288 4650 292
rect 4686 288 4690 292
rect 4798 288 4802 292
rect 4910 288 4914 292
rect 5094 288 5098 292
rect 5190 288 5194 292
rect 222 278 226 282
rect 454 278 458 282
rect 1334 278 1338 282
rect 1398 278 1402 282
rect 1710 278 1714 282
rect 1742 278 1746 282
rect 3238 278 3242 282
rect 3358 278 3362 282
rect 3910 278 3914 282
rect 4190 278 4194 282
rect 4294 278 4298 282
rect 4582 278 4586 282
rect 46 268 50 272
rect 102 268 106 272
rect 158 268 162 272
rect 190 268 194 272
rect 318 268 322 272
rect 358 268 362 272
rect 446 268 450 272
rect 478 268 482 272
rect 582 268 586 272
rect 38 258 42 262
rect 110 258 114 262
rect 150 258 154 262
rect 182 258 186 262
rect 222 259 226 263
rect 638 268 642 272
rect 662 268 666 272
rect 694 268 698 272
rect 718 268 722 272
rect 726 268 730 272
rect 782 268 786 272
rect 798 268 802 272
rect 910 268 914 272
rect 982 268 986 272
rect 1062 268 1066 272
rect 1078 268 1082 272
rect 1110 268 1114 272
rect 1214 268 1218 272
rect 1230 268 1234 272
rect 1262 268 1266 272
rect 1270 268 1274 272
rect 1350 268 1354 272
rect 1462 268 1466 272
rect 1478 268 1482 272
rect 1502 268 1506 272
rect 1526 268 1530 272
rect 1534 268 1538 272
rect 1550 268 1554 272
rect 310 258 314 262
rect 374 258 378 262
rect 422 258 426 262
rect 438 258 442 262
rect 502 258 506 262
rect 566 258 570 262
rect 598 258 602 262
rect 606 258 610 262
rect 614 258 618 262
rect 630 258 634 262
rect 670 258 674 262
rect 686 258 690 262
rect 734 258 738 262
rect 774 258 778 262
rect 814 259 818 263
rect 910 259 914 263
rect 990 258 994 262
rect 1030 258 1034 262
rect 1094 258 1098 262
rect 1102 258 1106 262
rect 1150 258 1154 262
rect 1174 258 1178 262
rect 1222 258 1226 262
rect 1278 258 1282 262
rect 1302 258 1306 262
rect 1326 258 1330 262
rect 1350 258 1354 262
rect 1374 258 1378 262
rect 1414 258 1418 262
rect 1446 259 1450 263
rect 1606 268 1610 272
rect 1750 268 1754 272
rect 1806 268 1810 272
rect 1926 268 1930 272
rect 1934 268 1938 272
rect 1958 268 1962 272
rect 1982 268 1986 272
rect 2014 268 2018 272
rect 2190 268 2194 272
rect 2230 268 2234 272
rect 2286 268 2290 272
rect 2302 268 2306 272
rect 2390 268 2394 272
rect 2446 268 2450 272
rect 2486 268 2490 272
rect 2550 268 2554 272
rect 2686 268 2690 272
rect 2718 268 2722 272
rect 2726 268 2730 272
rect 2758 268 2762 272
rect 2774 268 2778 272
rect 2790 268 2794 272
rect 2902 268 2906 272
rect 2934 268 2938 272
rect 2974 268 2978 272
rect 3006 268 3010 272
rect 3078 268 3082 272
rect 3150 268 3154 272
rect 3206 268 3210 272
rect 3318 268 3322 272
rect 3366 268 3370 272
rect 3422 268 3426 272
rect 3446 268 3450 272
rect 3534 268 3538 272
rect 3550 268 3554 272
rect 3678 268 3682 272
rect 1494 258 1498 262
rect 1582 258 1586 262
rect 1598 258 1602 262
rect 1606 258 1610 262
rect 1662 259 1666 263
rect 1686 258 1690 262
rect 1758 258 1762 262
rect 1798 258 1802 262
rect 1846 258 1850 262
rect 1870 258 1874 262
rect 1966 258 1970 262
rect 2014 258 2018 262
rect 2054 258 2058 262
rect 2078 258 2082 262
rect 2166 258 2170 262
rect 2238 258 2242 262
rect 2246 258 2250 262
rect 2286 258 2290 262
rect 2318 259 2322 263
rect 2398 258 2402 262
rect 2438 258 2442 262
rect 2510 258 2514 262
rect 2598 258 2602 262
rect 2614 258 2618 262
rect 2686 258 2690 262
rect 2694 258 2698 262
rect 2710 258 2714 262
rect 2734 258 2738 262
rect 2806 259 2810 263
rect 2878 258 2882 262
rect 2902 258 2906 262
rect 2942 258 2946 262
rect 2958 258 2962 262
rect 2982 258 2986 262
rect 2998 258 3002 262
rect 3014 258 3018 262
rect 3062 259 3066 263
rect 3158 258 3162 262
rect 3198 258 3202 262
rect 3254 258 3258 262
rect 3262 258 3266 262
rect 3310 258 3314 262
rect 3342 258 3346 262
rect 3366 258 3370 262
rect 3414 258 3418 262
rect 3518 259 3522 263
rect 3558 258 3562 262
rect 3590 258 3594 262
rect 3630 258 3634 262
rect 3662 259 3666 263
rect 3718 268 3722 272
rect 3726 268 3730 272
rect 3758 268 3762 272
rect 3838 268 3842 272
rect 3894 268 3898 272
rect 4022 268 4026 272
rect 4198 268 4202 272
rect 4206 268 4210 272
rect 4262 268 4266 272
rect 4278 268 4282 272
rect 3694 258 3698 262
rect 3710 258 3714 262
rect 3726 258 3730 262
rect 3750 258 3754 262
rect 3782 258 3786 262
rect 3838 258 3842 262
rect 3886 258 3890 262
rect 3950 258 3954 262
rect 3974 258 3978 262
rect 4014 258 4018 262
rect 4046 258 4050 262
rect 4102 258 4106 262
rect 4126 258 4130 262
rect 4198 258 4202 262
rect 4254 258 4258 262
rect 4302 258 4306 262
rect 4382 258 4386 262
rect 4398 268 4402 272
rect 4454 268 4458 272
rect 4510 268 4514 272
rect 4662 268 4666 272
rect 4702 278 4706 282
rect 4806 278 4810 282
rect 4974 278 4978 282
rect 4726 268 4730 272
rect 4782 268 4786 272
rect 4894 268 4898 272
rect 5110 268 5114 272
rect 4398 258 4402 262
rect 4406 258 4410 262
rect 4446 258 4450 262
rect 4526 259 4530 263
rect 4590 258 4594 262
rect 4670 258 4674 262
rect 4718 258 4722 262
rect 4734 258 4738 262
rect 4774 258 4778 262
rect 4790 258 4794 262
rect 4870 258 4874 262
rect 4942 258 4946 262
rect 4974 259 4978 263
rect 5038 258 5042 262
rect 5062 258 5066 262
rect 5134 258 5138 262
rect 110 248 114 252
rect 134 248 138 252
rect 614 248 618 252
rect 646 248 650 252
rect 662 248 666 252
rect 702 248 706 252
rect 1014 248 1018 252
rect 1062 248 1066 252
rect 1238 248 1242 252
rect 1246 248 1250 252
rect 1278 248 1282 252
rect 1294 248 1298 252
rect 1478 248 1482 252
rect 1510 248 1514 252
rect 1550 248 1554 252
rect 1598 248 1602 252
rect 1614 248 1618 252
rect 1798 248 1802 252
rect 1910 248 1914 252
rect 1950 248 1954 252
rect 2414 248 2418 252
rect 2438 248 2442 252
rect 2678 248 2682 252
rect 2694 248 2698 252
rect 2942 248 2946 252
rect 2998 248 3002 252
rect 3014 248 3018 252
rect 3030 248 3034 252
rect 3174 248 3178 252
rect 3398 248 3402 252
rect 3430 248 3434 252
rect 3694 248 3698 252
rect 3750 248 3754 252
rect 3782 248 3786 252
rect 3910 248 3914 252
rect 4038 248 4042 252
rect 4182 248 4186 252
rect 4214 248 4218 252
rect 4230 248 4234 252
rect 4238 248 4242 252
rect 4366 248 4370 252
rect 94 238 98 242
rect 166 238 170 242
rect 294 238 298 242
rect 558 238 562 242
rect 758 238 762 242
rect 1078 238 1082 242
rect 1630 238 1634 242
rect 1726 238 1730 242
rect 1774 238 1778 242
rect 1814 238 1818 242
rect 1990 238 1994 242
rect 2022 238 2026 242
rect 2222 238 2226 242
rect 2262 238 2266 242
rect 2366 238 2370 242
rect 2758 238 2762 242
rect 2854 238 2858 242
rect 2934 238 2938 242
rect 3470 238 3474 242
rect 3734 238 3738 242
rect 4422 238 4426 242
rect 4750 238 4754 242
rect 4830 238 4834 242
rect 182 218 186 222
rect 310 218 314 222
rect 734 218 738 222
rect 878 218 882 222
rect 1310 218 1314 222
rect 1942 218 1946 222
rect 2894 218 2898 222
rect 2958 218 2962 222
rect 3198 218 3202 222
rect 3374 218 3378 222
rect 4446 218 4450 222
rect 4774 218 4778 222
rect 538 203 542 207
rect 545 203 549 207
rect 1562 203 1566 207
rect 1569 203 1573 207
rect 2586 203 2590 207
rect 2593 203 2597 207
rect 3610 203 3614 207
rect 3617 203 3621 207
rect 4634 203 4638 207
rect 4641 203 4645 207
rect 94 188 98 192
rect 326 188 330 192
rect 422 188 426 192
rect 694 188 698 192
rect 782 188 786 192
rect 1046 188 1050 192
rect 1398 188 1402 192
rect 1558 188 1562 192
rect 1830 188 1834 192
rect 2118 188 2122 192
rect 2726 188 2730 192
rect 2926 188 2930 192
rect 3078 188 3082 192
rect 3110 188 3114 192
rect 3222 188 3226 192
rect 3342 188 3346 192
rect 3534 188 3538 192
rect 3782 188 3786 192
rect 3958 188 3962 192
rect 4054 188 4058 192
rect 4214 188 4218 192
rect 4398 188 4402 192
rect 4406 188 4410 192
rect 4542 188 4546 192
rect 4814 188 4818 192
rect 4910 188 4914 192
rect 5102 188 5106 192
rect 190 178 194 182
rect 1190 178 1194 182
rect 1918 178 1922 182
rect 2702 178 2706 182
rect 5006 178 5010 182
rect 702 168 706 172
rect 758 168 762 172
rect 854 168 858 172
rect 950 168 954 172
rect 1174 168 1178 172
rect 1222 168 1226 172
rect 1358 168 1362 172
rect 1430 168 1434 172
rect 1686 168 1690 172
rect 1702 168 1706 172
rect 1766 168 1770 172
rect 1886 168 1890 172
rect 2102 168 2106 172
rect 2222 168 2226 172
rect 2254 168 2258 172
rect 2326 168 2330 172
rect 2342 168 2346 172
rect 2438 168 2442 172
rect 2646 168 2650 172
rect 2814 168 2818 172
rect 3494 168 3498 172
rect 3678 168 3682 172
rect 3854 168 3858 172
rect 4094 168 4098 172
rect 4638 168 4642 172
rect 4766 168 4770 172
rect 4870 168 4874 172
rect 198 158 202 162
rect 286 158 290 162
rect 38 148 42 152
rect 134 148 138 152
rect 198 148 202 152
rect 214 148 218 152
rect 230 148 234 152
rect 262 148 266 152
rect 278 148 282 152
rect 302 148 306 152
rect 366 148 370 152
rect 438 148 442 152
rect 446 148 450 152
rect 462 158 466 162
rect 494 158 498 162
rect 566 158 570 162
rect 598 158 602 162
rect 478 148 482 152
rect 510 148 514 152
rect 550 148 554 152
rect 582 148 586 152
rect 638 148 642 152
rect 702 148 706 152
rect 742 148 746 152
rect 822 158 826 162
rect 1094 158 1098 162
rect 798 148 802 152
rect 838 148 842 152
rect 854 148 858 152
rect 894 148 898 152
rect 918 148 922 152
rect 990 148 994 152
rect 1070 148 1074 152
rect 1094 148 1098 152
rect 1134 148 1138 152
rect 1206 148 1210 152
rect 1270 148 1274 152
rect 1294 158 1298 162
rect 1310 148 1314 152
rect 1334 148 1338 152
rect 1374 148 1378 152
rect 1414 148 1418 152
rect 1718 158 1722 162
rect 1734 158 1738 162
rect 1750 158 1754 162
rect 1774 158 1778 162
rect 1846 158 1850 162
rect 1446 148 1450 152
rect 1454 148 1458 152
rect 1494 147 1498 151
rect 1582 148 1586 152
rect 1646 148 1650 152
rect 1718 148 1722 152
rect 1750 148 1754 152
rect 1790 148 1794 152
rect 1822 148 1826 152
rect 1862 148 1866 152
rect 2134 158 2138 162
rect 2150 158 2154 162
rect 2190 158 2194 162
rect 2310 158 2314 162
rect 2654 158 2658 162
rect 2686 158 2690 162
rect 1902 148 1906 152
rect 1950 148 1954 152
rect 1974 148 1978 152
rect 2046 148 2050 152
rect 2134 148 2138 152
rect 2158 148 2162 152
rect 2166 148 2170 152
rect 2174 148 2178 152
rect 2206 148 2210 152
rect 2222 148 2226 152
rect 2238 148 2242 152
rect 2278 148 2282 152
rect 2294 148 2298 152
rect 2310 148 2314 152
rect 2326 148 2330 152
rect 14 138 18 142
rect 110 138 114 142
rect 158 138 162 142
rect 222 138 226 142
rect 238 138 242 142
rect 310 138 314 142
rect 430 138 434 142
rect 486 138 490 142
rect 518 138 522 142
rect 542 138 546 142
rect 574 138 578 142
rect 614 138 618 142
rect 734 138 738 142
rect 790 138 794 142
rect 798 138 802 142
rect 822 138 826 142
rect 830 138 834 142
rect 870 138 874 142
rect 1062 138 1066 142
rect 1198 138 1202 142
rect 1230 138 1234 142
rect 1254 138 1258 142
rect 1262 138 1266 142
rect 1278 138 1282 142
rect 1318 138 1322 142
rect 1326 138 1330 142
rect 1342 138 1346 142
rect 1382 138 1386 142
rect 1406 138 1410 142
rect 1462 138 1466 142
rect 1478 138 1482 142
rect 1606 138 1610 142
rect 1622 138 1626 142
rect 1710 138 1714 142
rect 1742 138 1746 142
rect 1798 138 1802 142
rect 1854 138 1858 142
rect 1878 138 1882 142
rect 1910 138 1914 142
rect 2126 138 2130 142
rect 2182 138 2186 142
rect 2214 138 2218 142
rect 2374 147 2378 151
rect 2478 148 2482 152
rect 2510 147 2514 151
rect 2598 148 2602 152
rect 2614 148 2618 152
rect 2654 148 2658 152
rect 2678 148 2682 152
rect 2710 148 2714 152
rect 2742 148 2746 152
rect 2766 158 2770 162
rect 2798 158 2802 162
rect 2830 158 2834 162
rect 2862 158 2866 162
rect 2902 158 2906 162
rect 2918 158 2922 162
rect 2782 148 2786 152
rect 2814 148 2818 152
rect 2846 148 2850 152
rect 2894 148 2898 152
rect 2966 148 2970 152
rect 3094 148 3098 152
rect 3142 148 3146 152
rect 3174 147 3178 151
rect 3206 148 3210 152
rect 3214 148 3218 152
rect 3238 148 3242 152
rect 3286 148 3290 152
rect 3374 148 3378 152
rect 3398 158 3402 162
rect 3422 158 3426 162
rect 3454 158 3458 162
rect 3638 158 3642 162
rect 3438 148 3442 152
rect 3494 148 3498 152
rect 3590 148 3594 152
rect 3814 158 3818 162
rect 3662 148 3666 152
rect 3726 148 3730 152
rect 3798 148 3802 152
rect 3830 148 3834 152
rect 3846 148 3850 152
rect 3886 148 3890 152
rect 3910 148 3914 152
rect 3998 148 4002 152
rect 4070 148 4074 152
rect 4190 158 4194 162
rect 4110 148 4114 152
rect 4142 148 4146 152
rect 4358 158 4362 162
rect 4742 158 4746 162
rect 4214 148 4218 152
rect 4238 148 4242 152
rect 4246 148 4250 152
rect 4254 148 4258 152
rect 4294 148 4298 152
rect 4326 147 4330 151
rect 4366 148 4370 152
rect 4374 148 4378 152
rect 4438 148 4442 152
rect 4446 148 4450 152
rect 4502 148 4506 152
rect 4598 148 4602 152
rect 4678 148 4682 152
rect 4702 147 4706 151
rect 4742 148 4746 152
rect 4782 148 4786 152
rect 4798 148 4802 152
rect 4830 148 4834 152
rect 4838 148 4842 152
rect 4854 148 4858 152
rect 4894 158 4898 162
rect 4894 148 4898 152
rect 4942 148 4946 152
rect 4966 148 4970 152
rect 5054 148 5058 152
rect 5134 148 5138 152
rect 5166 147 5170 151
rect 2246 138 2250 142
rect 2278 138 2282 142
rect 2286 138 2290 142
rect 2318 138 2322 142
rect 2358 138 2362 142
rect 2678 138 2682 142
rect 2710 138 2714 142
rect 2734 138 2738 142
rect 2750 138 2754 142
rect 2790 138 2794 142
rect 2822 138 2826 142
rect 2854 138 2858 142
rect 2886 138 2890 142
rect 2974 138 2978 142
rect 3022 138 3026 142
rect 3262 138 3266 142
rect 3382 138 3386 142
rect 3414 138 3418 142
rect 3446 138 3450 142
rect 3470 138 3474 142
rect 3590 138 3594 142
rect 3598 138 3602 142
rect 3654 138 3658 142
rect 3670 138 3674 142
rect 3742 138 3746 142
rect 3790 138 3794 142
rect 3814 138 3818 142
rect 3822 138 3826 142
rect 3950 138 3954 142
rect 3974 138 3978 142
rect 4062 138 4066 142
rect 4078 138 4082 142
rect 4118 138 4122 142
rect 4166 138 4170 142
rect 4174 138 4178 142
rect 4222 138 4226 142
rect 4230 138 4234 142
rect 4382 138 4386 142
rect 4598 138 4602 142
rect 4734 138 4738 142
rect 4790 138 4794 142
rect 4846 138 4850 142
rect 4902 138 4906 142
rect 5062 138 5066 142
rect 62 128 66 132
rect 278 128 282 132
rect 318 128 322 132
rect 358 128 362 132
rect 982 128 986 132
rect 1126 128 1130 132
rect 1390 128 1394 132
rect 1638 128 1642 132
rect 1806 128 1810 132
rect 2190 128 2194 132
rect 2718 128 2722 132
rect 3518 128 3522 132
rect 3774 128 3778 132
rect 3950 128 3954 132
rect 4390 128 4394 132
rect 246 118 250 122
rect 494 118 498 122
rect 566 118 570 122
rect 598 118 602 122
rect 1774 118 1778 122
rect 2254 118 2258 122
rect 2446 118 2450 122
rect 2830 118 2834 122
rect 2862 118 2866 122
rect 3422 118 3426 122
rect 4518 118 4522 122
rect 1050 103 1054 107
rect 1057 103 1061 107
rect 2074 103 2078 107
rect 2081 103 2085 107
rect 3098 103 3102 107
rect 3105 103 3109 107
rect 4114 103 4118 107
rect 4121 103 4125 107
rect 14 88 18 92
rect 310 88 314 92
rect 406 88 410 92
rect 534 88 538 92
rect 646 88 650 92
rect 654 88 658 92
rect 902 88 906 92
rect 1070 88 1074 92
rect 1206 88 1210 92
rect 1302 88 1306 92
rect 1326 88 1330 92
rect 1526 88 1530 92
rect 1694 88 1698 92
rect 1702 88 1706 92
rect 1798 88 1802 92
rect 1990 88 1994 92
rect 2014 88 2018 92
rect 2334 88 2338 92
rect 2430 88 2434 92
rect 2526 88 2530 92
rect 2534 88 2538 92
rect 2718 88 2722 92
rect 2886 88 2890 92
rect 2982 88 2986 92
rect 3102 88 3106 92
rect 3254 88 3258 92
rect 3438 88 3442 92
rect 3630 88 3634 92
rect 4190 88 4194 92
rect 4510 88 4514 92
rect 4526 88 4530 92
rect 4550 88 4554 92
rect 4590 88 4594 92
rect 4622 88 4626 92
rect 4806 88 4810 92
rect 4814 88 4818 92
rect 5006 88 5010 92
rect 5022 88 5026 92
rect 5054 88 5058 92
rect 5174 88 5178 92
rect 502 78 506 82
rect 718 78 722 82
rect 1358 78 1362 82
rect 1598 78 1602 82
rect 2790 78 2794 82
rect 3166 78 3170 82
rect 78 68 82 72
rect 142 68 146 72
rect 150 68 154 72
rect 230 68 234 72
rect 326 68 330 72
rect 358 68 362 72
rect 414 68 418 72
rect 454 68 458 72
rect 566 68 570 72
rect 614 68 618 72
rect 750 68 754 72
rect 806 68 810 72
rect 910 68 914 72
rect 942 68 946 72
rect 982 68 986 72
rect 1070 68 1074 72
rect 1126 68 1130 72
rect 1222 68 1226 72
rect 1318 68 1322 72
rect 1366 68 1370 72
rect 1446 68 1450 72
rect 1494 68 1498 72
rect 1542 68 1546 72
rect 1614 68 1618 72
rect 1638 68 1642 72
rect 1782 68 1786 72
rect 1822 68 1826 72
rect 1830 68 1834 72
rect 1894 68 1898 72
rect 1910 68 1914 72
rect 1958 68 1962 72
rect 2054 68 2058 72
rect 2102 68 2106 72
rect 2166 68 2170 72
rect 2174 68 2178 72
rect 2238 68 2242 72
rect 2254 68 2258 72
rect 2350 68 2354 72
rect 2446 68 2450 72
rect 2494 68 2498 72
rect 2614 68 2618 72
rect 2630 68 2634 72
rect 2670 68 2674 72
rect 2678 68 2682 72
rect 2750 68 2754 72
rect 2838 68 2842 72
rect 2934 68 2938 72
rect 2998 68 3002 72
rect 3046 68 3050 72
rect 214 58 218 62
rect 246 59 250 63
rect 358 58 362 62
rect 422 58 426 62
rect 430 58 434 62
rect 478 58 482 62
rect 598 58 602 62
rect 718 59 722 63
rect 758 58 762 62
rect 766 58 770 62
rect 798 58 802 62
rect 846 58 850 62
rect 870 58 874 62
rect 918 58 922 62
rect 934 58 938 62
rect 950 58 954 62
rect 1006 58 1010 62
rect 1110 58 1114 62
rect 1150 58 1154 62
rect 1246 58 1250 62
rect 1310 58 1314 62
rect 1342 58 1346 62
rect 1430 58 1434 62
rect 1470 58 1474 62
rect 1534 58 1538 62
rect 1566 58 1570 62
rect 1582 58 1586 62
rect 1630 59 1634 63
rect 1766 59 1770 63
rect 1798 58 1802 62
rect 1814 58 1818 62
rect 1934 58 1938 62
rect 1998 58 2002 62
rect 2022 58 2026 62
rect 2046 58 2050 62
rect 2062 58 2066 62
rect 2278 58 2282 62
rect 2374 58 2378 62
rect 2470 58 2474 62
rect 2598 59 2602 63
rect 2686 58 2690 62
rect 2734 58 2738 62
rect 2742 58 2746 62
rect 2766 58 2770 62
rect 2774 58 2778 62
rect 2822 59 2826 63
rect 3078 68 3082 72
rect 3206 68 3210 72
rect 3230 78 3234 82
rect 3446 78 3450 82
rect 3478 78 3482 82
rect 4294 78 4298 82
rect 4598 78 4602 82
rect 3470 68 3474 72
rect 3502 68 3506 72
rect 3534 68 3538 72
rect 3654 68 3658 72
rect 3710 68 3714 72
rect 3790 68 3794 72
rect 3854 68 3858 72
rect 3870 68 3874 72
rect 3982 68 3986 72
rect 2942 58 2946 62
rect 3014 58 3018 62
rect 3038 58 3042 62
rect 3054 58 3058 62
rect 3070 58 3074 62
rect 3166 59 3170 63
rect 3198 58 3202 62
rect 3230 58 3234 62
rect 3246 58 3250 62
rect 3318 59 3322 63
rect 4014 68 4018 72
rect 4022 68 4026 72
rect 4054 68 4058 72
rect 4110 68 4114 72
rect 4198 68 4202 72
rect 3382 58 3386 62
rect 3406 58 3410 62
rect 3462 58 3466 62
rect 3494 58 3498 62
rect 3502 58 3506 62
rect 3526 58 3530 62
rect 3574 58 3578 62
rect 3598 58 3602 62
rect 3662 58 3666 62
rect 3670 58 3674 62
rect 3702 58 3706 62
rect 3718 58 3722 62
rect 3902 58 3906 62
rect 3966 58 3970 62
rect 3974 58 3978 62
rect 3990 58 3994 62
rect 4006 58 4010 62
rect 4014 58 4018 62
rect 4030 58 4034 62
rect 4038 58 4042 62
rect 4062 58 4066 62
rect 4126 59 4130 63
rect 4230 68 4234 72
rect 4342 68 4346 72
rect 4358 68 4362 72
rect 4414 68 4418 72
rect 4462 68 4466 72
rect 4574 68 4578 72
rect 4702 68 4706 72
rect 4758 68 4762 72
rect 4838 68 4842 72
rect 4910 68 4914 72
rect 4958 68 4962 72
rect 5118 68 5122 72
rect 4206 58 4210 62
rect 4222 58 4226 62
rect 4238 58 4242 62
rect 4318 58 4322 62
rect 4366 58 4370 62
rect 4406 58 4410 62
rect 4446 59 4450 63
rect 4542 58 4546 62
rect 4566 58 4570 62
rect 4582 58 4586 62
rect 4686 59 4690 63
rect 4750 58 4754 62
rect 4830 58 4834 62
rect 4854 58 4858 62
rect 4950 58 4954 62
rect 5038 58 5042 62
rect 438 48 442 52
rect 782 48 786 52
rect 934 48 938 52
rect 950 48 954 52
rect 966 48 970 52
rect 2030 48 2034 52
rect 2646 48 2650 52
rect 2702 48 2706 52
rect 3022 48 3026 52
rect 3038 48 3042 52
rect 3054 48 3058 52
rect 3446 48 3450 52
rect 3478 48 3482 52
rect 3510 48 3514 52
rect 3686 48 3690 52
rect 3958 48 3962 52
rect 4046 48 4050 52
rect 4062 48 4066 52
rect 4094 48 4098 52
rect 4222 48 4226 52
rect 4238 48 4242 52
rect 4366 48 4370 52
rect 4382 48 4386 52
rect 4390 48 4394 52
rect 4406 48 4410 52
rect 4550 48 4554 52
rect 4814 48 4818 52
rect 2686 38 2690 42
rect 3950 38 3954 42
rect 3990 38 3994 42
rect 2094 18 2098 22
rect 538 3 542 7
rect 545 3 549 7
rect 1562 3 1566 7
rect 1569 3 1573 7
rect 2586 3 2590 7
rect 2593 3 2597 7
rect 3610 3 3614 7
rect 3617 3 3621 7
rect 4634 3 4638 7
rect 4641 3 4645 7
<< metal2 >>
rect 1294 4928 1298 4932
rect 2406 4931 2410 4932
rect 2406 4928 2417 4931
rect 1048 4903 1050 4907
rect 1054 4903 1057 4907
rect 1061 4903 1064 4907
rect 970 4888 974 4891
rect 846 4882 849 4888
rect 1254 4882 1257 4888
rect 834 4878 838 4881
rect 874 4878 878 4881
rect 230 4872 233 4878
rect 286 4872 289 4878
rect 78 4832 81 4868
rect 182 4862 185 4868
rect 214 4863 217 4868
rect 138 4858 142 4861
rect 246 4862 249 4868
rect 258 4858 262 4861
rect 154 4818 158 4821
rect 14 4742 17 4818
rect 190 4792 193 4848
rect 246 4842 249 4848
rect 206 4772 209 4818
rect 98 4768 102 4771
rect 134 4762 137 4768
rect 42 4748 46 4751
rect 14 4672 17 4738
rect 102 4712 105 4738
rect 110 4722 113 4748
rect 118 4742 121 4748
rect 134 4732 137 4758
rect 154 4748 158 4751
rect 162 4738 166 4741
rect 162 4728 166 4731
rect 174 4712 177 4718
rect 6 4552 9 4588
rect 14 4542 17 4668
rect 38 4662 41 4668
rect 46 4542 49 4588
rect 54 4552 57 4708
rect 94 4692 97 4698
rect 102 4682 105 4708
rect 182 4692 185 4738
rect 134 4682 137 4688
rect 190 4672 193 4748
rect 206 4702 209 4768
rect 246 4742 249 4748
rect 222 4721 225 4738
rect 214 4718 225 4721
rect 262 4722 265 4858
rect 270 4822 273 4868
rect 318 4792 321 4858
rect 374 4832 377 4868
rect 366 4812 369 4818
rect 342 4772 345 4808
rect 366 4792 369 4808
rect 310 4752 313 4758
rect 310 4742 313 4748
rect 306 4718 310 4721
rect 214 4672 217 4718
rect 122 4668 126 4671
rect 110 4662 113 4668
rect 146 4658 150 4661
rect 102 4652 105 4658
rect 94 4552 97 4558
rect 14 4472 17 4538
rect 22 4502 25 4528
rect 38 4462 41 4518
rect 46 4362 49 4538
rect 54 4422 57 4548
rect 70 4542 73 4548
rect 94 4492 97 4498
rect 102 4482 105 4648
rect 110 4472 113 4658
rect 166 4552 169 4668
rect 190 4642 193 4658
rect 246 4642 249 4658
rect 254 4652 257 4668
rect 262 4662 265 4718
rect 310 4692 313 4708
rect 318 4691 321 4748
rect 342 4692 345 4738
rect 318 4688 326 4691
rect 310 4672 313 4688
rect 318 4672 321 4678
rect 302 4662 305 4668
rect 266 4658 273 4661
rect 262 4642 265 4648
rect 262 4592 265 4628
rect 190 4552 193 4568
rect 270 4562 273 4658
rect 286 4652 289 4658
rect 278 4572 281 4578
rect 302 4552 305 4558
rect 310 4552 313 4668
rect 318 4572 321 4668
rect 326 4662 329 4688
rect 334 4552 337 4668
rect 350 4652 353 4718
rect 358 4671 361 4748
rect 366 4721 369 4738
rect 382 4732 385 4818
rect 422 4752 425 4878
rect 454 4872 457 4878
rect 598 4872 601 4878
rect 714 4868 718 4871
rect 986 4868 990 4871
rect 582 4862 585 4868
rect 570 4858 574 4861
rect 686 4862 689 4868
rect 366 4718 377 4721
rect 374 4672 377 4718
rect 358 4668 366 4671
rect 366 4662 369 4668
rect 374 4642 377 4668
rect 382 4662 385 4728
rect 398 4692 401 4747
rect 430 4712 433 4818
rect 478 4792 481 4858
rect 614 4852 617 4859
rect 706 4858 710 4861
rect 638 4852 641 4858
rect 578 4848 582 4851
rect 530 4818 534 4821
rect 502 4772 505 4818
rect 536 4803 538 4807
rect 542 4803 545 4807
rect 549 4803 552 4807
rect 558 4792 561 4848
rect 574 4772 577 4798
rect 614 4752 617 4758
rect 638 4752 641 4848
rect 694 4842 697 4858
rect 714 4848 721 4851
rect 678 4802 681 4818
rect 674 4778 678 4781
rect 686 4762 689 4768
rect 710 4762 713 4838
rect 718 4792 721 4848
rect 726 4772 729 4778
rect 702 4752 705 4758
rect 470 4732 473 4738
rect 434 4678 449 4681
rect 446 4672 449 4678
rect 462 4672 465 4718
rect 470 4682 473 4698
rect 478 4692 481 4748
rect 526 4732 529 4738
rect 434 4668 438 4671
rect 390 4662 393 4668
rect 418 4658 422 4661
rect 446 4652 449 4668
rect 118 4492 121 4548
rect 166 4542 169 4548
rect 150 4482 153 4518
rect 110 4462 113 4468
rect 130 4458 134 4461
rect 102 4422 105 4458
rect 6 4352 9 4358
rect 34 4348 38 4351
rect 6 4262 9 4348
rect 46 4342 49 4358
rect 54 4352 57 4368
rect 86 4351 89 4358
rect 22 4322 25 4328
rect 22 4192 25 4278
rect 46 4272 49 4338
rect 70 4292 73 4338
rect 70 4272 73 4288
rect 58 4258 62 4261
rect 30 4151 33 4218
rect 94 4212 97 4418
rect 150 4362 153 4478
rect 166 4472 169 4538
rect 214 4472 217 4478
rect 246 4468 254 4471
rect 158 4352 161 4368
rect 166 4342 169 4458
rect 190 4452 193 4458
rect 246 4431 249 4468
rect 278 4462 281 4548
rect 326 4542 329 4548
rect 318 4532 321 4538
rect 290 4488 294 4491
rect 258 4458 262 4461
rect 282 4448 286 4451
rect 262 4442 265 4448
rect 246 4428 257 4431
rect 186 4358 190 4361
rect 234 4348 238 4351
rect 146 4318 150 4321
rect 142 4272 145 4278
rect 166 4272 169 4338
rect 186 4328 190 4331
rect 126 4232 129 4268
rect 94 4192 97 4198
rect 90 4188 94 4191
rect 62 4152 65 4158
rect 142 4152 145 4268
rect 174 4262 177 4318
rect 206 4192 209 4338
rect 246 4332 249 4418
rect 254 4392 257 4428
rect 318 4362 321 4488
rect 334 4472 337 4528
rect 350 4522 353 4558
rect 374 4552 377 4558
rect 366 4542 369 4548
rect 382 4542 385 4578
rect 414 4542 417 4547
rect 398 4532 401 4538
rect 382 4482 385 4488
rect 422 4482 425 4538
rect 330 4468 334 4471
rect 350 4463 353 4468
rect 398 4462 401 4478
rect 422 4472 425 4478
rect 410 4468 414 4471
rect 430 4462 433 4568
rect 462 4562 465 4658
rect 486 4632 489 4668
rect 518 4662 521 4668
rect 498 4658 502 4661
rect 514 4648 518 4651
rect 526 4642 529 4728
rect 550 4722 553 4738
rect 558 4702 561 4748
rect 678 4742 681 4748
rect 686 4712 689 4748
rect 710 4712 713 4758
rect 726 4752 729 4758
rect 722 4738 726 4741
rect 566 4672 569 4708
rect 734 4692 737 4758
rect 538 4668 542 4671
rect 478 4531 481 4618
rect 518 4552 521 4628
rect 490 4548 494 4551
rect 518 4542 521 4548
rect 498 4538 502 4541
rect 526 4532 529 4638
rect 536 4603 538 4607
rect 542 4603 545 4607
rect 549 4603 552 4607
rect 566 4542 569 4668
rect 582 4622 585 4688
rect 682 4678 686 4681
rect 742 4672 745 4868
rect 786 4858 790 4861
rect 850 4858 854 4861
rect 766 4852 769 4858
rect 770 4748 774 4751
rect 750 4702 753 4748
rect 758 4742 761 4748
rect 770 4738 774 4741
rect 750 4682 753 4698
rect 782 4682 785 4798
rect 806 4762 809 4768
rect 794 4758 798 4761
rect 794 4748 798 4751
rect 798 4732 801 4738
rect 798 4712 801 4728
rect 798 4682 801 4688
rect 806 4682 809 4748
rect 814 4672 817 4858
rect 830 4832 833 4858
rect 862 4832 865 4868
rect 878 4862 881 4868
rect 894 4852 897 4868
rect 910 4852 913 4859
rect 822 4762 825 4768
rect 854 4751 857 4758
rect 658 4668 665 4671
rect 594 4658 598 4661
rect 654 4622 657 4658
rect 638 4618 646 4621
rect 478 4528 489 4531
rect 474 4518 478 4521
rect 398 4362 401 4458
rect 298 4358 302 4361
rect 274 4348 278 4351
rect 258 4338 262 4341
rect 214 4172 217 4318
rect 238 4292 241 4328
rect 262 4272 265 4278
rect 286 4272 289 4318
rect 246 4262 249 4268
rect 286 4252 289 4258
rect 222 4182 225 4218
rect 270 4162 273 4208
rect 222 4152 225 4158
rect 210 4148 214 4151
rect 38 4062 41 4068
rect 62 4062 65 4148
rect 134 4142 137 4148
rect 142 4142 145 4148
rect 234 4138 238 4141
rect 98 4088 102 4091
rect 142 4072 145 4138
rect 150 4082 153 4088
rect 166 4072 169 4078
rect 122 4068 126 4071
rect 62 3952 65 4058
rect 102 4052 105 4058
rect 98 3968 102 3971
rect 110 3952 113 4068
rect 246 4062 249 4158
rect 302 4152 305 4158
rect 294 4142 297 4148
rect 266 4138 270 4141
rect 286 4132 289 4138
rect 278 4082 281 4118
rect 310 4072 313 4338
rect 334 4332 337 4338
rect 326 4242 329 4318
rect 374 4272 377 4358
rect 382 4292 385 4348
rect 398 4342 401 4348
rect 430 4332 433 4458
rect 438 4452 441 4458
rect 446 4452 449 4458
rect 454 4441 457 4468
rect 486 4462 489 4528
rect 454 4438 465 4441
rect 446 4342 449 4348
rect 462 4342 465 4438
rect 470 4352 473 4358
rect 494 4352 497 4468
rect 502 4462 505 4518
rect 550 4492 553 4528
rect 518 4462 521 4468
rect 536 4403 538 4407
rect 542 4403 545 4407
rect 549 4403 552 4407
rect 566 4392 569 4418
rect 574 4412 577 4468
rect 582 4462 585 4618
rect 638 4572 641 4618
rect 662 4612 665 4668
rect 710 4662 713 4668
rect 766 4662 769 4668
rect 674 4658 678 4661
rect 738 4658 742 4661
rect 670 4648 678 4651
rect 670 4592 673 4648
rect 702 4642 705 4658
rect 650 4578 654 4581
rect 658 4568 662 4571
rect 590 4542 593 4548
rect 614 4472 617 4538
rect 590 4452 593 4458
rect 630 4452 633 4459
rect 598 4442 601 4448
rect 574 4362 577 4368
rect 598 4362 601 4408
rect 598 4352 601 4358
rect 614 4352 617 4438
rect 622 4372 625 4398
rect 638 4352 641 4478
rect 578 4348 582 4351
rect 646 4342 649 4528
rect 642 4338 646 4341
rect 426 4318 430 4321
rect 414 4282 417 4318
rect 362 4268 366 4271
rect 374 4262 377 4268
rect 394 4258 398 4261
rect 366 4242 369 4258
rect 326 4162 329 4218
rect 350 4162 353 4238
rect 382 4162 385 4198
rect 414 4192 417 4278
rect 542 4272 545 4338
rect 602 4288 606 4291
rect 422 4262 425 4268
rect 430 4182 433 4258
rect 438 4252 441 4258
rect 446 4221 449 4248
rect 454 4232 457 4268
rect 554 4258 558 4261
rect 574 4252 577 4288
rect 594 4268 598 4271
rect 550 4222 553 4228
rect 446 4218 457 4221
rect 426 4158 441 4161
rect 318 4142 321 4158
rect 438 4152 441 4158
rect 370 4148 374 4151
rect 426 4148 430 4151
rect 394 4138 398 4141
rect 426 4138 430 4141
rect 342 4132 345 4138
rect 134 3952 137 4058
rect 190 4052 193 4058
rect 230 3991 233 4038
rect 222 3988 233 3991
rect 98 3948 102 3951
rect 138 3948 142 3951
rect 38 3942 41 3948
rect 38 3862 41 3918
rect 62 3862 65 3948
rect 110 3942 113 3948
rect 122 3938 126 3941
rect 150 3932 153 3968
rect 162 3948 166 3951
rect 190 3942 193 3948
rect 222 3942 225 3988
rect 246 3952 249 3958
rect 166 3932 169 3938
rect 174 3922 177 3928
rect 206 3902 209 3928
rect 94 3892 97 3898
rect 106 3888 110 3891
rect 198 3882 201 3888
rect 262 3882 265 4018
rect 270 3892 273 4058
rect 302 4052 305 4058
rect 278 4042 281 4048
rect 318 4032 321 4068
rect 334 4062 337 4068
rect 326 4052 329 4058
rect 310 3962 313 4008
rect 342 3992 345 4118
rect 358 4062 361 4138
rect 374 4122 377 4138
rect 454 4092 457 4218
rect 470 4152 473 4158
rect 494 4152 497 4178
rect 510 4162 513 4218
rect 536 4203 538 4207
rect 542 4203 545 4207
rect 549 4203 552 4207
rect 478 4142 481 4148
rect 462 4112 465 4118
rect 486 4092 489 4138
rect 498 4088 502 4091
rect 382 4062 385 4068
rect 330 3938 334 3941
rect 334 3922 337 3928
rect 306 3918 310 3921
rect 182 3872 185 3878
rect 262 3862 265 3868
rect 278 3862 281 3868
rect 166 3852 169 3859
rect 226 3858 230 3861
rect 246 3852 249 3858
rect 222 3842 225 3848
rect 206 3832 209 3838
rect 246 3802 249 3848
rect 302 3822 305 3858
rect 318 3852 321 3918
rect 326 3862 329 3868
rect 334 3792 337 3818
rect 134 3752 137 3778
rect 342 3762 345 3898
rect 350 3762 353 4018
rect 374 4012 377 4058
rect 422 4052 425 4078
rect 450 4068 454 4071
rect 438 4042 441 4058
rect 454 4052 457 4058
rect 382 3962 385 3978
rect 398 3962 401 4018
rect 406 3962 409 3988
rect 462 3962 465 4058
rect 470 4042 473 4068
rect 478 4052 481 4088
rect 486 4072 489 4088
rect 510 4082 513 4118
rect 518 4092 521 4158
rect 566 4152 569 4158
rect 586 4148 590 4151
rect 526 4142 529 4148
rect 530 4118 534 4121
rect 494 4072 497 4078
rect 590 4072 593 4088
rect 614 4072 617 4338
rect 662 4302 665 4568
rect 686 4552 689 4558
rect 674 4548 678 4551
rect 678 4532 681 4538
rect 678 4442 681 4468
rect 694 4442 697 4618
rect 726 4572 729 4618
rect 758 4602 761 4658
rect 774 4652 777 4668
rect 814 4662 817 4668
rect 822 4662 825 4738
rect 846 4672 849 4708
rect 838 4662 841 4668
rect 854 4662 857 4678
rect 766 4572 769 4578
rect 790 4572 793 4618
rect 718 4562 721 4568
rect 754 4548 761 4551
rect 702 4542 705 4548
rect 746 4538 750 4541
rect 702 4482 705 4538
rect 734 4532 737 4538
rect 750 4522 753 4528
rect 758 4522 761 4548
rect 702 4462 705 4468
rect 714 4458 718 4461
rect 726 4452 729 4518
rect 750 4492 753 4518
rect 758 4482 761 4518
rect 766 4502 769 4568
rect 774 4542 777 4548
rect 790 4532 793 4548
rect 798 4542 801 4658
rect 822 4622 825 4658
rect 842 4648 846 4651
rect 854 4642 857 4648
rect 862 4632 865 4828
rect 878 4752 881 4848
rect 914 4768 918 4771
rect 958 4742 961 4838
rect 1014 4762 1017 4768
rect 886 4682 889 4688
rect 870 4642 873 4648
rect 902 4622 905 4658
rect 806 4582 809 4618
rect 798 4492 801 4538
rect 762 4478 766 4481
rect 734 4462 737 4468
rect 678 4342 681 4438
rect 694 4402 697 4418
rect 690 4348 694 4351
rect 694 4282 697 4288
rect 710 4271 713 4418
rect 738 4378 742 4381
rect 750 4362 753 4438
rect 726 4272 729 4278
rect 710 4268 721 4271
rect 654 4262 657 4268
rect 662 4142 665 4268
rect 710 4252 713 4258
rect 718 4162 721 4268
rect 734 4262 737 4268
rect 742 4262 745 4328
rect 750 4282 753 4308
rect 734 4212 737 4258
rect 758 4251 761 4398
rect 766 4381 769 4478
rect 782 4472 785 4478
rect 806 4472 809 4538
rect 814 4522 817 4548
rect 806 4432 809 4458
rect 766 4378 777 4381
rect 766 4362 769 4368
rect 774 4352 777 4378
rect 798 4372 801 4378
rect 806 4342 809 4348
rect 766 4292 769 4338
rect 758 4248 766 4251
rect 774 4242 777 4338
rect 814 4272 817 4438
rect 822 4362 825 4618
rect 834 4568 838 4571
rect 902 4562 905 4618
rect 918 4562 921 4718
rect 966 4692 969 4748
rect 1046 4742 1049 4858
rect 1070 4822 1073 4868
rect 1150 4862 1153 4868
rect 1190 4862 1193 4878
rect 1250 4868 1254 4871
rect 1234 4858 1238 4861
rect 1234 4838 1238 4841
rect 1070 4712 1073 4748
rect 1126 4732 1129 4818
rect 1214 4771 1217 4838
rect 1246 4832 1249 4868
rect 1270 4842 1273 4878
rect 1286 4862 1289 4868
rect 1294 4862 1297 4928
rect 2072 4903 2074 4907
rect 2078 4903 2081 4907
rect 2085 4903 2088 4907
rect 2414 4892 2417 4928
rect 3190 4928 3194 4932
rect 3096 4903 3098 4907
rect 3102 4903 3105 4907
rect 3109 4903 3112 4907
rect 2306 4888 2310 4891
rect 2270 4882 2273 4888
rect 1834 4878 1838 4881
rect 1502 4872 1505 4878
rect 1774 4872 1777 4878
rect 1554 4868 1558 4871
rect 1682 4868 1686 4871
rect 1354 4859 1358 4862
rect 1482 4859 1486 4862
rect 1214 4768 1225 4771
rect 1186 4758 1190 4761
rect 1150 4742 1153 4748
rect 1048 4703 1050 4707
rect 1054 4703 1057 4707
rect 1061 4703 1064 4707
rect 1086 4672 1089 4728
rect 1126 4702 1129 4718
rect 1134 4672 1137 4728
rect 1166 4692 1169 4718
rect 1158 4682 1161 4688
rect 1174 4682 1177 4758
rect 1186 4748 1190 4751
rect 1222 4742 1225 4768
rect 1286 4752 1289 4858
rect 1294 4852 1297 4858
rect 1294 4832 1297 4848
rect 1310 4822 1313 4828
rect 1314 4748 1318 4751
rect 1182 4682 1185 4738
rect 1206 4732 1209 4738
rect 1194 4718 1198 4721
rect 1246 4692 1249 4748
rect 1270 4732 1273 4738
rect 1262 4692 1265 4708
rect 1238 4682 1241 4688
rect 1278 4682 1281 4698
rect 1154 4668 1158 4671
rect 934 4663 937 4668
rect 942 4572 945 4668
rect 1006 4652 1009 4668
rect 1014 4652 1017 4658
rect 994 4638 998 4641
rect 954 4568 958 4571
rect 962 4558 966 4561
rect 990 4552 993 4638
rect 1022 4632 1025 4668
rect 850 4548 854 4551
rect 894 4542 897 4547
rect 842 4538 846 4541
rect 862 4532 865 4538
rect 878 4482 881 4538
rect 862 4442 865 4448
rect 870 4392 873 4468
rect 882 4458 889 4461
rect 886 4432 889 4458
rect 878 4422 881 4428
rect 838 4362 841 4388
rect 822 4352 825 4358
rect 834 4338 838 4341
rect 854 4322 857 4338
rect 870 4332 873 4388
rect 846 4282 849 4318
rect 886 4292 889 4347
rect 894 4342 897 4478
rect 930 4468 934 4471
rect 942 4462 945 4498
rect 966 4462 969 4548
rect 982 4532 985 4538
rect 902 4442 905 4448
rect 902 4282 905 4438
rect 918 4322 921 4458
rect 934 4452 937 4458
rect 974 4452 977 4518
rect 990 4512 993 4518
rect 982 4472 985 4508
rect 1018 4468 1022 4471
rect 982 4442 985 4458
rect 1002 4448 1006 4451
rect 1014 4422 1017 4458
rect 958 4372 961 4418
rect 1030 4392 1033 4548
rect 1070 4542 1073 4668
rect 1190 4662 1193 4668
rect 1082 4658 1086 4661
rect 1202 4658 1206 4661
rect 1218 4658 1222 4661
rect 1142 4652 1145 4658
rect 1134 4642 1137 4648
rect 1142 4612 1145 4648
rect 1198 4612 1201 4648
rect 1230 4642 1233 4678
rect 1254 4662 1257 4668
rect 1246 4622 1249 4658
rect 1048 4503 1050 4507
rect 1054 4503 1057 4507
rect 1061 4503 1064 4507
rect 1038 4402 1041 4458
rect 990 4362 993 4368
rect 1002 4358 1006 4361
rect 1014 4352 1017 4358
rect 986 4348 990 4351
rect 958 4332 961 4338
rect 966 4322 969 4348
rect 994 4338 998 4341
rect 782 4262 785 4268
rect 798 4262 801 4268
rect 830 4262 833 4268
rect 878 4262 881 4268
rect 810 4258 814 4261
rect 758 4202 761 4218
rect 782 4192 785 4248
rect 822 4232 825 4258
rect 854 4252 857 4258
rect 870 4252 873 4258
rect 738 4168 742 4171
rect 674 4148 678 4151
rect 626 4088 630 4091
rect 538 4068 542 4071
rect 582 4062 585 4068
rect 518 4052 521 4058
rect 530 4048 534 4051
rect 494 4042 497 4048
rect 574 4042 577 4048
rect 536 4003 538 4007
rect 542 4003 545 4007
rect 549 4003 552 4007
rect 362 3958 366 3961
rect 362 3948 366 3951
rect 374 3942 377 3958
rect 406 3952 409 3958
rect 442 3948 446 3951
rect 454 3942 457 3958
rect 462 3952 465 3958
rect 542 3952 545 3958
rect 590 3952 593 4058
rect 606 4048 614 4051
rect 598 3962 601 4018
rect 606 3992 609 4048
rect 630 3991 633 4078
rect 638 4062 641 4138
rect 662 4092 665 4138
rect 694 4092 697 4098
rect 742 4092 745 4158
rect 750 4142 753 4148
rect 758 4131 761 4148
rect 766 4142 769 4168
rect 806 4162 809 4188
rect 838 4152 841 4158
rect 846 4152 849 4218
rect 894 4162 897 4278
rect 902 4262 905 4268
rect 918 4262 921 4278
rect 950 4272 953 4318
rect 970 4278 974 4281
rect 990 4272 993 4328
rect 998 4272 1001 4318
rect 934 4262 937 4268
rect 958 4262 961 4268
rect 910 4152 913 4198
rect 926 4192 929 4258
rect 990 4242 993 4268
rect 998 4262 1001 4268
rect 934 4192 937 4238
rect 786 4148 790 4151
rect 822 4142 825 4148
rect 750 4128 761 4131
rect 830 4132 833 4148
rect 878 4141 881 4148
rect 878 4138 894 4141
rect 918 4132 921 4138
rect 682 4068 686 4071
rect 670 4062 673 4068
rect 710 4062 713 4078
rect 638 4022 641 4058
rect 646 4052 649 4058
rect 734 4052 737 4068
rect 718 4042 721 4048
rect 742 4042 745 4048
rect 750 4042 753 4128
rect 774 4072 777 4088
rect 626 3988 633 3991
rect 726 3961 729 4018
rect 742 3992 745 4038
rect 758 4032 761 4068
rect 722 3958 729 3961
rect 614 3952 617 3958
rect 678 3952 681 3958
rect 734 3942 737 3948
rect 774 3942 777 4068
rect 798 4062 801 4068
rect 846 3992 849 4118
rect 878 4092 881 4128
rect 886 4122 889 4128
rect 858 4088 862 4091
rect 854 4078 862 4081
rect 854 4072 857 4078
rect 886 4072 889 4118
rect 898 4068 902 4071
rect 914 4068 918 4071
rect 862 4052 865 4068
rect 926 4062 929 4148
rect 886 4042 889 4058
rect 918 4052 921 4058
rect 942 4042 945 4208
rect 950 4172 953 4218
rect 982 4162 985 4218
rect 1006 4162 1009 4318
rect 1014 4242 1017 4248
rect 954 4158 958 4161
rect 1022 4152 1025 4368
rect 1030 4252 1033 4348
rect 1038 4342 1041 4388
rect 1070 4342 1073 4538
rect 1102 4472 1105 4478
rect 1094 4462 1097 4468
rect 1086 4402 1089 4418
rect 1098 4348 1102 4351
rect 1094 4312 1097 4338
rect 1110 4322 1113 4458
rect 1126 4452 1129 4518
rect 1134 4492 1137 4548
rect 1126 4392 1129 4448
rect 1142 4332 1145 4608
rect 1158 4552 1161 4558
rect 1182 4492 1185 4608
rect 1198 4562 1201 4568
rect 1214 4562 1217 4568
rect 1222 4542 1225 4578
rect 1246 4562 1249 4568
rect 1234 4548 1238 4551
rect 1190 4512 1193 4518
rect 1158 4472 1161 4488
rect 1170 4468 1174 4471
rect 1190 4462 1193 4468
rect 1166 4432 1169 4458
rect 1186 4448 1198 4451
rect 1202 4448 1206 4451
rect 1166 4352 1169 4428
rect 1174 4352 1177 4358
rect 1166 4342 1169 4348
rect 1158 4332 1161 4338
rect 1182 4322 1185 4358
rect 1190 4332 1193 4388
rect 1206 4342 1209 4398
rect 1214 4392 1217 4538
rect 1242 4528 1246 4531
rect 1222 4462 1225 4468
rect 1230 4462 1233 4518
rect 1238 4472 1241 4478
rect 1230 4452 1233 4458
rect 1270 4452 1273 4459
rect 1226 4358 1230 4361
rect 1214 4342 1217 4348
rect 1230 4342 1233 4348
rect 1262 4342 1265 4347
rect 1214 4331 1217 4338
rect 1206 4328 1217 4331
rect 1048 4303 1050 4307
rect 1054 4303 1057 4307
rect 1061 4303 1064 4307
rect 1094 4282 1097 4308
rect 1050 4268 1054 4271
rect 1098 4259 1102 4262
rect 1150 4262 1153 4318
rect 1166 4272 1169 4288
rect 1190 4272 1193 4278
rect 1170 4268 1174 4271
rect 1038 4252 1041 4258
rect 1054 4252 1057 4258
rect 1166 4252 1169 4258
rect 1186 4248 1190 4251
rect 1154 4238 1158 4241
rect 1170 4188 1174 4191
rect 1198 4181 1201 4318
rect 1206 4292 1209 4328
rect 1206 4252 1209 4258
rect 1190 4178 1201 4181
rect 1046 4152 1049 4168
rect 1182 4162 1185 4168
rect 1110 4152 1113 4158
rect 986 4148 990 4151
rect 1178 4148 1182 4151
rect 950 4132 953 4148
rect 1014 4142 1017 4148
rect 986 4138 990 4141
rect 1170 4138 1174 4141
rect 950 4062 953 4108
rect 786 3948 790 3951
rect 410 3938 414 3941
rect 470 3938 478 3941
rect 594 3938 598 3941
rect 398 3932 401 3938
rect 366 3872 369 3878
rect 374 3862 377 3868
rect 390 3852 393 3918
rect 410 3878 417 3881
rect 414 3862 417 3878
rect 402 3848 406 3851
rect 362 3818 366 3821
rect 374 3812 377 3818
rect 310 3752 313 3758
rect 38 3748 46 3751
rect 6 3692 9 3718
rect 38 3692 41 3748
rect 6 3682 9 3688
rect 86 3672 89 3738
rect 206 3732 209 3738
rect 238 3692 241 3747
rect 46 3662 49 3668
rect 54 3662 57 3668
rect 26 3658 30 3661
rect 6 3542 9 3598
rect 86 3542 89 3668
rect 94 3662 97 3678
rect 174 3672 177 3678
rect 150 3642 153 3648
rect 6 3501 9 3538
rect 6 3498 17 3501
rect 6 3452 9 3488
rect 14 3341 17 3498
rect 62 3472 65 3518
rect 86 3472 89 3538
rect 110 3492 113 3548
rect 70 3463 73 3468
rect 118 3462 121 3628
rect 150 3552 153 3568
rect 158 3542 161 3668
rect 166 3632 169 3658
rect 190 3642 193 3648
rect 190 3612 193 3638
rect 198 3551 201 3558
rect 182 3542 185 3548
rect 166 3522 169 3528
rect 126 3472 129 3498
rect 166 3472 169 3478
rect 154 3468 158 3471
rect 174 3462 177 3518
rect 190 3482 193 3488
rect 106 3458 110 3461
rect 166 3458 174 3461
rect 102 3442 105 3448
rect 118 3422 121 3458
rect 134 3452 137 3458
rect 150 3432 153 3438
rect 158 3432 161 3458
rect 10 3338 17 3341
rect 94 3342 97 3348
rect 6 3262 9 3338
rect 14 3241 17 3298
rect 62 3272 65 3318
rect 78 3312 81 3328
rect 78 3302 81 3308
rect 110 3262 113 3318
rect 118 3292 121 3338
rect 126 3302 129 3348
rect 166 3332 169 3458
rect 198 3442 201 3528
rect 206 3461 209 3658
rect 214 3472 217 3668
rect 222 3662 225 3668
rect 230 3662 233 3668
rect 222 3502 225 3658
rect 246 3572 249 3738
rect 298 3718 302 3721
rect 270 3682 273 3718
rect 302 3712 305 3718
rect 310 3682 313 3748
rect 382 3742 385 3748
rect 390 3742 393 3828
rect 422 3822 425 3938
rect 430 3892 433 3938
rect 438 3882 441 3918
rect 470 3912 473 3938
rect 566 3932 569 3938
rect 670 3932 673 3938
rect 482 3918 486 3921
rect 566 3872 569 3928
rect 742 3922 745 3938
rect 662 3892 665 3898
rect 490 3868 494 3871
rect 486 3862 489 3868
rect 478 3822 481 3858
rect 414 3792 417 3818
rect 406 3782 409 3788
rect 430 3762 433 3798
rect 410 3748 414 3751
rect 354 3738 358 3741
rect 238 3482 241 3488
rect 246 3482 249 3568
rect 226 3478 230 3481
rect 226 3468 230 3471
rect 206 3458 214 3461
rect 202 3438 206 3441
rect 214 3432 217 3458
rect 246 3442 249 3448
rect 226 3378 230 3381
rect 238 3362 241 3368
rect 174 3352 177 3358
rect 230 3342 233 3348
rect 238 3332 241 3348
rect 134 3272 137 3278
rect 158 3272 161 3328
rect 118 3262 121 3268
rect 70 3252 73 3259
rect 162 3258 166 3261
rect 106 3248 110 3251
rect 10 3238 17 3241
rect 62 3162 65 3168
rect 74 3158 78 3161
rect 86 3152 89 3248
rect 110 3172 113 3218
rect 110 3158 118 3161
rect 22 3142 25 3148
rect 6 3092 9 3128
rect 6 3082 9 3088
rect 38 3061 41 3118
rect 38 3058 46 3061
rect 10 2978 14 2981
rect 14 2932 17 2948
rect 54 2922 57 3138
rect 62 3042 65 3148
rect 102 3142 105 3148
rect 94 3132 97 3138
rect 110 3092 113 3158
rect 174 3152 177 3258
rect 118 3142 121 3148
rect 122 3128 126 3131
rect 174 3082 177 3088
rect 86 3062 89 3068
rect 118 3062 121 3068
rect 126 3062 129 3078
rect 158 3062 161 3078
rect 170 3058 174 3061
rect 70 2951 73 2958
rect 86 2942 89 3058
rect 102 2982 105 3048
rect 150 2982 153 3018
rect 10 2888 14 2891
rect 70 2863 73 2898
rect 86 2882 89 2938
rect 102 2932 105 2978
rect 182 2952 185 3288
rect 214 3282 217 3288
rect 222 3272 225 3298
rect 198 3152 201 3158
rect 206 3072 209 3128
rect 206 3062 209 3068
rect 206 2952 209 3038
rect 178 2948 182 2951
rect 118 2922 121 2948
rect 126 2942 129 2948
rect 150 2942 153 2948
rect 198 2942 201 2948
rect 142 2922 145 2938
rect 158 2892 161 2928
rect 190 2902 193 2918
rect 86 2872 89 2878
rect 102 2862 105 2868
rect 134 2862 137 2888
rect 158 2872 161 2878
rect 182 2862 185 2888
rect 110 2851 113 2858
rect 102 2848 113 2851
rect 6 2742 9 2748
rect 74 2738 78 2741
rect 38 2662 41 2668
rect 62 2662 65 2718
rect 102 2682 105 2848
rect 126 2702 129 2818
rect 134 2742 137 2748
rect 142 2672 145 2838
rect 158 2742 161 2748
rect 182 2742 185 2748
rect 122 2668 126 2671
rect 142 2662 145 2668
rect 150 2662 153 2668
rect 182 2662 185 2688
rect 194 2678 198 2681
rect 206 2672 209 2948
rect 214 2942 217 3108
rect 222 2942 225 3268
rect 230 3262 233 3328
rect 254 3302 257 3658
rect 278 3652 281 3668
rect 318 3662 321 3738
rect 398 3732 401 3738
rect 334 3702 337 3728
rect 350 3682 353 3718
rect 366 3702 369 3718
rect 358 3692 361 3698
rect 362 3658 366 3661
rect 278 3602 281 3648
rect 318 3572 321 3578
rect 262 3562 265 3568
rect 294 3562 297 3568
rect 330 3558 334 3561
rect 302 3552 305 3558
rect 290 3548 294 3551
rect 270 3532 273 3538
rect 278 3522 281 3548
rect 278 3472 281 3478
rect 262 3462 265 3468
rect 302 3462 305 3468
rect 262 3442 265 3448
rect 318 3432 321 3548
rect 326 3482 329 3538
rect 262 3372 265 3378
rect 254 3262 257 3288
rect 262 3282 265 3368
rect 278 3352 281 3428
rect 326 3362 329 3458
rect 278 3262 281 3348
rect 286 3322 289 3338
rect 286 3282 289 3288
rect 302 3282 305 3338
rect 318 3311 321 3347
rect 326 3342 329 3358
rect 310 3308 321 3311
rect 310 3292 313 3308
rect 318 3272 321 3298
rect 342 3292 345 3658
rect 374 3652 377 3688
rect 390 3632 393 3668
rect 406 3662 409 3688
rect 422 3661 425 3758
rect 430 3752 433 3758
rect 446 3732 449 3738
rect 446 3662 449 3668
rect 422 3658 430 3661
rect 438 3642 441 3658
rect 462 3651 465 3818
rect 486 3742 489 3858
rect 554 3818 561 3821
rect 536 3803 538 3807
rect 542 3803 545 3807
rect 549 3803 552 3807
rect 502 3692 505 3748
rect 558 3732 561 3818
rect 542 3702 545 3718
rect 482 3668 486 3671
rect 474 3658 478 3661
rect 462 3648 473 3651
rect 354 3558 358 3561
rect 354 3538 358 3541
rect 374 3532 377 3608
rect 382 3572 385 3618
rect 398 3552 401 3638
rect 454 3632 457 3648
rect 418 3618 422 3621
rect 454 3582 457 3618
rect 470 3592 473 3648
rect 486 3592 489 3658
rect 446 3562 449 3568
rect 410 3558 414 3561
rect 430 3552 433 3558
rect 502 3552 505 3648
rect 510 3572 513 3698
rect 566 3672 569 3868
rect 590 3792 593 3868
rect 718 3862 721 3918
rect 742 3902 745 3918
rect 774 3872 777 3938
rect 822 3871 825 3988
rect 838 3962 841 3968
rect 846 3942 849 3978
rect 874 3968 878 3971
rect 854 3952 857 3958
rect 866 3948 870 3951
rect 850 3938 854 3941
rect 814 3868 825 3871
rect 838 3882 841 3908
rect 838 3872 841 3878
rect 878 3872 881 3968
rect 726 3862 729 3868
rect 814 3862 817 3868
rect 602 3858 606 3861
rect 786 3858 790 3861
rect 866 3858 870 3861
rect 702 3832 705 3858
rect 822 3852 825 3858
rect 686 3792 689 3818
rect 590 3762 593 3788
rect 654 3762 657 3768
rect 710 3752 713 3758
rect 742 3752 745 3788
rect 686 3742 689 3748
rect 574 3672 577 3718
rect 562 3658 566 3661
rect 526 3592 529 3638
rect 536 3603 538 3607
rect 542 3603 545 3607
rect 549 3603 552 3607
rect 606 3592 609 3658
rect 630 3592 633 3698
rect 642 3668 646 3671
rect 582 3552 585 3558
rect 398 3542 401 3548
rect 358 3492 361 3528
rect 366 3472 369 3518
rect 386 3468 390 3471
rect 378 3458 382 3461
rect 298 3268 302 3271
rect 330 3268 334 3271
rect 242 3258 246 3261
rect 230 3192 233 3258
rect 254 3252 257 3258
rect 246 3242 249 3248
rect 270 3232 273 3238
rect 278 3232 281 3258
rect 278 3152 281 3168
rect 286 3102 289 3268
rect 270 3072 273 3078
rect 310 3072 313 3238
rect 238 3063 241 3068
rect 286 3062 289 3068
rect 294 3062 297 3068
rect 278 2952 281 2958
rect 214 2912 217 2938
rect 222 2772 225 2848
rect 122 2658 126 2661
rect 62 2572 65 2658
rect 190 2652 193 2658
rect 158 2642 161 2648
rect 62 2552 65 2568
rect 126 2552 129 2558
rect 42 2548 46 2551
rect 102 2542 105 2548
rect 134 2542 137 2548
rect 166 2542 169 2568
rect 190 2552 193 2598
rect 206 2552 209 2668
rect 214 2662 217 2698
rect 222 2662 225 2678
rect 230 2662 233 2938
rect 238 2932 241 2948
rect 238 2921 241 2928
rect 238 2918 249 2921
rect 246 2912 249 2918
rect 238 2892 241 2898
rect 254 2872 257 2938
rect 318 2922 321 3268
rect 346 3258 350 3261
rect 326 3212 329 3258
rect 362 3248 366 3251
rect 374 3242 377 3458
rect 398 3452 401 3458
rect 406 3452 409 3538
rect 422 3522 425 3538
rect 414 3472 417 3478
rect 438 3462 441 3538
rect 454 3512 457 3548
rect 494 3542 497 3548
rect 482 3538 486 3541
rect 462 3472 465 3478
rect 446 3468 454 3471
rect 446 3462 449 3468
rect 470 3462 473 3498
rect 526 3462 529 3528
rect 542 3512 545 3548
rect 566 3522 569 3538
rect 582 3482 585 3538
rect 598 3492 601 3588
rect 610 3548 614 3551
rect 614 3532 617 3538
rect 478 3458 502 3461
rect 538 3458 542 3461
rect 478 3451 481 3458
rect 442 3448 481 3451
rect 422 3442 425 3448
rect 406 3372 409 3388
rect 386 3368 390 3371
rect 390 3302 393 3348
rect 398 3342 401 3348
rect 406 3332 409 3368
rect 422 3342 425 3358
rect 446 3352 449 3358
rect 494 3332 497 3418
rect 506 3368 510 3371
rect 526 3362 529 3458
rect 566 3452 569 3458
rect 574 3442 577 3458
rect 558 3412 561 3418
rect 536 3403 538 3407
rect 542 3403 545 3407
rect 549 3403 552 3407
rect 546 3368 550 3371
rect 514 3358 518 3361
rect 522 3348 526 3351
rect 582 3351 585 3478
rect 622 3472 625 3558
rect 638 3532 641 3658
rect 646 3652 649 3658
rect 654 3632 657 3738
rect 670 3732 673 3738
rect 662 3652 665 3718
rect 670 3652 673 3708
rect 678 3672 681 3738
rect 718 3672 721 3718
rect 726 3702 729 3738
rect 750 3682 753 3758
rect 766 3752 769 3778
rect 774 3772 777 3818
rect 806 3782 809 3818
rect 886 3802 889 4038
rect 894 3952 897 3978
rect 942 3972 945 4018
rect 950 3942 953 3948
rect 902 3882 905 3938
rect 918 3912 921 3938
rect 942 3882 945 3938
rect 958 3912 961 4118
rect 966 4062 969 4068
rect 974 4042 977 4138
rect 1006 4072 1009 4118
rect 982 3972 985 3988
rect 926 3872 929 3878
rect 962 3868 966 3871
rect 982 3851 985 3878
rect 978 3848 985 3851
rect 974 3842 977 3848
rect 922 3838 926 3841
rect 894 3772 897 3788
rect 774 3732 777 3748
rect 758 3672 761 3718
rect 782 3692 785 3748
rect 814 3742 817 3758
rect 798 3732 801 3738
rect 790 3702 793 3718
rect 814 3682 817 3688
rect 822 3682 825 3698
rect 830 3692 833 3747
rect 894 3742 897 3768
rect 902 3742 905 3768
rect 910 3752 913 3798
rect 918 3752 921 3828
rect 934 3812 937 3818
rect 934 3762 937 3798
rect 950 3782 953 3818
rect 966 3762 969 3818
rect 954 3758 958 3761
rect 990 3752 993 4018
rect 998 4012 1001 4058
rect 1006 4052 1009 4058
rect 1014 3971 1017 4058
rect 1022 3992 1025 4008
rect 1014 3968 1022 3971
rect 1038 3961 1041 4118
rect 1048 4103 1050 4107
rect 1054 4103 1057 4107
rect 1061 4103 1064 4107
rect 1086 4072 1089 4138
rect 1054 3992 1057 4068
rect 1062 4062 1065 4068
rect 1126 4062 1129 4068
rect 1142 4062 1145 4088
rect 1154 4068 1158 4071
rect 1154 4058 1158 4061
rect 1130 4048 1145 4051
rect 1122 4018 1129 4021
rect 1098 3968 1102 3971
rect 1030 3958 1041 3961
rect 1126 3962 1129 4018
rect 1142 3992 1145 4048
rect 1166 4022 1169 4118
rect 1182 4092 1185 4148
rect 1174 3982 1177 4018
rect 998 3922 1001 3928
rect 998 3862 1001 3868
rect 1006 3862 1009 3868
rect 1014 3852 1017 3948
rect 1030 3872 1033 3958
rect 1042 3948 1046 3951
rect 1062 3942 1065 3948
rect 1048 3903 1050 3907
rect 1054 3903 1057 3907
rect 1061 3903 1064 3907
rect 1022 3862 1025 3868
rect 1062 3862 1065 3868
rect 998 3792 1001 3848
rect 1030 3832 1033 3858
rect 1054 3852 1057 3858
rect 1010 3758 1014 3761
rect 974 3742 977 3748
rect 982 3742 985 3748
rect 946 3738 950 3741
rect 990 3722 993 3738
rect 862 3692 865 3718
rect 838 3672 841 3688
rect 854 3672 857 3678
rect 686 3642 689 3668
rect 910 3662 913 3668
rect 934 3662 937 3678
rect 950 3662 953 3668
rect 958 3662 961 3718
rect 970 3678 974 3681
rect 714 3658 718 3661
rect 762 3658 766 3661
rect 890 3658 894 3661
rect 978 3658 982 3661
rect 646 3592 649 3618
rect 646 3512 649 3548
rect 654 3532 657 3568
rect 682 3548 686 3551
rect 638 3472 641 3478
rect 646 3472 649 3488
rect 598 3452 601 3458
rect 618 3448 622 3451
rect 654 3442 657 3458
rect 670 3452 673 3458
rect 678 3452 681 3468
rect 686 3442 689 3538
rect 694 3492 697 3558
rect 710 3462 713 3618
rect 654 3422 657 3428
rect 606 3391 609 3418
rect 578 3348 585 3351
rect 598 3388 609 3391
rect 598 3352 601 3388
rect 574 3342 577 3348
rect 514 3338 526 3341
rect 582 3322 585 3338
rect 382 3272 385 3278
rect 342 3202 345 3218
rect 374 3192 377 3228
rect 342 3172 345 3178
rect 326 3162 329 3168
rect 350 3152 353 3188
rect 398 3162 401 3308
rect 414 3282 417 3288
rect 346 3148 350 3151
rect 326 3138 334 3141
rect 326 3062 329 3138
rect 358 3122 361 3158
rect 422 3152 425 3298
rect 598 3292 601 3338
rect 494 3272 497 3288
rect 598 3272 601 3278
rect 522 3258 526 3261
rect 430 3192 433 3258
rect 578 3238 582 3241
rect 478 3212 481 3218
rect 454 3182 457 3208
rect 454 3172 457 3178
rect 470 3152 473 3158
rect 526 3152 529 3228
rect 536 3203 538 3207
rect 542 3203 545 3207
rect 549 3203 552 3207
rect 566 3162 569 3168
rect 490 3148 494 3151
rect 390 3132 393 3148
rect 526 3142 529 3148
rect 410 3138 414 3141
rect 482 3138 486 3141
rect 382 3072 385 3128
rect 390 3092 393 3118
rect 406 3112 409 3118
rect 422 3102 425 3138
rect 338 3058 342 3061
rect 326 3042 329 3058
rect 334 2981 337 3018
rect 342 2992 345 3058
rect 374 3052 377 3058
rect 390 3052 393 3078
rect 414 3072 417 3098
rect 418 3068 422 3071
rect 418 3058 422 3061
rect 406 3052 409 3058
rect 358 3032 361 3038
rect 326 2978 337 2981
rect 326 2892 329 2978
rect 338 2968 342 2971
rect 358 2952 361 2988
rect 390 2972 393 3018
rect 406 2972 409 3048
rect 430 3032 433 3058
rect 398 2968 406 2971
rect 390 2962 393 2968
rect 370 2958 374 2961
rect 362 2938 366 2941
rect 334 2928 342 2931
rect 334 2892 337 2928
rect 342 2918 350 2921
rect 342 2902 345 2918
rect 342 2872 345 2898
rect 398 2882 401 2968
rect 406 2952 409 2968
rect 430 2952 433 2978
rect 454 2952 457 3068
rect 462 3062 465 3078
rect 470 3062 473 3128
rect 470 2952 473 2958
rect 418 2938 422 2941
rect 462 2932 465 2948
rect 478 2941 481 3118
rect 486 3072 489 3138
rect 502 3082 505 3128
rect 518 3092 521 3118
rect 486 2972 489 3018
rect 486 2952 489 2968
rect 494 2962 497 2968
rect 518 2962 521 2968
rect 526 2961 529 3108
rect 550 3102 553 3148
rect 582 3132 585 3148
rect 598 3122 601 3268
rect 606 3262 609 3298
rect 622 3292 625 3348
rect 630 3302 633 3418
rect 694 3382 697 3448
rect 726 3431 729 3578
rect 734 3552 737 3558
rect 798 3552 801 3578
rect 834 3548 838 3551
rect 758 3472 761 3548
rect 806 3542 809 3548
rect 846 3542 849 3658
rect 878 3652 881 3658
rect 942 3652 945 3658
rect 990 3652 993 3658
rect 894 3632 897 3648
rect 790 3512 793 3518
rect 718 3428 729 3431
rect 734 3432 737 3458
rect 742 3452 745 3458
rect 710 3372 713 3378
rect 662 3362 665 3368
rect 690 3348 694 3351
rect 646 3342 649 3348
rect 614 3262 617 3268
rect 646 3262 649 3338
rect 678 3322 681 3328
rect 686 3312 689 3338
rect 654 3282 657 3308
rect 682 3288 686 3291
rect 710 3282 713 3328
rect 718 3292 721 3428
rect 726 3402 729 3418
rect 746 3378 750 3381
rect 782 3362 785 3468
rect 798 3462 801 3528
rect 806 3372 809 3538
rect 870 3532 873 3628
rect 878 3562 881 3568
rect 902 3562 905 3618
rect 918 3572 921 3618
rect 926 3562 929 3648
rect 998 3642 1001 3748
rect 1022 3742 1025 3768
rect 1062 3762 1065 3848
rect 1070 3842 1073 3948
rect 1110 3942 1113 3948
rect 1078 3912 1081 3938
rect 1094 3932 1097 3938
rect 1102 3932 1105 3938
rect 1118 3912 1121 3948
rect 1106 3888 1110 3891
rect 1118 3882 1121 3888
rect 1126 3882 1129 3958
rect 1142 3952 1145 3968
rect 1150 3902 1153 3978
rect 1182 3972 1185 4088
rect 1190 4072 1193 4178
rect 1198 4162 1201 4168
rect 1206 4162 1209 4238
rect 1214 4152 1217 4328
rect 1222 4282 1225 4328
rect 1230 4292 1233 4318
rect 1246 4312 1249 4338
rect 1222 4262 1225 4278
rect 1262 4272 1265 4278
rect 1222 4242 1225 4248
rect 1222 4172 1225 4188
rect 1222 4152 1225 4158
rect 1222 4132 1225 4138
rect 1170 3968 1174 3971
rect 1158 3962 1161 3968
rect 1142 3882 1145 3888
rect 1150 3881 1153 3898
rect 1146 3878 1153 3881
rect 1158 3882 1161 3938
rect 1174 3932 1177 3938
rect 1166 3872 1169 3878
rect 1182 3872 1185 3958
rect 1190 3952 1193 4058
rect 1214 4052 1217 4118
rect 1230 4092 1233 4208
rect 1246 4152 1249 4258
rect 1246 4132 1249 4148
rect 1254 4142 1257 4268
rect 1278 4162 1281 4678
rect 1286 4562 1289 4738
rect 1326 4732 1329 4808
rect 1334 4792 1337 4858
rect 1358 4752 1361 4758
rect 1374 4752 1377 4858
rect 1414 4812 1417 4818
rect 1350 4742 1353 4748
rect 1374 4742 1377 4748
rect 1398 4742 1401 4748
rect 1302 4702 1305 4718
rect 1302 4672 1305 4678
rect 1318 4671 1321 4718
rect 1334 4682 1337 4688
rect 1318 4668 1329 4671
rect 1314 4658 1318 4661
rect 1286 4542 1289 4558
rect 1294 4542 1297 4548
rect 1286 4292 1289 4358
rect 1294 4352 1297 4458
rect 1302 4421 1305 4658
rect 1326 4652 1329 4668
rect 1350 4621 1353 4738
rect 1374 4672 1377 4738
rect 1374 4662 1377 4668
rect 1386 4658 1390 4661
rect 1350 4618 1361 4621
rect 1310 4502 1313 4618
rect 1358 4552 1361 4618
rect 1414 4582 1417 4808
rect 1422 4762 1425 4818
rect 1502 4772 1505 4868
rect 1518 4841 1521 4868
rect 1598 4862 1601 4868
rect 1510 4838 1521 4841
rect 1538 4858 1542 4861
rect 1498 4748 1502 4751
rect 1454 4702 1457 4718
rect 1430 4682 1433 4688
rect 1470 4672 1473 4678
rect 1454 4662 1457 4668
rect 1446 4652 1449 4658
rect 1430 4642 1433 4648
rect 1422 4572 1425 4638
rect 1446 4592 1449 4638
rect 1346 4548 1350 4551
rect 1378 4548 1382 4551
rect 1450 4548 1454 4551
rect 1358 4542 1361 4548
rect 1470 4542 1473 4668
rect 1498 4658 1502 4661
rect 1510 4622 1513 4838
rect 1526 4792 1529 4858
rect 1542 4782 1545 4848
rect 1622 4832 1625 4858
rect 1654 4812 1657 4818
rect 1560 4803 1562 4807
rect 1566 4803 1569 4807
rect 1573 4803 1576 4807
rect 1554 4768 1558 4771
rect 1518 4752 1521 4768
rect 1566 4752 1569 4778
rect 1606 4762 1609 4768
rect 1626 4758 1638 4761
rect 1498 4548 1502 4551
rect 1370 4538 1374 4541
rect 1402 4538 1406 4541
rect 1450 4538 1454 4541
rect 1342 4512 1345 4518
rect 1346 4478 1350 4481
rect 1358 4472 1361 4538
rect 1398 4512 1401 4528
rect 1414 4442 1417 4518
rect 1422 4472 1425 4478
rect 1438 4462 1441 4498
rect 1510 4472 1513 4478
rect 1498 4468 1502 4471
rect 1430 4452 1433 4458
rect 1494 4452 1497 4458
rect 1478 4442 1481 4448
rect 1302 4418 1313 4421
rect 1294 4342 1297 4348
rect 1310 4272 1313 4418
rect 1334 4392 1337 4408
rect 1366 4392 1369 4418
rect 1334 4352 1337 4358
rect 1318 4318 1326 4321
rect 1306 4268 1310 4271
rect 1318 4262 1321 4318
rect 1326 4262 1329 4268
rect 1286 4252 1289 4258
rect 1262 4122 1265 4138
rect 1294 4122 1297 4258
rect 1314 4248 1318 4251
rect 1326 4212 1329 4258
rect 1334 4191 1337 4348
rect 1366 4342 1369 4348
rect 1390 4342 1393 4348
rect 1346 4328 1350 4331
rect 1342 4282 1345 4288
rect 1358 4192 1361 4268
rect 1374 4192 1377 4298
rect 1382 4272 1385 4328
rect 1454 4322 1457 4418
rect 1470 4372 1473 4378
rect 1486 4362 1489 4368
rect 1434 4288 1438 4291
rect 1382 4252 1385 4258
rect 1334 4188 1345 4191
rect 1330 4178 1334 4181
rect 1342 4152 1345 4188
rect 1382 4152 1385 4238
rect 1406 4162 1409 4288
rect 1446 4282 1449 4318
rect 1470 4302 1473 4348
rect 1478 4342 1481 4358
rect 1502 4352 1505 4458
rect 1486 4342 1489 4348
rect 1498 4258 1502 4261
rect 1510 4261 1513 4388
rect 1518 4342 1521 4728
rect 1558 4632 1561 4668
rect 1558 4622 1561 4628
rect 1566 4622 1569 4718
rect 1574 4682 1577 4758
rect 1594 4748 1598 4751
rect 1634 4748 1638 4751
rect 1622 4742 1625 4748
rect 1662 4742 1665 4868
rect 1758 4863 1761 4868
rect 1674 4858 1678 4861
rect 1790 4862 1793 4868
rect 1670 4772 1673 4808
rect 1686 4792 1689 4848
rect 1790 4842 1793 4848
rect 1694 4812 1697 4818
rect 1702 4762 1705 4838
rect 1710 4832 1713 4838
rect 1674 4748 1678 4751
rect 1702 4742 1705 4748
rect 1634 4738 1638 4741
rect 1598 4722 1601 4738
rect 1606 4692 1609 4738
rect 1662 4732 1665 4738
rect 1638 4682 1641 4698
rect 1650 4678 1654 4681
rect 1594 4658 1598 4661
rect 1582 4652 1585 4658
rect 1622 4652 1625 4658
rect 1598 4631 1601 4648
rect 1606 4642 1609 4648
rect 1598 4628 1609 4631
rect 1550 4592 1553 4618
rect 1560 4603 1562 4607
rect 1566 4603 1569 4607
rect 1573 4603 1576 4607
rect 1582 4532 1585 4618
rect 1606 4592 1609 4628
rect 1590 4572 1593 4588
rect 1622 4552 1625 4628
rect 1602 4548 1606 4551
rect 1630 4542 1633 4588
rect 1638 4542 1641 4548
rect 1614 4532 1617 4538
rect 1602 4528 1609 4531
rect 1550 4512 1553 4518
rect 1558 4472 1561 4518
rect 1606 4492 1609 4528
rect 1594 4468 1598 4471
rect 1614 4452 1617 4518
rect 1622 4472 1625 4478
rect 1622 4452 1625 4458
rect 1566 4422 1569 4428
rect 1560 4403 1562 4407
rect 1566 4403 1569 4407
rect 1573 4403 1576 4407
rect 1582 4342 1585 4418
rect 1598 4342 1601 4347
rect 1534 4322 1537 4328
rect 1574 4272 1577 4308
rect 1510 4258 1518 4261
rect 1286 4102 1289 4118
rect 1302 4112 1305 4148
rect 1310 4142 1313 4148
rect 1358 4142 1361 4148
rect 1322 4128 1326 4131
rect 1362 4128 1366 4131
rect 1222 4082 1225 4088
rect 1310 4072 1313 4108
rect 1262 4062 1265 4068
rect 1250 4058 1254 4061
rect 1198 3992 1201 4018
rect 1230 4012 1233 4018
rect 1238 3992 1241 4048
rect 1198 3962 1201 3968
rect 1214 3962 1217 3968
rect 1198 3952 1201 3958
rect 1206 3942 1209 3958
rect 1230 3952 1233 3978
rect 1246 3962 1249 4058
rect 1294 4042 1297 4059
rect 1254 4032 1257 4038
rect 1278 3992 1281 3998
rect 1254 3982 1257 3988
rect 1190 3892 1193 3938
rect 1198 3882 1201 3888
rect 1142 3862 1145 3868
rect 1090 3858 1094 3861
rect 1106 3858 1110 3861
rect 1006 3682 1009 3688
rect 1014 3662 1017 3718
rect 1030 3702 1033 3748
rect 1022 3662 1025 3688
rect 1038 3672 1041 3738
rect 1070 3712 1073 3738
rect 1048 3703 1050 3707
rect 1054 3703 1057 3707
rect 1061 3703 1064 3707
rect 1078 3672 1081 3818
rect 1094 3742 1097 3808
rect 1102 3752 1105 3768
rect 1110 3722 1113 3858
rect 1134 3762 1137 3818
rect 1142 3802 1145 3858
rect 1122 3758 1126 3761
rect 1150 3752 1153 3838
rect 1158 3792 1161 3848
rect 1166 3812 1169 3858
rect 1174 3842 1177 3858
rect 1206 3852 1209 3938
rect 1190 3791 1193 3838
rect 1214 3812 1217 3918
rect 1186 3788 1193 3791
rect 1126 3722 1129 3748
rect 1142 3732 1145 3738
rect 1118 3702 1121 3718
rect 1102 3672 1105 3678
rect 1094 3662 1097 3668
rect 1126 3662 1129 3668
rect 1134 3662 1137 3718
rect 1150 3662 1153 3748
rect 1174 3742 1177 3748
rect 1230 3732 1233 3948
rect 1238 3922 1241 3938
rect 1262 3932 1265 3938
rect 1238 3752 1241 3888
rect 1246 3742 1249 3868
rect 1262 3863 1265 3888
rect 1278 3872 1281 3938
rect 1294 3882 1297 4018
rect 1310 3992 1313 4038
rect 1322 3948 1326 3951
rect 1302 3942 1305 3948
rect 1302 3872 1305 3938
rect 1310 3882 1313 3898
rect 1318 3892 1321 3908
rect 1342 3902 1345 4128
rect 1382 4122 1385 4148
rect 1422 4142 1425 4238
rect 1394 4138 1398 4141
rect 1386 4088 1390 4091
rect 1370 4068 1374 4071
rect 1382 4042 1385 4078
rect 1398 4062 1401 4118
rect 1406 4091 1409 4118
rect 1422 4112 1425 4138
rect 1406 4088 1417 4091
rect 1406 4072 1409 4078
rect 1414 4072 1417 4088
rect 1438 4082 1441 4258
rect 1454 4162 1457 4218
rect 1450 4148 1454 4151
rect 1410 4058 1414 4061
rect 1430 4052 1433 4068
rect 1462 4062 1465 4098
rect 1494 4072 1497 4158
rect 1510 4132 1513 4138
rect 1506 4118 1510 4121
rect 1518 4082 1521 4258
rect 1550 4242 1553 4248
rect 1574 4222 1577 4268
rect 1582 4262 1585 4288
rect 1614 4282 1617 4448
rect 1630 4352 1633 4538
rect 1646 4492 1649 4618
rect 1654 4512 1657 4528
rect 1646 4462 1649 4468
rect 1642 4448 1646 4451
rect 1642 4348 1646 4351
rect 1650 4338 1654 4341
rect 1630 4332 1633 4338
rect 1590 4262 1593 4268
rect 1610 4248 1614 4251
rect 1560 4203 1562 4207
rect 1566 4203 1569 4207
rect 1573 4203 1576 4207
rect 1526 4162 1529 4168
rect 1526 4142 1529 4148
rect 1518 4062 1521 4068
rect 1490 4058 1494 4061
rect 1326 3852 1329 3858
rect 1334 3852 1337 3878
rect 1350 3862 1353 3908
rect 1366 3902 1369 3948
rect 1390 3942 1393 3948
rect 1370 3888 1374 3891
rect 1390 3872 1393 3928
rect 1398 3892 1401 3898
rect 1362 3868 1366 3871
rect 1358 3862 1361 3868
rect 1362 3848 1366 3851
rect 1350 3842 1353 3848
rect 1302 3782 1305 3818
rect 1326 3762 1329 3768
rect 1298 3758 1302 3761
rect 1306 3748 1310 3751
rect 1306 3738 1310 3741
rect 1166 3672 1169 3678
rect 1034 3658 1038 3661
rect 1114 3658 1118 3661
rect 1150 3652 1153 3658
rect 1082 3648 1086 3651
rect 1186 3648 1190 3651
rect 934 3592 937 3628
rect 902 3552 905 3558
rect 882 3548 886 3551
rect 818 3528 822 3531
rect 846 3492 849 3528
rect 854 3512 857 3528
rect 862 3512 865 3518
rect 842 3488 846 3491
rect 870 3472 873 3528
rect 846 3462 849 3468
rect 862 3462 865 3468
rect 842 3448 846 3451
rect 782 3352 785 3358
rect 802 3348 806 3351
rect 726 3342 729 3348
rect 734 3301 737 3348
rect 746 3338 750 3341
rect 730 3298 737 3301
rect 654 3272 657 3278
rect 670 3262 673 3268
rect 698 3258 702 3261
rect 630 3242 633 3248
rect 646 3172 649 3258
rect 662 3252 665 3258
rect 634 3148 638 3151
rect 614 3112 617 3128
rect 550 3091 553 3098
rect 550 3088 561 3091
rect 542 3063 545 3088
rect 536 3003 538 3007
rect 542 3003 545 3007
rect 549 3003 552 3007
rect 558 2992 561 3088
rect 574 3062 577 3108
rect 606 3082 609 3088
rect 566 2972 569 2978
rect 574 2962 577 3058
rect 526 2958 534 2961
rect 474 2938 481 2941
rect 414 2882 417 2918
rect 362 2868 366 2871
rect 394 2868 398 2871
rect 254 2852 257 2868
rect 278 2862 281 2868
rect 350 2842 353 2858
rect 374 2842 377 2848
rect 414 2792 417 2858
rect 430 2852 433 2868
rect 242 2768 246 2771
rect 238 2748 246 2751
rect 238 2672 241 2748
rect 246 2692 249 2738
rect 262 2732 265 2768
rect 366 2762 369 2768
rect 254 2682 257 2718
rect 278 2692 281 2748
rect 298 2747 302 2750
rect 426 2748 430 2751
rect 326 2742 329 2748
rect 382 2742 385 2748
rect 398 2742 401 2748
rect 310 2682 313 2718
rect 238 2662 241 2668
rect 262 2662 265 2668
rect 270 2662 273 2668
rect 230 2652 233 2658
rect 250 2588 254 2591
rect 294 2582 297 2658
rect 318 2592 321 2678
rect 274 2548 278 2551
rect 106 2528 110 2531
rect 98 2518 102 2521
rect 134 2512 137 2538
rect 142 2532 145 2538
rect 150 2522 153 2528
rect 150 2502 153 2518
rect 146 2488 150 2491
rect 10 2468 14 2471
rect 22 2462 25 2488
rect 30 2452 33 2468
rect 114 2459 118 2462
rect 134 2462 137 2468
rect 182 2462 185 2468
rect 6 2372 9 2378
rect 10 2288 14 2291
rect 62 2272 65 2348
rect 86 2342 89 2458
rect 206 2392 209 2548
rect 294 2542 297 2568
rect 318 2542 321 2548
rect 326 2542 329 2738
rect 354 2718 358 2721
rect 374 2692 377 2718
rect 398 2682 401 2738
rect 446 2702 449 2918
rect 458 2858 462 2861
rect 354 2668 358 2671
rect 334 2662 337 2668
rect 366 2662 369 2668
rect 406 2662 409 2668
rect 246 2492 249 2508
rect 254 2492 257 2528
rect 214 2432 217 2459
rect 230 2452 233 2468
rect 246 2462 249 2488
rect 262 2462 265 2518
rect 270 2492 273 2538
rect 334 2492 337 2658
rect 342 2602 345 2618
rect 382 2552 385 2558
rect 390 2542 393 2578
rect 430 2552 433 2578
rect 438 2552 441 2618
rect 470 2562 473 2688
rect 478 2662 481 2938
rect 494 2862 497 2918
rect 502 2891 505 2958
rect 514 2948 518 2951
rect 526 2932 529 2938
rect 502 2888 510 2891
rect 558 2872 561 2958
rect 566 2942 569 2948
rect 574 2902 577 2938
rect 582 2912 585 2948
rect 606 2942 609 3038
rect 614 3022 617 3078
rect 630 3052 633 3078
rect 650 3068 654 3071
rect 670 3062 673 3218
rect 690 3158 697 3161
rect 686 3142 689 3148
rect 682 3118 686 3121
rect 694 3092 697 3158
rect 702 3152 705 3228
rect 710 3161 713 3278
rect 718 3272 721 3288
rect 726 3262 729 3298
rect 782 3272 785 3348
rect 830 3272 833 3448
rect 838 3371 841 3388
rect 870 3372 873 3468
rect 878 3382 881 3548
rect 918 3542 921 3558
rect 838 3368 849 3371
rect 846 3362 849 3368
rect 878 3342 881 3358
rect 898 3348 902 3351
rect 862 3332 865 3338
rect 854 3272 857 3318
rect 870 3272 873 3278
rect 738 3268 742 3271
rect 774 3263 777 3268
rect 850 3258 854 3261
rect 742 3252 745 3258
rect 734 3162 737 3238
rect 710 3158 718 3161
rect 774 3152 777 3158
rect 798 3152 801 3188
rect 862 3172 865 3258
rect 878 3252 881 3268
rect 902 3262 905 3288
rect 910 3272 913 3518
rect 918 3332 921 3538
rect 926 3482 929 3558
rect 934 3472 937 3548
rect 942 3522 945 3538
rect 950 3502 953 3548
rect 970 3518 974 3521
rect 982 3492 985 3538
rect 990 3532 993 3538
rect 942 3452 945 3488
rect 990 3472 993 3508
rect 958 3462 961 3468
rect 1006 3462 1009 3588
rect 994 3458 998 3461
rect 982 3402 985 3418
rect 958 3372 961 3378
rect 966 3352 969 3398
rect 926 3292 929 3348
rect 934 3282 937 3298
rect 950 3282 953 3288
rect 966 3272 969 3348
rect 982 3332 985 3368
rect 998 3342 1001 3358
rect 974 3302 977 3318
rect 982 3282 985 3318
rect 982 3272 985 3278
rect 922 3268 926 3271
rect 890 3258 894 3261
rect 886 3192 889 3248
rect 834 3158 838 3161
rect 702 3142 705 3148
rect 806 3142 809 3148
rect 814 3142 817 3158
rect 738 3138 742 3141
rect 762 3138 766 3141
rect 678 3072 681 3078
rect 702 3072 705 3088
rect 710 3082 713 3118
rect 718 3092 721 3138
rect 838 3132 841 3148
rect 786 3118 790 3121
rect 726 3092 729 3118
rect 730 3078 734 3081
rect 690 3048 694 3051
rect 622 3032 625 3038
rect 670 2962 673 3018
rect 662 2951 665 2958
rect 686 2952 689 2958
rect 662 2948 670 2951
rect 598 2872 601 2918
rect 638 2902 641 2948
rect 678 2942 681 2948
rect 718 2942 721 3018
rect 726 2958 734 2961
rect 726 2952 729 2958
rect 734 2942 737 2948
rect 654 2932 657 2938
rect 646 2921 649 2928
rect 646 2918 657 2921
rect 654 2892 657 2918
rect 642 2888 646 2891
rect 494 2842 497 2848
rect 490 2758 494 2761
rect 494 2748 502 2751
rect 514 2748 518 2751
rect 494 2662 497 2748
rect 494 2652 497 2658
rect 398 2542 401 2548
rect 478 2542 481 2618
rect 486 2562 489 2568
rect 494 2552 497 2568
rect 502 2562 505 2718
rect 514 2668 518 2671
rect 526 2671 529 2868
rect 538 2858 542 2861
rect 558 2852 561 2868
rect 586 2858 590 2861
rect 536 2803 538 2807
rect 542 2803 545 2807
rect 549 2803 552 2807
rect 646 2802 649 2878
rect 662 2862 665 2938
rect 678 2892 681 2928
rect 702 2892 705 2918
rect 670 2882 673 2888
rect 702 2862 705 2868
rect 606 2792 609 2798
rect 662 2782 665 2858
rect 694 2842 697 2858
rect 694 2832 697 2838
rect 542 2692 545 2758
rect 550 2742 553 2758
rect 562 2748 566 2751
rect 582 2742 585 2768
rect 658 2748 662 2751
rect 574 2722 577 2728
rect 582 2712 585 2738
rect 578 2688 582 2691
rect 526 2668 534 2671
rect 522 2648 526 2651
rect 534 2632 537 2668
rect 536 2603 538 2607
rect 542 2603 545 2607
rect 549 2603 552 2607
rect 530 2568 534 2571
rect 490 2538 494 2541
rect 514 2538 518 2541
rect 414 2522 417 2528
rect 378 2518 382 2521
rect 374 2482 377 2488
rect 310 2462 313 2468
rect 302 2452 305 2458
rect 94 2351 97 2358
rect 126 2342 129 2388
rect 166 2362 169 2368
rect 182 2362 185 2368
rect 154 2358 158 2361
rect 154 2348 158 2351
rect 214 2351 217 2358
rect 134 2331 137 2348
rect 126 2328 137 2331
rect 62 2152 65 2268
rect 70 2263 73 2278
rect 118 2272 121 2278
rect 106 2268 110 2271
rect 126 2262 129 2328
rect 134 2292 137 2308
rect 110 2162 113 2258
rect 134 2252 137 2288
rect 158 2272 161 2338
rect 166 2272 169 2348
rect 230 2342 233 2448
rect 274 2368 278 2371
rect 286 2352 289 2448
rect 318 2352 321 2368
rect 326 2352 329 2358
rect 342 2352 345 2418
rect 358 2362 361 2368
rect 366 2361 369 2478
rect 382 2462 385 2468
rect 398 2452 401 2468
rect 422 2462 425 2508
rect 446 2492 449 2538
rect 466 2528 470 2531
rect 454 2512 457 2518
rect 494 2492 497 2528
rect 502 2462 505 2488
rect 534 2482 537 2548
rect 558 2542 561 2648
rect 574 2642 577 2668
rect 606 2592 609 2618
rect 574 2552 577 2558
rect 582 2552 585 2568
rect 622 2562 625 2588
rect 638 2551 641 2748
rect 710 2742 713 2848
rect 718 2832 721 2848
rect 650 2738 654 2741
rect 646 2682 649 2738
rect 702 2692 705 2698
rect 646 2652 649 2659
rect 638 2548 646 2551
rect 566 2512 569 2518
rect 590 2482 593 2548
rect 638 2542 641 2548
rect 502 2442 505 2458
rect 478 2392 481 2418
rect 378 2368 382 2371
rect 490 2368 494 2371
rect 366 2358 377 2361
rect 374 2352 377 2358
rect 306 2318 310 2321
rect 290 2288 294 2291
rect 6 2142 9 2148
rect 10 2088 14 2091
rect 62 1992 65 2148
rect 90 2147 94 2150
rect 118 2092 121 2118
rect 150 2082 153 2188
rect 158 2182 161 2268
rect 166 2262 169 2268
rect 190 2241 193 2258
rect 230 2252 233 2258
rect 190 2238 201 2241
rect 198 2232 201 2238
rect 162 2148 166 2151
rect 182 2132 185 2138
rect 158 2082 161 2088
rect 70 2063 73 2078
rect 114 2068 118 2071
rect 86 2012 89 2068
rect 134 2062 137 2068
rect 166 2061 169 2098
rect 178 2068 182 2071
rect 166 2058 174 2061
rect 102 2052 105 2058
rect 182 2052 185 2068
rect 190 2052 193 2078
rect 158 2042 161 2048
rect 198 2031 201 2228
rect 254 2221 257 2258
rect 254 2218 265 2221
rect 218 2168 222 2171
rect 250 2168 254 2171
rect 230 2152 233 2158
rect 242 2148 246 2151
rect 214 2072 217 2108
rect 222 2092 225 2138
rect 230 2112 233 2148
rect 234 2088 238 2091
rect 226 2078 230 2081
rect 206 2042 209 2048
rect 198 2028 209 2031
rect 134 1992 137 2008
rect 182 1952 185 1978
rect 10 1938 14 1941
rect 74 1938 78 1941
rect 6 1882 9 1888
rect 14 1861 17 1938
rect 6 1858 17 1861
rect 6 1832 9 1858
rect 6 1742 9 1828
rect 62 1792 65 1868
rect 102 1862 105 1868
rect 118 1862 121 1948
rect 70 1852 73 1859
rect 106 1848 110 1851
rect 126 1842 129 1868
rect 134 1852 137 1878
rect 158 1872 161 1898
rect 174 1882 177 1888
rect 166 1872 169 1878
rect 154 1858 158 1861
rect 142 1852 145 1858
rect 166 1792 169 1798
rect 86 1742 89 1748
rect 66 1738 70 1741
rect 6 1672 9 1738
rect 102 1711 105 1747
rect 182 1742 185 1938
rect 190 1862 193 1868
rect 198 1752 201 1938
rect 206 1862 209 2028
rect 222 1922 225 2058
rect 238 1962 241 1968
rect 246 1952 249 2108
rect 262 2072 265 2218
rect 270 2152 273 2258
rect 294 2212 297 2268
rect 302 2262 305 2268
rect 326 2252 329 2288
rect 302 2242 305 2248
rect 278 2142 281 2178
rect 310 2142 313 2147
rect 334 2142 337 2338
rect 342 2272 345 2348
rect 350 2282 353 2348
rect 366 2342 369 2348
rect 374 2331 377 2348
rect 366 2328 377 2331
rect 358 2302 361 2318
rect 350 2272 353 2278
rect 366 2262 369 2328
rect 390 2302 393 2358
rect 430 2352 433 2368
rect 478 2361 481 2368
rect 478 2358 502 2361
rect 502 2342 505 2348
rect 490 2338 494 2341
rect 406 2322 409 2338
rect 382 2263 385 2298
rect 406 2272 409 2318
rect 510 2312 513 2478
rect 542 2462 545 2478
rect 590 2462 593 2468
rect 530 2458 534 2461
rect 554 2458 561 2461
rect 536 2403 538 2407
rect 542 2403 545 2407
rect 549 2403 552 2407
rect 558 2382 561 2458
rect 602 2458 606 2461
rect 574 2452 577 2458
rect 602 2448 606 2451
rect 566 2382 569 2418
rect 530 2368 534 2371
rect 446 2292 449 2298
rect 454 2282 457 2288
rect 470 2282 473 2298
rect 502 2292 505 2298
rect 478 2282 481 2288
rect 514 2268 518 2271
rect 346 2258 350 2261
rect 370 2188 374 2191
rect 390 2142 393 2268
rect 470 2262 473 2268
rect 526 2262 529 2338
rect 542 2292 545 2378
rect 574 2352 577 2368
rect 550 2348 558 2351
rect 550 2302 553 2348
rect 558 2338 566 2341
rect 486 2232 489 2258
rect 542 2232 545 2248
rect 536 2203 538 2207
rect 542 2203 545 2207
rect 549 2203 552 2207
rect 410 2148 414 2151
rect 262 2012 265 2068
rect 270 2042 273 2058
rect 254 1982 257 1988
rect 278 1982 281 2138
rect 294 2132 297 2138
rect 370 2128 374 2131
rect 278 1962 281 1968
rect 294 1952 297 2118
rect 326 2082 329 2088
rect 390 2072 393 2138
rect 422 2092 425 2188
rect 462 2072 465 2178
rect 474 2168 478 2171
rect 510 2162 513 2168
rect 498 2148 502 2151
rect 478 2112 481 2138
rect 486 2112 489 2148
rect 434 2068 438 2071
rect 342 2012 345 2068
rect 366 2052 369 2058
rect 250 1938 254 1941
rect 222 1872 225 1918
rect 246 1892 249 1928
rect 294 1922 297 1948
rect 302 1942 305 1978
rect 422 1952 425 2058
rect 302 1902 305 1938
rect 342 1932 345 1948
rect 206 1812 209 1858
rect 214 1752 217 1868
rect 222 1862 225 1868
rect 238 1852 241 1868
rect 262 1822 265 1858
rect 270 1852 273 1868
rect 262 1752 265 1758
rect 94 1708 105 1711
rect 6 1601 9 1668
rect 78 1662 81 1698
rect 94 1692 97 1708
rect 126 1682 129 1718
rect 158 1682 161 1738
rect 178 1728 182 1731
rect 166 1712 169 1718
rect 90 1668 94 1671
rect 110 1662 113 1668
rect 182 1662 185 1718
rect 190 1692 193 1738
rect 222 1732 225 1738
rect 210 1728 214 1731
rect 222 1692 225 1728
rect 6 1598 17 1601
rect 14 1142 17 1598
rect 62 1552 65 1618
rect 98 1568 102 1571
rect 42 1548 46 1551
rect 62 1532 65 1548
rect 102 1542 105 1548
rect 110 1542 113 1658
rect 190 1621 193 1688
rect 254 1682 257 1728
rect 270 1702 273 1848
rect 258 1678 262 1681
rect 266 1658 270 1661
rect 190 1618 201 1621
rect 122 1548 126 1551
rect 62 1462 65 1528
rect 94 1482 97 1488
rect 102 1472 105 1538
rect 110 1512 113 1538
rect 134 1512 137 1548
rect 150 1532 153 1568
rect 166 1532 169 1538
rect 42 1458 46 1461
rect 122 1458 126 1461
rect 110 1442 113 1458
rect 134 1452 137 1488
rect 166 1482 169 1528
rect 174 1472 177 1508
rect 182 1492 185 1547
rect 190 1482 193 1488
rect 98 1378 102 1381
rect 102 1362 105 1368
rect 50 1348 54 1351
rect 62 1322 65 1348
rect 102 1342 105 1348
rect 62 1262 65 1318
rect 98 1288 102 1291
rect 102 1262 105 1268
rect 110 1262 113 1438
rect 118 1342 121 1348
rect 126 1342 129 1388
rect 134 1372 137 1378
rect 150 1362 153 1458
rect 134 1352 137 1358
rect 150 1352 153 1358
rect 114 1258 121 1261
rect 38 1252 41 1258
rect 62 1192 65 1258
rect 110 1242 113 1248
rect 110 1152 113 1158
rect 10 1138 14 1141
rect 86 1132 89 1138
rect 62 1122 65 1128
rect 38 1062 41 1078
rect 62 1062 65 1118
rect 46 952 49 1058
rect 94 1052 97 1088
rect 102 1062 105 1068
rect 110 1051 113 1068
rect 106 1048 113 1051
rect 118 1062 121 1258
rect 134 1252 137 1288
rect 150 1262 153 1348
rect 158 1272 161 1468
rect 170 1458 174 1461
rect 182 1451 185 1468
rect 174 1448 185 1451
rect 198 1462 201 1618
rect 246 1592 249 1618
rect 254 1492 257 1628
rect 278 1552 281 1818
rect 302 1772 305 1868
rect 310 1862 313 1918
rect 334 1872 337 1928
rect 382 1892 385 1898
rect 370 1888 374 1891
rect 374 1872 377 1878
rect 390 1872 393 1878
rect 398 1872 401 1918
rect 406 1892 409 1928
rect 414 1892 417 1908
rect 402 1858 406 1861
rect 422 1852 425 1888
rect 318 1782 321 1788
rect 326 1752 329 1818
rect 358 1772 361 1778
rect 338 1758 342 1761
rect 326 1702 329 1738
rect 358 1722 361 1768
rect 374 1742 377 1748
rect 382 1742 385 1748
rect 370 1678 374 1681
rect 382 1672 385 1738
rect 398 1682 401 1738
rect 422 1702 425 1838
rect 430 1771 433 2068
rect 442 2058 446 2061
rect 474 2058 481 2061
rect 458 2048 462 2051
rect 438 2042 441 2048
rect 470 2042 473 2048
rect 454 1952 457 2028
rect 470 1952 473 1958
rect 446 1942 449 1948
rect 438 1922 441 1928
rect 446 1892 449 1918
rect 442 1868 446 1871
rect 446 1802 449 1848
rect 454 1842 457 1948
rect 462 1902 465 1938
rect 478 1931 481 2058
rect 486 2052 489 2078
rect 494 2072 497 2138
rect 526 2122 529 2148
rect 558 2142 561 2338
rect 590 2292 593 2318
rect 582 2272 585 2278
rect 566 2262 569 2268
rect 598 2262 601 2398
rect 606 2352 609 2358
rect 614 2352 617 2518
rect 622 2452 625 2498
rect 630 2492 633 2518
rect 638 2472 641 2528
rect 646 2512 649 2518
rect 662 2502 665 2668
rect 686 2662 689 2668
rect 710 2662 713 2688
rect 722 2678 726 2681
rect 734 2672 737 2868
rect 742 2852 745 3118
rect 750 2962 753 2978
rect 758 2962 761 3088
rect 774 3062 777 3098
rect 798 3062 801 3088
rect 822 3052 825 3118
rect 838 3112 841 3128
rect 842 3088 846 3091
rect 854 3062 857 3158
rect 862 3142 865 3168
rect 874 3148 878 3151
rect 894 3132 897 3218
rect 902 3192 905 3258
rect 958 3181 961 3268
rect 1002 3258 1006 3261
rect 966 3252 969 3258
rect 1014 3232 1017 3648
rect 1034 3618 1038 3621
rect 1022 3552 1025 3578
rect 1038 3542 1041 3618
rect 1134 3602 1137 3638
rect 1138 3568 1142 3571
rect 1150 3562 1153 3618
rect 1054 3542 1057 3548
rect 1048 3503 1050 3507
rect 1054 3503 1057 3507
rect 1061 3503 1064 3507
rect 1046 3472 1049 3488
rect 1062 3462 1065 3468
rect 1070 3462 1073 3558
rect 1134 3552 1137 3558
rect 1182 3551 1185 3568
rect 1078 3472 1081 3548
rect 1166 3542 1169 3548
rect 1126 3532 1129 3538
rect 1118 3512 1121 3518
rect 1042 3458 1046 3461
rect 1030 3442 1033 3458
rect 1022 3382 1025 3418
rect 1022 3352 1025 3358
rect 1070 3352 1073 3458
rect 1094 3452 1097 3508
rect 1110 3442 1113 3458
rect 1082 3368 1086 3371
rect 1106 3358 1110 3361
rect 1106 3348 1110 3351
rect 1106 3338 1110 3341
rect 1030 3272 1033 3338
rect 1048 3303 1050 3307
rect 1054 3303 1057 3307
rect 1061 3303 1064 3307
rect 1070 3302 1073 3338
rect 1118 3292 1121 3468
rect 1126 3462 1129 3518
rect 1166 3472 1169 3538
rect 1190 3462 1193 3498
rect 1126 3352 1129 3358
rect 1134 3352 1137 3438
rect 1142 3412 1145 3418
rect 1158 3362 1161 3368
rect 1146 3358 1150 3361
rect 1174 3352 1177 3398
rect 1166 3342 1169 3348
rect 1126 3292 1129 3338
rect 1134 3292 1137 3338
rect 990 3212 993 3228
rect 1054 3182 1057 3258
rect 1078 3192 1081 3268
rect 1142 3252 1145 3258
rect 958 3178 969 3181
rect 902 3162 905 3178
rect 918 3142 921 3158
rect 950 3142 953 3148
rect 862 3072 865 3078
rect 870 3062 873 3068
rect 878 3062 881 3118
rect 886 3102 889 3118
rect 890 3088 894 3091
rect 838 3052 841 3058
rect 830 2992 833 3038
rect 894 3032 897 3078
rect 910 3062 913 3118
rect 934 3072 937 3118
rect 942 3072 945 3078
rect 958 3072 961 3118
rect 954 3058 961 3061
rect 902 2992 905 3058
rect 942 3042 945 3058
rect 958 3032 961 3058
rect 934 3022 937 3028
rect 802 2978 806 2981
rect 778 2958 782 2961
rect 778 2948 782 2951
rect 806 2942 809 2958
rect 910 2952 913 2968
rect 918 2952 921 2978
rect 818 2948 822 2951
rect 882 2948 886 2951
rect 946 2948 950 2951
rect 794 2938 798 2941
rect 782 2932 785 2938
rect 762 2868 766 2871
rect 774 2862 777 2908
rect 806 2892 809 2938
rect 814 2862 817 2948
rect 838 2942 841 2948
rect 926 2932 929 2938
rect 958 2932 961 3018
rect 966 2952 969 3178
rect 1046 3162 1049 3168
rect 1094 3152 1097 3248
rect 1126 3242 1129 3248
rect 1110 3202 1113 3218
rect 994 3148 998 3151
rect 982 3122 985 3128
rect 974 3012 977 3068
rect 982 3062 985 3088
rect 1014 3061 1017 3128
rect 1030 3062 1033 3108
rect 1048 3103 1050 3107
rect 1054 3103 1057 3107
rect 1061 3103 1064 3107
rect 1078 3092 1081 3138
rect 1094 3081 1097 3148
rect 1102 3142 1105 3188
rect 1114 3178 1118 3181
rect 1138 3178 1142 3181
rect 1126 3152 1129 3158
rect 1150 3152 1153 3268
rect 1174 3262 1177 3288
rect 1182 3262 1185 3278
rect 1190 3262 1193 3318
rect 1198 3301 1201 3728
rect 1262 3672 1265 3738
rect 1278 3712 1281 3738
rect 1290 3718 1294 3721
rect 1222 3662 1225 3668
rect 1210 3658 1214 3661
rect 1254 3632 1257 3659
rect 1214 3622 1217 3628
rect 1278 3612 1281 3708
rect 1246 3592 1249 3598
rect 1274 3588 1278 3591
rect 1230 3432 1233 3438
rect 1206 3358 1214 3361
rect 1206 3332 1209 3358
rect 1218 3348 1230 3351
rect 1230 3332 1233 3338
rect 1238 3322 1241 3588
rect 1286 3562 1289 3598
rect 1250 3548 1254 3551
rect 1302 3542 1305 3688
rect 1318 3642 1321 3648
rect 1326 3592 1329 3708
rect 1334 3692 1337 3828
rect 1350 3752 1353 3798
rect 1362 3768 1366 3771
rect 1342 3742 1345 3748
rect 1362 3738 1366 3741
rect 1350 3662 1353 3698
rect 1366 3672 1369 3678
rect 1382 3602 1385 3858
rect 1402 3848 1406 3851
rect 1414 3842 1417 4018
rect 1422 3862 1425 3988
rect 1446 3972 1449 4018
rect 1454 3982 1457 4058
rect 1474 4028 1478 4031
rect 1490 3948 1494 3951
rect 1490 3938 1494 3941
rect 1430 3902 1433 3938
rect 1430 3872 1433 3898
rect 1462 3882 1465 3888
rect 1450 3878 1454 3881
rect 1470 3872 1473 3898
rect 1442 3868 1446 3871
rect 1482 3868 1486 3871
rect 1482 3858 1486 3861
rect 1494 3852 1497 3918
rect 1502 3902 1505 4058
rect 1526 4052 1529 4118
rect 1534 4092 1537 4158
rect 1582 4152 1585 4218
rect 1614 4212 1617 4248
rect 1638 4242 1641 4268
rect 1646 4262 1649 4298
rect 1662 4251 1665 4618
rect 1694 4612 1697 4738
rect 1710 4731 1713 4828
rect 1734 4792 1737 4838
rect 1750 4772 1753 4808
rect 1726 4742 1729 4768
rect 1806 4752 1809 4878
rect 1818 4868 1822 4871
rect 1814 4792 1817 4858
rect 1886 4822 1889 4868
rect 1734 4742 1737 4748
rect 1702 4728 1713 4731
rect 1702 4672 1705 4728
rect 1710 4682 1713 4718
rect 1706 4658 1710 4661
rect 1670 4552 1673 4588
rect 1710 4542 1713 4548
rect 1686 4472 1689 4538
rect 1718 4532 1721 4738
rect 1726 4722 1729 4738
rect 1790 4732 1793 4748
rect 1770 4668 1774 4671
rect 1806 4662 1809 4738
rect 1814 4702 1817 4788
rect 1950 4782 1953 4818
rect 1850 4748 1854 4751
rect 1850 4718 1854 4721
rect 1862 4712 1865 4738
rect 1870 4732 1873 4738
rect 1786 4658 1790 4661
rect 1810 4658 1814 4661
rect 1774 4632 1777 4658
rect 1794 4648 1798 4651
rect 1814 4642 1817 4648
rect 1798 4622 1801 4638
rect 1762 4618 1766 4621
rect 1802 4618 1809 4621
rect 1790 4542 1793 4588
rect 1798 4552 1801 4558
rect 1778 4538 1782 4541
rect 1750 4482 1753 4518
rect 1766 4512 1769 4518
rect 1774 4501 1777 4528
rect 1766 4498 1777 4501
rect 1678 4463 1681 4468
rect 1686 4422 1689 4468
rect 1694 4392 1697 4448
rect 1710 4372 1713 4418
rect 1670 4342 1673 4348
rect 1662 4248 1673 4251
rect 1630 4162 1633 4198
rect 1550 4062 1553 4068
rect 1558 4052 1561 4148
rect 1606 4142 1609 4148
rect 1630 4142 1633 4148
rect 1566 4122 1569 4128
rect 1606 4062 1609 4108
rect 1638 4102 1641 4238
rect 1662 4232 1665 4238
rect 1658 4148 1662 4151
rect 1670 4142 1673 4248
rect 1678 4242 1681 4338
rect 1686 4312 1689 4348
rect 1694 4332 1697 4348
rect 1726 4342 1729 4438
rect 1738 4418 1742 4421
rect 1750 4352 1753 4358
rect 1694 4302 1697 4328
rect 1686 4262 1689 4288
rect 1698 4268 1702 4271
rect 1758 4271 1761 4488
rect 1766 4482 1769 4498
rect 1790 4462 1793 4538
rect 1798 4472 1801 4538
rect 1806 4482 1809 4618
rect 1822 4612 1825 4668
rect 1834 4638 1838 4641
rect 1830 4552 1833 4638
rect 1814 4532 1817 4548
rect 1770 4458 1774 4461
rect 1778 4448 1782 4451
rect 1790 4372 1793 4418
rect 1798 4402 1801 4458
rect 1822 4452 1825 4518
rect 1878 4482 1881 4738
rect 1886 4712 1889 4748
rect 1902 4722 1905 4728
rect 1918 4691 1921 4738
rect 1910 4688 1921 4691
rect 1942 4692 1945 4748
rect 1910 4682 1913 4688
rect 1910 4672 1913 4678
rect 1950 4672 1953 4768
rect 1958 4752 1961 4878
rect 1974 4872 1977 4878
rect 2002 4858 2006 4861
rect 2058 4838 2062 4841
rect 2038 4752 2041 4758
rect 2054 4752 2057 4818
rect 2078 4812 2081 4868
rect 2094 4862 2097 4868
rect 2122 4858 2126 4861
rect 2086 4822 2089 4858
rect 2114 4838 2118 4841
rect 2118 4782 2121 4838
rect 2002 4748 2006 4751
rect 2046 4742 2049 4748
rect 2054 4742 2057 4748
rect 2086 4742 2089 4778
rect 2102 4751 2105 4758
rect 2022 4732 2025 4738
rect 2014 4722 2017 4728
rect 2030 4722 2033 4728
rect 1998 4712 2001 4718
rect 1990 4708 1998 4711
rect 1894 4663 1897 4668
rect 1958 4662 1961 4668
rect 1974 4662 1977 4698
rect 1946 4658 1950 4661
rect 1954 4648 1958 4651
rect 1926 4642 1929 4648
rect 1942 4642 1945 4648
rect 1974 4642 1977 4658
rect 1982 4632 1985 4668
rect 1886 4551 1889 4558
rect 1918 4542 1921 4628
rect 1926 4562 1929 4568
rect 1950 4562 1953 4578
rect 1970 4568 1974 4571
rect 1990 4562 1993 4708
rect 2022 4682 2025 4708
rect 1998 4662 2001 4668
rect 2038 4662 2041 4668
rect 2014 4632 2017 4658
rect 2038 4602 2041 4658
rect 1934 4558 1942 4561
rect 1902 4512 1905 4538
rect 1918 4532 1921 4538
rect 1926 4532 1929 4548
rect 1934 4472 1937 4558
rect 2046 4552 2049 4738
rect 2134 4722 2137 4868
rect 2150 4772 2153 4868
rect 2174 4862 2177 4878
rect 2382 4872 2385 4878
rect 2258 4868 2262 4871
rect 2298 4868 2302 4871
rect 2250 4858 2254 4861
rect 2150 4752 2153 4768
rect 2174 4742 2177 4768
rect 2182 4762 2185 4768
rect 2190 4751 2193 4858
rect 2254 4832 2257 4838
rect 2230 4792 2233 4818
rect 2202 4768 2206 4771
rect 2202 4758 2206 4761
rect 2226 4758 2230 4761
rect 2186 4748 2193 4751
rect 2166 4722 2169 4728
rect 2072 4703 2074 4707
rect 2078 4703 2081 4707
rect 2085 4703 2088 4707
rect 2102 4692 2105 4718
rect 2174 4712 2177 4738
rect 2222 4721 2225 4748
rect 2246 4742 2249 4748
rect 2262 4742 2265 4868
rect 2270 4842 2273 4848
rect 2230 4732 2233 4738
rect 2214 4718 2225 4721
rect 2214 4702 2217 4718
rect 2058 4688 2062 4691
rect 2134 4672 2137 4678
rect 2058 4668 2062 4671
rect 2158 4662 2161 4678
rect 2074 4658 2078 4661
rect 2118 4652 2121 4658
rect 2214 4642 2217 4698
rect 2238 4682 2241 4688
rect 2234 4668 2238 4671
rect 2102 4612 2105 4618
rect 2086 4562 2089 4568
rect 2030 4542 2033 4548
rect 2126 4542 2129 4548
rect 1978 4538 1982 4541
rect 2098 4538 2102 4541
rect 1966 4532 1969 4538
rect 2114 4528 2118 4531
rect 1842 4468 1846 4471
rect 1922 4468 1926 4471
rect 1846 4452 1849 4458
rect 1834 4448 1838 4451
rect 1822 4432 1825 4448
rect 1854 4442 1857 4458
rect 1910 4452 1913 4458
rect 1890 4448 1894 4451
rect 1930 4438 1934 4441
rect 1814 4382 1817 4418
rect 1810 4368 1814 4371
rect 1822 4352 1825 4378
rect 1846 4362 1849 4368
rect 1834 4348 1838 4351
rect 1766 4302 1769 4338
rect 1766 4282 1769 4298
rect 1798 4282 1801 4288
rect 1758 4268 1769 4271
rect 1690 4258 1694 4261
rect 1758 4252 1761 4258
rect 1690 4248 1694 4251
rect 1698 4228 1702 4231
rect 1710 4162 1713 4168
rect 1726 4162 1729 4198
rect 1734 4162 1737 4208
rect 1686 4152 1689 4158
rect 1714 4148 1718 4151
rect 1646 4092 1649 4138
rect 1694 4132 1697 4148
rect 1702 4142 1705 4148
rect 1750 4132 1753 4138
rect 1758 4122 1761 4128
rect 1670 4112 1673 4118
rect 1742 4102 1745 4118
rect 1630 4072 1633 4078
rect 1538 4048 1542 4051
rect 1534 3992 1537 4048
rect 1566 4032 1569 4058
rect 1614 4052 1617 4058
rect 1560 4003 1562 4007
rect 1566 4003 1569 4007
rect 1573 4003 1576 4007
rect 1598 3992 1601 4018
rect 1654 3992 1657 4058
rect 1538 3978 1542 3981
rect 1606 3972 1609 3978
rect 1542 3962 1545 3968
rect 1582 3942 1585 3948
rect 1562 3938 1566 3941
rect 1590 3922 1593 3948
rect 1618 3938 1622 3941
rect 1546 3918 1550 3921
rect 1590 3912 1593 3918
rect 1638 3912 1641 3938
rect 1646 3932 1649 3938
rect 1654 3932 1657 3948
rect 1534 3862 1537 3888
rect 1558 3862 1561 3868
rect 1502 3852 1505 3858
rect 1442 3848 1446 3851
rect 1510 3842 1513 3858
rect 1582 3842 1585 3848
rect 1522 3818 1526 3821
rect 1560 3803 1562 3807
rect 1566 3803 1569 3807
rect 1573 3803 1576 3807
rect 1418 3748 1422 3751
rect 1390 3662 1393 3678
rect 1414 3672 1417 3738
rect 1446 3692 1449 3778
rect 1462 3762 1465 3788
rect 1590 3762 1593 3908
rect 1598 3862 1601 3908
rect 1642 3878 1646 3881
rect 1614 3872 1617 3878
rect 1622 3862 1625 3868
rect 1654 3862 1657 3878
rect 1642 3858 1646 3861
rect 1606 3832 1609 3858
rect 1638 3842 1641 3848
rect 1662 3831 1665 3978
rect 1670 3962 1673 3968
rect 1678 3952 1681 4098
rect 1766 4072 1769 4268
rect 1806 4251 1809 4318
rect 1814 4262 1817 4338
rect 1846 4272 1849 4298
rect 1826 4268 1830 4271
rect 1806 4248 1814 4251
rect 1786 4068 1790 4071
rect 1758 4062 1761 4068
rect 1722 4058 1726 4061
rect 1746 4058 1750 4061
rect 1774 4042 1777 4058
rect 1798 4052 1801 4118
rect 1686 3972 1689 3978
rect 1710 3972 1713 4018
rect 1726 3952 1729 3958
rect 1678 3942 1681 3948
rect 1686 3922 1689 3948
rect 1726 3932 1729 3938
rect 1710 3882 1713 3918
rect 1734 3882 1737 3968
rect 1742 3881 1745 4018
rect 1754 3938 1758 3941
rect 1766 3932 1769 3938
rect 1742 3878 1750 3881
rect 1694 3852 1697 3878
rect 1774 3862 1777 3978
rect 1806 3961 1809 4218
rect 1822 4202 1825 4218
rect 1822 4151 1825 4168
rect 1838 4132 1841 4138
rect 1854 4122 1857 4128
rect 1822 4072 1825 4088
rect 1814 4032 1817 4068
rect 1834 4058 1838 4061
rect 1846 4052 1849 4098
rect 1854 3982 1857 4068
rect 1862 4032 1865 4418
rect 1870 4352 1873 4418
rect 1878 4341 1881 4428
rect 1942 4422 1945 4458
rect 1950 4432 1953 4468
rect 1910 4362 1913 4368
rect 1902 4352 1905 4358
rect 1874 4338 1881 4341
rect 1870 4161 1873 4338
rect 1886 4332 1889 4338
rect 1882 4258 1886 4261
rect 1882 4168 1886 4171
rect 1870 4158 1881 4161
rect 1870 4142 1873 4148
rect 1862 3962 1865 4008
rect 1870 3992 1873 4138
rect 1878 4122 1881 4158
rect 1910 4152 1913 4308
rect 1918 4292 1921 4318
rect 1918 4182 1921 4238
rect 1926 4232 1929 4338
rect 1942 4292 1945 4408
rect 1950 4392 1953 4428
rect 1958 4412 1961 4468
rect 1982 4462 1985 4468
rect 1990 4462 1993 4518
rect 2022 4512 2025 4528
rect 2010 4488 2014 4491
rect 2022 4472 2025 4508
rect 2072 4503 2074 4507
rect 2078 4503 2081 4507
rect 2085 4503 2088 4507
rect 2134 4482 2137 4548
rect 2142 4532 2145 4558
rect 2158 4552 2161 4588
rect 2190 4562 2193 4568
rect 2166 4552 2169 4558
rect 2154 4548 2158 4551
rect 2186 4538 2190 4541
rect 2206 4532 2209 4548
rect 2154 4528 2158 4531
rect 2214 4531 2217 4638
rect 2222 4562 2225 4568
rect 2230 4551 2233 4618
rect 2238 4572 2241 4648
rect 2246 4612 2249 4738
rect 2270 4682 2273 4778
rect 2278 4752 2281 4758
rect 2286 4682 2289 4768
rect 2294 4682 2297 4858
rect 2302 4812 2305 4868
rect 2362 4859 2366 4862
rect 2398 4862 2401 4888
rect 2462 4872 2465 4878
rect 2598 4872 2601 4878
rect 2894 4872 2897 4878
rect 3070 4872 3073 4878
rect 2426 4868 2430 4871
rect 2690 4868 2694 4871
rect 2730 4868 2734 4871
rect 2478 4863 2481 4868
rect 2442 4858 2446 4861
rect 2814 4862 2817 4868
rect 2506 4858 2510 4861
rect 2706 4858 2710 4861
rect 2786 4858 2790 4861
rect 2834 4858 2838 4861
rect 2322 4768 2326 4771
rect 2342 4752 2345 4858
rect 2362 4768 2366 4771
rect 2330 4738 2334 4741
rect 2342 4672 2345 4748
rect 2350 4692 2353 4758
rect 2374 4742 2377 4748
rect 2366 4672 2369 4708
rect 2266 4668 2270 4671
rect 2322 4668 2326 4671
rect 2374 4662 2377 4668
rect 2298 4658 2302 4661
rect 2330 4658 2334 4661
rect 2254 4572 2257 4658
rect 2382 4632 2385 4748
rect 2390 4692 2393 4738
rect 2422 4701 2425 4858
rect 2446 4842 2449 4848
rect 2502 4792 2505 4838
rect 2482 4768 2486 4771
rect 2502 4752 2505 4758
rect 2510 4752 2513 4858
rect 2550 4852 2553 4858
rect 2654 4822 2657 4858
rect 2686 4842 2689 4848
rect 2670 4832 2673 4838
rect 2538 4818 2542 4821
rect 2518 4772 2521 4818
rect 2566 4762 2569 4818
rect 2584 4803 2586 4807
rect 2590 4803 2593 4807
rect 2597 4803 2600 4807
rect 2654 4752 2657 4818
rect 2694 4772 2697 4858
rect 2702 4842 2705 4848
rect 2702 4752 2705 4768
rect 2718 4762 2721 4768
rect 2710 4758 2718 4761
rect 2450 4748 2454 4751
rect 2554 4748 2558 4751
rect 2430 4742 2433 4748
rect 2494 4722 2497 4738
rect 2418 4698 2425 4701
rect 2414 4662 2417 4698
rect 2422 4672 2425 4678
rect 2510 4672 2513 4748
rect 2542 4742 2545 4748
rect 2562 4738 2566 4741
rect 2526 4732 2529 4738
rect 2402 4658 2406 4661
rect 2482 4658 2486 4661
rect 2394 4638 2398 4641
rect 2426 4638 2430 4641
rect 2222 4548 2233 4551
rect 2270 4552 2273 4608
rect 2278 4562 2281 4618
rect 2222 4542 2225 4548
rect 2270 4542 2273 4548
rect 2238 4532 2241 4538
rect 2214 4528 2225 4531
rect 2174 4492 2177 4518
rect 2190 4512 2193 4518
rect 2222 4492 2225 4528
rect 2038 4472 2041 4478
rect 2242 4468 2246 4471
rect 1998 4462 2001 4468
rect 1966 4442 1969 4458
rect 2006 4372 2009 4468
rect 2030 4462 2033 4468
rect 2254 4462 2257 4498
rect 2022 4432 2025 4458
rect 2062 4392 2065 4458
rect 2150 4452 2153 4459
rect 2182 4442 2185 4458
rect 2246 4452 2249 4458
rect 2062 4352 2065 4378
rect 2078 4362 2081 4368
rect 2086 4352 2089 4418
rect 2094 4411 2097 4418
rect 2094 4408 2105 4411
rect 1958 4302 1961 4328
rect 1966 4312 1969 4348
rect 2054 4342 2057 4348
rect 2062 4342 2065 4348
rect 2094 4342 2097 4388
rect 1958 4272 1961 4298
rect 1982 4262 1985 4338
rect 2038 4322 2041 4328
rect 2014 4318 2022 4321
rect 1998 4292 2001 4308
rect 2014 4282 2017 4318
rect 1990 4262 1993 4268
rect 1970 4258 1974 4261
rect 1958 4222 1961 4258
rect 1918 4172 1921 4178
rect 1890 4138 1894 4141
rect 1886 4062 1889 4068
rect 1894 4062 1897 4068
rect 1902 3982 1905 4058
rect 1910 4031 1913 4148
rect 1934 4142 1937 4148
rect 1942 4142 1945 4168
rect 1958 4151 1961 4218
rect 1966 4162 1969 4168
rect 1958 4148 1969 4151
rect 1918 4082 1921 4088
rect 1934 4072 1937 4118
rect 1910 4028 1918 4031
rect 1898 3968 1902 3971
rect 1798 3958 1809 3961
rect 1842 3958 1846 3961
rect 1782 3952 1785 3958
rect 1790 3922 1793 3928
rect 1798 3881 1801 3958
rect 1790 3878 1801 3881
rect 1806 3922 1809 3948
rect 1814 3942 1817 3948
rect 1822 3942 1825 3958
rect 1790 3872 1793 3878
rect 1798 3862 1801 3868
rect 1754 3858 1758 3861
rect 1662 3828 1673 3831
rect 1494 3742 1497 3748
rect 1518 3742 1521 3748
rect 1478 3722 1481 3738
rect 1470 3691 1473 3718
rect 1470 3688 1481 3691
rect 1470 3672 1473 3678
rect 1458 3668 1462 3671
rect 1478 3662 1481 3688
rect 1510 3672 1513 3698
rect 1590 3682 1593 3758
rect 1646 3752 1649 3758
rect 1606 3702 1609 3718
rect 1598 3672 1601 3678
rect 1522 3668 1526 3671
rect 1466 3658 1470 3661
rect 1482 3648 1494 3651
rect 1310 3562 1313 3578
rect 1354 3568 1358 3571
rect 1314 3548 1318 3551
rect 1294 3502 1297 3518
rect 1270 3492 1273 3498
rect 1250 3488 1254 3491
rect 1286 3482 1289 3488
rect 1262 3462 1265 3468
rect 1250 3458 1254 3461
rect 1286 3412 1289 3478
rect 1302 3472 1305 3518
rect 1306 3458 1310 3461
rect 1318 3452 1321 3458
rect 1318 3402 1321 3418
rect 1254 3312 1257 3348
rect 1278 3332 1281 3358
rect 1294 3352 1297 3368
rect 1318 3362 1321 3368
rect 1198 3298 1209 3301
rect 1206 3282 1209 3298
rect 1174 3252 1177 3258
rect 1198 3242 1201 3278
rect 1254 3262 1257 3278
rect 1270 3262 1273 3288
rect 1294 3271 1297 3348
rect 1302 3332 1305 3338
rect 1310 3292 1313 3358
rect 1294 3268 1305 3271
rect 1314 3268 1318 3271
rect 1226 3258 1230 3261
rect 1290 3258 1294 3261
rect 1110 3142 1113 3148
rect 1134 3142 1137 3148
rect 1142 3142 1145 3148
rect 1158 3141 1161 3158
rect 1166 3152 1169 3158
rect 1182 3152 1185 3158
rect 1190 3152 1193 3218
rect 1198 3172 1201 3198
rect 1158 3138 1166 3141
rect 1194 3138 1198 3141
rect 1118 3092 1121 3118
rect 1086 3078 1097 3081
rect 1014 3058 1022 3061
rect 990 3052 993 3058
rect 998 3022 1001 3058
rect 966 2942 969 2948
rect 974 2942 977 2988
rect 862 2922 865 2928
rect 862 2862 865 2898
rect 870 2862 873 2868
rect 902 2862 905 2868
rect 910 2862 913 2878
rect 942 2872 945 2888
rect 934 2862 937 2868
rect 950 2862 953 2908
rect 958 2902 961 2918
rect 982 2872 985 2948
rect 998 2911 1001 3008
rect 1014 2982 1017 3018
rect 1038 3012 1041 3068
rect 1038 2992 1041 2998
rect 1014 2952 1017 2968
rect 1022 2952 1025 2958
rect 1070 2952 1073 3038
rect 1042 2948 1046 2951
rect 1006 2922 1009 2948
rect 1070 2932 1073 2948
rect 990 2908 1001 2911
rect 990 2872 993 2908
rect 998 2882 1001 2888
rect 778 2858 782 2861
rect 758 2852 761 2858
rect 870 2842 873 2858
rect 758 2812 761 2818
rect 790 2802 793 2818
rect 802 2758 806 2761
rect 818 2748 822 2751
rect 742 2722 745 2748
rect 814 2732 817 2738
rect 798 2681 801 2718
rect 790 2678 801 2681
rect 718 2592 721 2658
rect 726 2622 729 2628
rect 710 2502 713 2547
rect 726 2542 729 2598
rect 750 2592 753 2608
rect 758 2602 761 2638
rect 742 2542 745 2548
rect 758 2512 761 2558
rect 766 2542 769 2618
rect 774 2592 777 2598
rect 774 2542 777 2548
rect 702 2482 705 2498
rect 770 2468 774 2471
rect 646 2462 649 2468
rect 702 2463 705 2468
rect 666 2458 670 2461
rect 638 2352 641 2448
rect 654 2422 657 2458
rect 666 2448 670 2451
rect 758 2392 761 2468
rect 782 2462 785 2618
rect 790 2602 793 2678
rect 798 2652 801 2658
rect 806 2632 809 2668
rect 782 2452 785 2458
rect 782 2422 785 2428
rect 766 2362 769 2418
rect 646 2352 649 2358
rect 790 2352 793 2578
rect 798 2562 801 2568
rect 806 2551 809 2598
rect 822 2582 825 2738
rect 854 2732 857 2758
rect 870 2752 873 2778
rect 870 2742 873 2748
rect 878 2742 881 2748
rect 866 2728 870 2731
rect 838 2722 841 2728
rect 846 2722 849 2728
rect 902 2692 905 2858
rect 982 2852 985 2858
rect 930 2848 934 2851
rect 934 2792 937 2838
rect 958 2782 961 2818
rect 970 2788 974 2791
rect 990 2762 993 2868
rect 1014 2862 1017 2928
rect 1048 2903 1050 2907
rect 1054 2903 1057 2907
rect 1061 2903 1064 2907
rect 1030 2862 1033 2878
rect 1054 2862 1057 2878
rect 1070 2871 1073 2918
rect 1062 2868 1073 2871
rect 1062 2862 1065 2868
rect 1070 2851 1073 2858
rect 1062 2848 1073 2851
rect 954 2748 958 2751
rect 978 2738 982 2741
rect 950 2682 953 2718
rect 874 2678 878 2681
rect 838 2672 841 2678
rect 982 2672 985 2678
rect 842 2658 846 2661
rect 950 2652 953 2659
rect 866 2648 870 2651
rect 846 2642 849 2648
rect 902 2632 905 2638
rect 830 2562 833 2608
rect 802 2548 809 2551
rect 814 2552 817 2558
rect 846 2552 849 2558
rect 862 2552 865 2578
rect 854 2542 857 2548
rect 870 2542 873 2618
rect 902 2542 905 2578
rect 910 2552 913 2578
rect 826 2538 830 2541
rect 882 2538 886 2541
rect 866 2528 870 2531
rect 882 2528 886 2531
rect 798 2522 801 2528
rect 798 2452 801 2488
rect 806 2462 809 2468
rect 814 2462 817 2488
rect 830 2472 833 2518
rect 830 2452 833 2458
rect 838 2452 841 2458
rect 854 2392 857 2478
rect 870 2462 873 2478
rect 886 2472 889 2478
rect 894 2462 897 2518
rect 902 2472 905 2538
rect 918 2532 921 2548
rect 922 2528 926 2531
rect 934 2521 937 2598
rect 966 2552 969 2668
rect 986 2658 990 2661
rect 990 2642 993 2648
rect 998 2611 1001 2818
rect 1046 2792 1049 2818
rect 1062 2752 1065 2848
rect 1078 2842 1081 3038
rect 1086 2892 1089 3078
rect 1094 3052 1097 3068
rect 1094 3032 1097 3048
rect 1102 3042 1105 3058
rect 1118 2962 1121 3018
rect 1110 2942 1113 2948
rect 1118 2942 1121 2948
rect 1094 2902 1097 2918
rect 1098 2878 1102 2881
rect 1110 2872 1113 2938
rect 1098 2858 1102 2861
rect 1122 2858 1126 2861
rect 1134 2792 1137 3138
rect 1142 3082 1145 3138
rect 1166 3062 1169 3088
rect 1174 3062 1177 3098
rect 1182 3072 1185 3128
rect 1206 3092 1209 3238
rect 1218 3178 1222 3181
rect 1238 3162 1241 3238
rect 1238 3152 1241 3158
rect 1234 3138 1238 3141
rect 1246 3112 1249 3218
rect 1258 3158 1262 3161
rect 1270 3122 1273 3258
rect 1302 3252 1305 3268
rect 1282 3248 1286 3251
rect 1302 3212 1305 3248
rect 1282 3178 1286 3181
rect 1282 3148 1286 3151
rect 1238 3092 1241 3108
rect 1278 3082 1281 3148
rect 1286 3132 1289 3138
rect 1302 3082 1305 3168
rect 1318 3151 1321 3178
rect 1326 3112 1329 3518
rect 1334 3452 1337 3498
rect 1350 3492 1353 3518
rect 1358 3492 1361 3568
rect 1406 3562 1409 3648
rect 1438 3552 1441 3628
rect 1458 3568 1462 3571
rect 1478 3552 1481 3598
rect 1490 3568 1494 3571
rect 1374 3482 1377 3548
rect 1486 3542 1489 3548
rect 1390 3502 1393 3518
rect 1402 3488 1406 3491
rect 1362 3478 1366 3481
rect 1414 3481 1417 3518
rect 1422 3502 1425 3538
rect 1430 3522 1433 3538
rect 1458 3518 1462 3521
rect 1414 3478 1425 3481
rect 1342 3452 1345 3478
rect 1358 3462 1361 3468
rect 1366 3442 1369 3458
rect 1382 3452 1385 3478
rect 1410 3468 1414 3471
rect 1394 3448 1398 3451
rect 1382 3442 1385 3448
rect 1350 3352 1353 3428
rect 1358 3362 1361 3418
rect 1406 3372 1409 3468
rect 1414 3422 1417 3458
rect 1414 3362 1417 3378
rect 1422 3361 1425 3478
rect 1462 3462 1465 3508
rect 1442 3458 1446 3461
rect 1430 3442 1433 3448
rect 1430 3402 1433 3438
rect 1422 3358 1430 3361
rect 1454 3361 1457 3428
rect 1462 3382 1465 3458
rect 1454 3358 1465 3361
rect 1334 3272 1337 3278
rect 1310 3092 1313 3108
rect 1210 3068 1214 3071
rect 1222 3062 1225 3068
rect 1286 3062 1289 3068
rect 1202 3058 1214 3061
rect 1142 3002 1145 3058
rect 1182 3052 1185 3058
rect 1194 3018 1198 3021
rect 1158 2982 1161 3018
rect 1190 2952 1193 2968
rect 1146 2948 1150 2951
rect 1146 2938 1150 2941
rect 1158 2932 1161 2948
rect 1182 2932 1185 2938
rect 1150 2861 1153 2928
rect 1222 2922 1225 3058
rect 1230 3032 1233 3058
rect 1254 3032 1257 3058
rect 1270 3042 1273 3058
rect 1166 2862 1169 2868
rect 1150 2858 1158 2861
rect 1174 2851 1177 2918
rect 1222 2882 1225 2888
rect 1182 2862 1185 2868
rect 1190 2862 1193 2868
rect 1230 2862 1233 2868
rect 1170 2848 1177 2851
rect 1142 2842 1145 2848
rect 1078 2742 1081 2748
rect 1102 2742 1105 2748
rect 1050 2738 1054 2741
rect 1046 2722 1049 2738
rect 1048 2703 1050 2707
rect 1054 2703 1057 2707
rect 1061 2703 1064 2707
rect 1030 2662 1033 2668
rect 1046 2662 1049 2678
rect 1062 2662 1065 2668
rect 1014 2652 1017 2658
rect 998 2608 1006 2611
rect 998 2551 1001 2558
rect 1014 2552 1017 2648
rect 1038 2562 1041 2568
rect 1034 2548 1038 2551
rect 926 2518 937 2521
rect 918 2492 921 2498
rect 906 2458 910 2461
rect 890 2448 894 2451
rect 862 2392 865 2448
rect 842 2368 846 2371
rect 814 2362 817 2368
rect 850 2358 854 2361
rect 614 2282 617 2348
rect 622 2342 625 2348
rect 630 2302 633 2348
rect 630 2262 633 2288
rect 618 2258 622 2261
rect 610 2248 614 2251
rect 574 2242 577 2248
rect 582 2192 585 2248
rect 598 2202 601 2218
rect 622 2192 625 2228
rect 638 2192 641 2338
rect 662 2322 665 2338
rect 694 2292 697 2348
rect 766 2332 769 2348
rect 674 2268 678 2271
rect 650 2258 654 2261
rect 678 2232 681 2258
rect 690 2248 694 2251
rect 702 2242 705 2268
rect 710 2262 713 2298
rect 742 2262 745 2318
rect 766 2301 769 2328
rect 782 2312 785 2328
rect 758 2298 769 2301
rect 726 2252 729 2258
rect 714 2248 718 2251
rect 582 2172 585 2188
rect 646 2172 649 2218
rect 682 2188 686 2191
rect 702 2182 705 2238
rect 614 2162 617 2168
rect 562 2138 566 2141
rect 590 2132 593 2158
rect 702 2152 705 2158
rect 642 2148 646 2151
rect 690 2148 694 2151
rect 746 2148 750 2151
rect 606 2142 609 2148
rect 630 2142 633 2148
rect 650 2128 654 2131
rect 494 2032 497 2068
rect 502 2062 505 2108
rect 522 2078 526 2081
rect 506 2048 510 2051
rect 534 2051 537 2078
rect 530 2048 537 2051
rect 486 1952 489 1958
rect 498 1948 502 1951
rect 518 1942 521 2008
rect 536 2003 538 2007
rect 542 2003 545 2007
rect 549 2003 552 2007
rect 542 1952 545 1958
rect 478 1928 486 1931
rect 486 1892 489 1928
rect 462 1862 465 1868
rect 470 1812 473 1858
rect 502 1832 505 1868
rect 470 1792 473 1808
rect 536 1803 538 1807
rect 542 1803 545 1807
rect 549 1803 552 1807
rect 430 1768 441 1771
rect 482 1768 486 1771
rect 430 1752 433 1758
rect 330 1668 334 1671
rect 382 1662 385 1668
rect 286 1592 289 1658
rect 310 1618 318 1621
rect 310 1572 313 1618
rect 262 1492 265 1518
rect 270 1512 273 1548
rect 326 1542 329 1548
rect 334 1542 337 1658
rect 374 1652 377 1658
rect 366 1592 369 1608
rect 422 1582 425 1698
rect 438 1672 441 1768
rect 542 1762 545 1768
rect 506 1748 510 1751
rect 486 1742 489 1748
rect 518 1742 521 1748
rect 494 1702 497 1738
rect 542 1732 545 1758
rect 494 1692 497 1698
rect 518 1682 521 1718
rect 498 1678 502 1681
rect 446 1662 449 1678
rect 470 1662 473 1678
rect 510 1672 513 1678
rect 490 1668 494 1671
rect 558 1662 561 2118
rect 582 2082 585 2118
rect 570 2058 574 2061
rect 598 2052 601 2118
rect 622 2062 625 2078
rect 646 2062 649 2098
rect 578 2048 582 2051
rect 566 1992 569 2018
rect 602 1968 606 1971
rect 638 1962 641 1968
rect 618 1958 622 1961
rect 618 1948 622 1951
rect 566 1932 569 1938
rect 606 1912 609 1938
rect 594 1868 598 1871
rect 646 1862 649 2058
rect 654 1952 657 2018
rect 662 2012 665 2138
rect 670 2042 673 2148
rect 678 2042 681 2048
rect 686 2042 689 2068
rect 694 2062 697 2108
rect 718 2102 721 2138
rect 702 2072 705 2078
rect 758 2072 761 2298
rect 766 2152 769 2268
rect 774 2201 777 2278
rect 790 2272 793 2338
rect 798 2322 801 2348
rect 786 2258 790 2261
rect 774 2198 785 2201
rect 766 2072 769 2118
rect 774 2072 777 2088
rect 710 2068 718 2071
rect 754 2068 758 2071
rect 654 1932 657 1948
rect 662 1942 665 2008
rect 694 1952 697 2058
rect 710 2052 713 2068
rect 718 2052 721 2058
rect 734 2022 737 2058
rect 746 2048 750 2051
rect 758 2012 761 2068
rect 782 2062 785 2198
rect 798 2162 801 2168
rect 806 2142 809 2268
rect 814 2262 817 2318
rect 822 2292 825 2358
rect 878 2352 881 2358
rect 886 2352 889 2408
rect 838 2301 841 2348
rect 874 2338 878 2341
rect 846 2332 849 2338
rect 834 2298 841 2301
rect 830 2272 833 2298
rect 846 2242 849 2268
rect 854 2262 857 2298
rect 870 2252 873 2278
rect 902 2272 905 2458
rect 926 2352 929 2518
rect 934 2482 937 2508
rect 982 2482 985 2538
rect 1014 2492 1017 2538
rect 1030 2532 1033 2538
rect 1038 2532 1041 2548
rect 1046 2521 1049 2658
rect 1054 2552 1057 2558
rect 1062 2542 1065 2658
rect 1070 2622 1073 2698
rect 1078 2672 1081 2738
rect 1090 2668 1097 2671
rect 1070 2552 1073 2618
rect 1078 2572 1081 2668
rect 1086 2652 1089 2658
rect 1094 2652 1097 2668
rect 1102 2662 1105 2678
rect 1118 2672 1121 2678
rect 1134 2652 1137 2659
rect 1142 2602 1145 2838
rect 1166 2752 1169 2788
rect 1158 2712 1161 2718
rect 1166 2702 1169 2748
rect 1174 2742 1177 2748
rect 1190 2742 1193 2798
rect 1210 2748 1214 2751
rect 1218 2738 1222 2741
rect 1182 2732 1185 2738
rect 1198 2712 1201 2728
rect 1198 2671 1201 2708
rect 1198 2668 1209 2671
rect 1198 2642 1201 2658
rect 1206 2652 1209 2668
rect 1182 2602 1185 2638
rect 1158 2578 1166 2581
rect 1038 2518 1049 2521
rect 950 2462 953 2468
rect 1038 2462 1041 2518
rect 1048 2503 1050 2507
rect 1054 2503 1057 2507
rect 1061 2503 1064 2507
rect 1050 2488 1054 2491
rect 982 2452 985 2459
rect 1078 2442 1081 2538
rect 1094 2482 1097 2568
rect 1146 2558 1150 2561
rect 1110 2542 1113 2548
rect 1102 2462 1105 2538
rect 1134 2532 1137 2558
rect 1158 2552 1161 2578
rect 1190 2552 1193 2558
rect 1198 2552 1201 2608
rect 1206 2552 1209 2568
rect 1166 2542 1169 2548
rect 1182 2542 1185 2548
rect 1154 2538 1158 2541
rect 1214 2532 1217 2548
rect 1126 2502 1129 2528
rect 1158 2492 1161 2498
rect 946 2388 950 2391
rect 1010 2348 1014 2351
rect 910 2312 913 2348
rect 918 2342 921 2348
rect 894 2262 897 2268
rect 918 2262 921 2268
rect 898 2248 902 2251
rect 910 2232 913 2258
rect 926 2231 929 2348
rect 934 2342 937 2348
rect 958 2302 961 2348
rect 946 2258 950 2261
rect 1006 2262 1009 2338
rect 1048 2303 1050 2307
rect 1054 2303 1057 2307
rect 1061 2303 1064 2307
rect 1046 2282 1049 2288
rect 982 2252 985 2259
rect 918 2228 929 2231
rect 842 2218 846 2221
rect 814 2152 817 2178
rect 822 2142 825 2148
rect 806 2081 809 2138
rect 814 2092 817 2118
rect 806 2078 817 2081
rect 802 2058 806 2061
rect 766 2052 769 2058
rect 794 2048 798 2051
rect 702 1952 705 1968
rect 798 1962 801 1968
rect 762 1958 766 1961
rect 662 1882 665 1938
rect 678 1932 681 1938
rect 570 1858 574 1861
rect 642 1858 646 1861
rect 574 1742 577 1748
rect 430 1642 433 1658
rect 470 1652 473 1658
rect 450 1648 454 1651
rect 486 1642 489 1658
rect 536 1603 538 1607
rect 542 1603 545 1607
rect 549 1603 552 1607
rect 366 1552 369 1558
rect 278 1522 281 1538
rect 334 1532 337 1538
rect 342 1502 345 1528
rect 382 1492 385 1558
rect 422 1552 425 1578
rect 550 1562 553 1568
rect 410 1548 414 1551
rect 442 1548 446 1551
rect 390 1502 393 1538
rect 422 1522 425 1538
rect 422 1512 425 1518
rect 166 1342 169 1408
rect 174 1392 177 1448
rect 198 1402 201 1458
rect 214 1452 217 1478
rect 294 1472 297 1478
rect 230 1468 238 1471
rect 274 1468 278 1471
rect 222 1422 225 1428
rect 230 1402 233 1468
rect 274 1458 278 1461
rect 222 1352 225 1368
rect 166 1292 169 1328
rect 190 1322 193 1338
rect 238 1292 241 1428
rect 246 1421 249 1458
rect 254 1432 257 1448
rect 310 1422 313 1459
rect 366 1432 369 1448
rect 370 1428 374 1431
rect 246 1418 257 1421
rect 254 1342 257 1418
rect 274 1388 278 1391
rect 290 1368 294 1371
rect 290 1348 294 1351
rect 278 1322 281 1338
rect 194 1288 198 1291
rect 182 1272 185 1278
rect 254 1272 257 1318
rect 226 1268 230 1271
rect 150 1152 153 1258
rect 126 1062 129 1068
rect 134 1062 137 1068
rect 150 1062 153 1148
rect 158 1072 161 1268
rect 166 1232 169 1248
rect 214 1242 217 1268
rect 234 1248 238 1251
rect 166 1192 169 1208
rect 238 1192 241 1238
rect 190 1162 193 1168
rect 186 1148 190 1151
rect 118 1021 121 1058
rect 134 1022 137 1038
rect 118 1018 129 1021
rect 98 988 102 991
rect 110 942 113 948
rect 14 872 17 938
rect 62 932 65 938
rect 98 888 102 891
rect 106 868 110 871
rect 14 742 17 868
rect 42 858 46 861
rect 110 802 113 858
rect 118 852 121 858
rect 126 802 129 1018
rect 134 992 137 1018
rect 158 982 161 1068
rect 166 1052 169 1078
rect 178 1068 182 1071
rect 190 1061 193 1148
rect 198 1142 201 1178
rect 206 1162 209 1168
rect 214 1152 217 1158
rect 198 1071 201 1138
rect 214 1082 217 1088
rect 198 1068 206 1071
rect 190 1058 198 1061
rect 182 1052 185 1058
rect 198 1052 201 1058
rect 214 1042 217 1048
rect 198 1032 201 1038
rect 194 988 198 991
rect 134 952 137 958
rect 134 852 137 888
rect 158 872 161 978
rect 198 942 201 968
rect 206 962 209 968
rect 214 951 217 1008
rect 210 948 217 951
rect 174 872 177 938
rect 150 862 153 868
rect 14 692 17 738
rect 38 732 41 748
rect 14 672 17 688
rect 14 542 17 618
rect 38 552 41 558
rect 14 482 17 488
rect 30 462 33 468
rect 38 452 41 458
rect 46 342 49 538
rect 54 462 57 798
rect 134 752 137 828
rect 94 722 97 738
rect 70 672 73 708
rect 102 702 105 748
rect 110 742 113 748
rect 150 732 153 738
rect 118 722 121 728
rect 86 672 89 678
rect 114 658 118 661
rect 98 568 102 571
rect 114 558 118 561
rect 98 538 102 541
rect 62 472 65 518
rect 54 352 57 418
rect 46 292 49 338
rect 46 272 49 288
rect 62 282 65 468
rect 86 462 89 478
rect 94 472 97 528
rect 102 472 105 508
rect 102 462 105 468
rect 74 458 78 461
rect 110 452 113 548
rect 126 472 129 698
rect 134 562 137 568
rect 150 552 153 568
rect 158 552 161 868
rect 198 852 201 938
rect 206 881 209 948
rect 206 878 214 881
rect 166 732 169 748
rect 166 692 169 728
rect 174 722 177 848
rect 182 792 185 818
rect 198 752 201 778
rect 206 772 209 858
rect 222 821 225 1148
rect 246 1142 249 1148
rect 230 1072 233 1138
rect 270 1132 273 1268
rect 278 1262 281 1308
rect 246 1122 249 1128
rect 270 1082 273 1128
rect 234 1068 238 1071
rect 278 1071 281 1148
rect 290 1138 294 1141
rect 270 1068 281 1071
rect 230 972 233 988
rect 222 818 233 821
rect 222 752 225 808
rect 174 702 177 718
rect 174 662 177 698
rect 182 672 185 748
rect 190 742 193 748
rect 230 742 233 818
rect 238 792 241 1058
rect 262 992 265 998
rect 270 972 273 1068
rect 278 1042 281 1058
rect 246 922 249 948
rect 258 938 262 941
rect 246 862 249 918
rect 254 892 257 928
rect 238 762 241 768
rect 258 758 262 761
rect 270 752 273 968
rect 286 872 289 878
rect 302 872 305 1398
rect 310 1372 313 1388
rect 326 1352 329 1358
rect 334 1342 337 1398
rect 382 1392 385 1448
rect 350 1352 353 1358
rect 346 1338 350 1341
rect 334 1292 337 1298
rect 350 1292 353 1328
rect 358 1312 361 1338
rect 366 1292 369 1318
rect 374 1302 377 1358
rect 390 1352 393 1498
rect 422 1482 425 1508
rect 446 1492 449 1538
rect 454 1522 457 1548
rect 506 1547 510 1550
rect 470 1522 473 1528
rect 398 1472 401 1478
rect 406 1422 409 1478
rect 334 1252 337 1288
rect 358 1282 361 1288
rect 366 1272 369 1288
rect 390 1262 393 1348
rect 398 1342 401 1398
rect 422 1392 425 1478
rect 450 1468 454 1471
rect 430 1452 433 1458
rect 430 1362 433 1368
rect 410 1348 414 1351
rect 426 1348 430 1351
rect 410 1338 414 1341
rect 346 1258 350 1261
rect 378 1258 382 1261
rect 390 1242 393 1248
rect 398 1222 401 1268
rect 406 1232 409 1238
rect 374 1192 377 1218
rect 366 1132 369 1138
rect 342 1082 345 1118
rect 318 952 321 988
rect 326 942 329 1078
rect 382 1071 385 1178
rect 390 1152 393 1188
rect 378 1068 385 1071
rect 406 1072 409 1088
rect 414 1072 417 1338
rect 446 1321 449 1448
rect 454 1402 457 1468
rect 462 1462 465 1498
rect 486 1492 489 1538
rect 494 1472 497 1488
rect 518 1462 521 1498
rect 462 1452 465 1458
rect 462 1362 465 1418
rect 478 1392 481 1438
rect 526 1392 529 1418
rect 536 1403 538 1407
rect 542 1403 545 1407
rect 549 1403 552 1407
rect 522 1388 526 1391
rect 466 1347 470 1350
rect 438 1318 449 1321
rect 462 1322 465 1328
rect 438 1292 441 1318
rect 450 1278 454 1281
rect 450 1268 454 1271
rect 450 1248 454 1251
rect 430 1192 433 1238
rect 462 1192 465 1308
rect 470 1262 473 1268
rect 486 1262 489 1288
rect 510 1262 513 1298
rect 442 1188 446 1191
rect 470 1152 473 1158
rect 502 1142 505 1228
rect 526 1192 529 1328
rect 550 1282 553 1358
rect 534 1252 537 1258
rect 558 1212 561 1658
rect 566 1542 569 1718
rect 574 1692 577 1708
rect 578 1668 582 1671
rect 606 1662 609 1668
rect 614 1662 617 1738
rect 622 1672 625 1748
rect 638 1672 641 1738
rect 654 1671 657 1868
rect 666 1859 670 1862
rect 702 1862 705 1868
rect 710 1862 713 1958
rect 790 1952 793 1958
rect 778 1938 782 1941
rect 758 1912 761 1918
rect 734 1882 737 1908
rect 746 1888 750 1891
rect 754 1868 758 1871
rect 722 1858 726 1861
rect 710 1852 713 1858
rect 730 1848 734 1851
rect 750 1822 753 1858
rect 766 1852 769 1918
rect 782 1892 785 1908
rect 790 1892 793 1938
rect 798 1922 801 1938
rect 806 1922 809 2048
rect 814 1932 817 2078
rect 822 2072 825 2128
rect 830 2062 833 2198
rect 842 2158 846 2161
rect 854 2152 857 2158
rect 846 2148 854 2151
rect 838 2062 841 2078
rect 846 2022 849 2148
rect 870 2142 873 2188
rect 886 2162 889 2218
rect 918 2202 921 2228
rect 918 2182 921 2188
rect 926 2162 929 2218
rect 934 2192 937 2218
rect 910 2152 913 2158
rect 906 2138 910 2141
rect 862 2132 865 2138
rect 894 2132 897 2138
rect 886 2112 889 2118
rect 854 2082 857 2088
rect 886 2072 889 2098
rect 822 1952 825 1958
rect 790 1872 793 1888
rect 802 1868 806 1871
rect 774 1852 777 1858
rect 782 1842 785 1848
rect 798 1832 801 1858
rect 814 1852 817 1868
rect 830 1862 833 2018
rect 838 1942 841 2008
rect 862 1992 865 2058
rect 854 1912 857 1948
rect 870 1882 873 2068
rect 910 2032 913 2058
rect 878 1952 881 1958
rect 886 1952 889 1958
rect 894 1952 897 1968
rect 902 1952 905 2028
rect 926 1971 929 2158
rect 942 2152 945 2158
rect 958 2152 961 2158
rect 938 2138 942 2141
rect 966 2141 969 2158
rect 982 2152 985 2178
rect 962 2138 969 2141
rect 974 2142 977 2148
rect 1006 2142 1009 2258
rect 1022 2142 1025 2147
rect 990 2132 993 2138
rect 974 2072 977 2128
rect 974 2052 977 2068
rect 982 2062 985 2108
rect 1006 2102 1009 2138
rect 1048 2103 1050 2107
rect 1054 2103 1057 2107
rect 1061 2103 1064 2107
rect 970 2038 974 2041
rect 982 2022 985 2028
rect 926 1968 937 1971
rect 922 1958 926 1961
rect 838 1872 841 1878
rect 882 1858 886 1861
rect 710 1762 713 1768
rect 738 1758 742 1761
rect 686 1742 689 1748
rect 694 1732 697 1758
rect 702 1741 705 1758
rect 758 1752 761 1818
rect 814 1802 817 1838
rect 838 1792 841 1798
rect 722 1748 726 1751
rect 774 1751 777 1758
rect 870 1752 873 1778
rect 878 1752 881 1768
rect 742 1742 745 1748
rect 702 1738 710 1741
rect 718 1732 721 1738
rect 686 1722 689 1728
rect 674 1718 678 1721
rect 702 1692 705 1718
rect 650 1668 657 1671
rect 686 1662 689 1668
rect 674 1658 678 1661
rect 578 1648 582 1651
rect 590 1612 593 1658
rect 598 1592 601 1648
rect 606 1632 609 1648
rect 614 1642 617 1648
rect 646 1641 649 1658
rect 654 1652 657 1658
rect 662 1652 665 1658
rect 710 1652 713 1658
rect 670 1642 673 1648
rect 646 1638 657 1641
rect 622 1592 625 1628
rect 646 1592 649 1598
rect 614 1562 617 1568
rect 654 1562 657 1638
rect 662 1592 665 1638
rect 602 1548 609 1551
rect 606 1542 609 1548
rect 634 1538 638 1541
rect 566 1522 569 1528
rect 574 1482 577 1488
rect 566 1392 569 1398
rect 582 1362 585 1538
rect 606 1472 609 1538
rect 638 1511 641 1528
rect 654 1522 657 1558
rect 630 1508 641 1511
rect 622 1492 625 1498
rect 630 1492 633 1508
rect 598 1462 601 1468
rect 606 1442 609 1458
rect 630 1452 633 1488
rect 646 1452 649 1458
rect 598 1362 601 1368
rect 570 1348 574 1351
rect 602 1348 606 1351
rect 574 1332 577 1338
rect 570 1288 574 1291
rect 590 1272 593 1278
rect 598 1262 601 1318
rect 536 1203 538 1207
rect 542 1203 545 1207
rect 549 1203 552 1207
rect 590 1162 593 1168
rect 578 1158 582 1161
rect 598 1152 601 1258
rect 606 1152 609 1338
rect 614 1292 617 1438
rect 622 1352 625 1358
rect 614 1248 622 1251
rect 614 1172 617 1248
rect 614 1152 617 1168
rect 630 1162 633 1388
rect 646 1362 649 1448
rect 654 1412 657 1468
rect 662 1461 665 1558
rect 670 1542 673 1588
rect 686 1562 689 1608
rect 686 1542 689 1558
rect 670 1492 673 1518
rect 702 1492 705 1547
rect 674 1468 678 1471
rect 698 1468 702 1471
rect 662 1458 673 1461
rect 662 1372 665 1448
rect 670 1352 673 1458
rect 678 1412 681 1468
rect 690 1458 694 1461
rect 702 1432 705 1468
rect 662 1292 665 1298
rect 678 1292 681 1368
rect 694 1342 697 1347
rect 710 1292 713 1638
rect 726 1602 729 1668
rect 734 1662 737 1738
rect 766 1692 769 1708
rect 754 1688 758 1691
rect 734 1642 737 1658
rect 734 1482 737 1508
rect 750 1492 753 1648
rect 758 1622 761 1648
rect 774 1612 777 1728
rect 886 1712 889 1758
rect 894 1752 897 1948
rect 926 1942 929 1948
rect 934 1942 937 1968
rect 954 1958 958 1961
rect 966 1952 969 1958
rect 990 1952 993 2058
rect 1022 2052 1025 2058
rect 1006 2042 1009 2048
rect 998 1952 1001 1998
rect 1014 1992 1017 1998
rect 918 1792 921 1838
rect 918 1748 926 1751
rect 902 1742 905 1748
rect 826 1678 830 1681
rect 782 1672 785 1678
rect 894 1672 897 1728
rect 782 1622 785 1658
rect 790 1632 793 1668
rect 806 1662 809 1668
rect 814 1632 817 1658
rect 782 1602 785 1618
rect 770 1578 774 1581
rect 774 1562 777 1568
rect 774 1548 782 1551
rect 766 1512 769 1518
rect 774 1492 777 1548
rect 830 1542 833 1668
rect 918 1662 921 1748
rect 942 1742 945 1838
rect 958 1822 961 1918
rect 966 1862 969 1948
rect 982 1942 985 1948
rect 974 1851 977 1918
rect 1014 1872 1017 1958
rect 1022 1891 1025 2048
rect 1030 2022 1033 2068
rect 1038 2042 1041 2048
rect 1054 2042 1057 2068
rect 1070 2032 1073 2318
rect 1094 2262 1097 2438
rect 1142 2362 1145 2448
rect 1166 2432 1169 2458
rect 1174 2412 1177 2518
rect 1182 2492 1185 2498
rect 1182 2472 1185 2488
rect 1206 2422 1209 2458
rect 1222 2422 1225 2668
rect 1230 2612 1233 2828
rect 1238 2762 1241 2998
rect 1286 2952 1289 3038
rect 1246 2942 1249 2948
rect 1270 2942 1273 2948
rect 1294 2922 1297 3058
rect 1302 2932 1305 3078
rect 1314 3058 1318 3061
rect 1326 3052 1329 3088
rect 1334 3072 1337 3258
rect 1350 3152 1353 3348
rect 1358 3342 1361 3348
rect 1430 3342 1433 3348
rect 1454 3342 1457 3348
rect 1462 3342 1465 3358
rect 1470 3342 1473 3528
rect 1478 3492 1481 3528
rect 1358 3262 1361 3318
rect 1382 3272 1385 3328
rect 1442 3318 1446 3321
rect 1410 3258 1414 3261
rect 1366 3232 1369 3258
rect 1358 3072 1361 3078
rect 1346 3068 1350 3071
rect 1374 3062 1377 3188
rect 1382 3162 1385 3168
rect 1422 3132 1425 3318
rect 1478 3292 1481 3428
rect 1486 3272 1489 3538
rect 1502 3502 1505 3618
rect 1510 3512 1513 3658
rect 1526 3652 1529 3658
rect 1558 3652 1561 3668
rect 1578 3658 1582 3661
rect 1526 3632 1529 3648
rect 1590 3632 1593 3668
rect 1582 3622 1585 3628
rect 1502 3462 1505 3478
rect 1526 3472 1529 3618
rect 1560 3603 1562 3607
rect 1566 3603 1569 3607
rect 1573 3603 1576 3607
rect 1590 3552 1593 3628
rect 1598 3622 1601 3658
rect 1614 3652 1617 3658
rect 1606 3581 1609 3618
rect 1606 3578 1617 3581
rect 1550 3522 1553 3548
rect 1554 3458 1558 3461
rect 1502 3362 1505 3458
rect 1582 3452 1585 3488
rect 1526 3362 1529 3378
rect 1494 3352 1497 3358
rect 1534 3352 1537 3398
rect 1542 3392 1545 3418
rect 1560 3403 1562 3407
rect 1566 3403 1569 3407
rect 1573 3403 1576 3407
rect 1546 3378 1550 3381
rect 1574 3372 1577 3378
rect 1498 3338 1502 3341
rect 1510 3332 1513 3348
rect 1526 3342 1529 3348
rect 1590 3342 1593 3538
rect 1606 3532 1609 3568
rect 1614 3561 1617 3578
rect 1622 3572 1625 3748
rect 1634 3738 1638 3741
rect 1662 3662 1665 3818
rect 1670 3762 1673 3828
rect 1702 3792 1705 3838
rect 1710 3832 1713 3858
rect 1742 3852 1745 3858
rect 1710 3781 1713 3828
rect 1702 3778 1713 3781
rect 1694 3762 1697 3768
rect 1670 3742 1673 3748
rect 1686 3742 1689 3748
rect 1614 3558 1622 3561
rect 1634 3548 1638 3551
rect 1622 3541 1625 3548
rect 1622 3538 1646 3541
rect 1606 3472 1609 3478
rect 1622 3462 1625 3518
rect 1602 3458 1606 3461
rect 1614 3452 1617 3458
rect 1654 3432 1657 3608
rect 1662 3592 1665 3598
rect 1670 3451 1673 3718
rect 1702 3682 1705 3778
rect 1730 3768 1734 3771
rect 1714 3738 1718 3741
rect 1718 3722 1721 3728
rect 1730 3718 1737 3721
rect 1726 3692 1729 3708
rect 1734 3671 1737 3718
rect 1742 3702 1745 3848
rect 1798 3842 1801 3858
rect 1806 3832 1809 3918
rect 1822 3882 1825 3888
rect 1814 3852 1817 3868
rect 1830 3851 1833 3918
rect 1826 3848 1833 3851
rect 1750 3782 1753 3788
rect 1766 3782 1769 3818
rect 1766 3762 1769 3768
rect 1750 3752 1753 3758
rect 1766 3722 1769 3738
rect 1726 3668 1737 3671
rect 1678 3652 1681 3658
rect 1686 3552 1689 3668
rect 1698 3558 1702 3561
rect 1678 3521 1681 3548
rect 1686 3532 1689 3538
rect 1710 3522 1713 3528
rect 1678 3518 1689 3521
rect 1666 3448 1673 3451
rect 1678 3462 1681 3478
rect 1678 3442 1681 3458
rect 1686 3432 1689 3518
rect 1702 3491 1705 3518
rect 1702 3488 1713 3491
rect 1694 3481 1697 3488
rect 1694 3478 1702 3481
rect 1710 3452 1713 3488
rect 1598 3402 1601 3418
rect 1638 3412 1641 3418
rect 1606 3342 1609 3347
rect 1474 3268 1478 3271
rect 1490 3258 1494 3261
rect 1446 3142 1449 3238
rect 1466 3228 1470 3231
rect 1478 3192 1481 3258
rect 1518 3252 1521 3258
rect 1502 3232 1505 3238
rect 1446 3132 1449 3138
rect 1346 3058 1350 3061
rect 1358 2972 1361 3058
rect 1382 3052 1385 3128
rect 1394 3118 1398 3121
rect 1454 3121 1457 3147
rect 1446 3118 1457 3121
rect 1406 3082 1409 3118
rect 1446 3092 1449 3118
rect 1418 3088 1422 3091
rect 1470 3082 1473 3158
rect 1486 3132 1489 3198
rect 1534 3182 1537 3338
rect 1542 3272 1545 3318
rect 1498 3158 1502 3161
rect 1502 3142 1505 3148
rect 1526 3142 1529 3148
rect 1514 3138 1518 3141
rect 1394 3078 1398 3081
rect 1434 3078 1438 3081
rect 1482 3078 1486 3081
rect 1390 3062 1393 3068
rect 1406 3062 1409 3078
rect 1510 3072 1513 3118
rect 1526 3082 1529 3128
rect 1534 3122 1537 3148
rect 1450 3068 1454 3071
rect 1366 2992 1369 3018
rect 1438 2982 1441 3068
rect 1534 3062 1537 3088
rect 1542 3082 1545 3268
rect 1550 3162 1553 3218
rect 1560 3203 1562 3207
rect 1566 3203 1569 3207
rect 1573 3203 1576 3207
rect 1590 3162 1593 3168
rect 1578 3158 1582 3161
rect 1586 3138 1590 3141
rect 1458 3058 1462 3061
rect 1462 3002 1465 3058
rect 1346 2958 1350 2961
rect 1362 2958 1366 2961
rect 1374 2952 1377 2958
rect 1330 2948 1334 2951
rect 1342 2942 1345 2948
rect 1314 2938 1318 2941
rect 1350 2922 1353 2938
rect 1302 2892 1305 2918
rect 1314 2868 1318 2871
rect 1270 2842 1273 2848
rect 1282 2838 1286 2841
rect 1294 2772 1297 2868
rect 1342 2862 1345 2888
rect 1350 2872 1353 2918
rect 1358 2892 1361 2948
rect 1406 2942 1409 2947
rect 1418 2938 1422 2941
rect 1346 2858 1353 2861
rect 1302 2832 1305 2858
rect 1330 2838 1334 2841
rect 1266 2758 1270 2761
rect 1238 2752 1241 2758
rect 1342 2752 1345 2848
rect 1350 2842 1353 2858
rect 1382 2852 1385 2868
rect 1390 2852 1393 2858
rect 1390 2762 1393 2798
rect 1350 2752 1353 2758
rect 1258 2748 1262 2751
rect 1262 2732 1265 2748
rect 1342 2742 1345 2748
rect 1278 2712 1281 2718
rect 1254 2672 1257 2708
rect 1238 2662 1241 2668
rect 1250 2658 1254 2661
rect 1230 2532 1233 2548
rect 1246 2462 1249 2468
rect 1230 2452 1233 2458
rect 1238 2452 1241 2458
rect 1186 2388 1190 2391
rect 1214 2372 1217 2418
rect 1102 2352 1105 2358
rect 1198 2352 1201 2368
rect 1210 2358 1214 2361
rect 1130 2348 1134 2351
rect 1210 2348 1214 2351
rect 1102 2342 1105 2348
rect 1110 2342 1113 2348
rect 1122 2338 1126 2341
rect 1114 2278 1121 2281
rect 1102 2272 1105 2278
rect 1118 2272 1121 2278
rect 1110 2262 1113 2268
rect 1078 2232 1081 2238
rect 1086 2162 1089 2168
rect 1094 2112 1097 2258
rect 1118 2242 1121 2258
rect 1118 2182 1121 2238
rect 1118 2132 1121 2158
rect 1126 2152 1129 2218
rect 1134 2182 1137 2338
rect 1150 2332 1153 2338
rect 1158 2332 1161 2338
rect 1150 2272 1153 2328
rect 1174 2312 1177 2348
rect 1202 2278 1206 2281
rect 1178 2268 1182 2271
rect 1214 2271 1217 2318
rect 1230 2302 1233 2338
rect 1238 2272 1241 2338
rect 1246 2272 1249 2458
rect 1206 2268 1217 2271
rect 1162 2258 1169 2261
rect 1194 2258 1198 2261
rect 1146 2248 1150 2251
rect 1154 2248 1158 2251
rect 1166 2232 1169 2258
rect 1206 2252 1209 2268
rect 1230 2262 1233 2268
rect 1214 2252 1217 2258
rect 1174 2192 1177 2238
rect 1238 2232 1241 2258
rect 1218 2218 1222 2221
rect 1150 2162 1153 2178
rect 1134 2152 1137 2158
rect 1182 2151 1185 2158
rect 1126 2132 1129 2138
rect 1094 2062 1097 2078
rect 1102 2072 1105 2118
rect 1122 2058 1126 2061
rect 1110 2042 1113 2058
rect 1098 2038 1102 2041
rect 1038 1962 1041 2028
rect 1030 1902 1033 1948
rect 1054 1942 1057 2008
rect 1110 1952 1113 2008
rect 1118 1952 1121 1998
rect 1134 1992 1137 2138
rect 1142 2062 1145 2138
rect 1166 2092 1169 2138
rect 1150 2072 1153 2078
rect 1166 2062 1169 2078
rect 1190 2072 1193 2078
rect 1206 2062 1209 2218
rect 1238 2092 1241 2228
rect 1246 2182 1249 2188
rect 1254 2162 1257 2378
rect 1262 2342 1265 2508
rect 1270 2352 1273 2648
rect 1286 2602 1289 2668
rect 1294 2652 1297 2658
rect 1346 2568 1350 2571
rect 1278 2552 1281 2558
rect 1302 2542 1305 2548
rect 1342 2492 1345 2548
rect 1278 2462 1281 2468
rect 1294 2462 1297 2468
rect 1302 2462 1305 2488
rect 1282 2448 1286 2451
rect 1302 2432 1305 2458
rect 1342 2452 1345 2488
rect 1286 2412 1289 2418
rect 1318 2412 1321 2418
rect 1290 2388 1294 2391
rect 1310 2391 1313 2408
rect 1310 2388 1321 2391
rect 1278 2381 1281 2388
rect 1278 2378 1289 2381
rect 1286 2372 1289 2378
rect 1278 2352 1281 2368
rect 1310 2352 1313 2378
rect 1318 2362 1321 2388
rect 1350 2352 1353 2508
rect 1358 2502 1361 2708
rect 1370 2668 1374 2671
rect 1390 2661 1393 2758
rect 1414 2742 1417 2918
rect 1386 2658 1393 2661
rect 1390 2652 1393 2658
rect 1398 2652 1401 2718
rect 1406 2712 1409 2738
rect 1430 2702 1433 2928
rect 1446 2882 1449 2888
rect 1450 2868 1454 2871
rect 1462 2862 1465 2908
rect 1470 2892 1473 3038
rect 1486 2992 1489 3048
rect 1498 3018 1502 3021
rect 1550 2982 1553 3118
rect 1598 3062 1601 3288
rect 1606 3272 1609 3328
rect 1610 3259 1614 3262
rect 1606 3152 1609 3238
rect 1614 3202 1617 3248
rect 1614 3152 1617 3198
rect 1630 3161 1633 3398
rect 1694 3392 1697 3448
rect 1666 3378 1670 3381
rect 1638 3352 1641 3368
rect 1678 3352 1681 3358
rect 1670 3272 1673 3278
rect 1650 3258 1654 3261
rect 1662 3252 1665 3258
rect 1646 3242 1649 3248
rect 1662 3192 1665 3248
rect 1670 3232 1673 3268
rect 1678 3192 1681 3348
rect 1686 3292 1689 3328
rect 1686 3202 1689 3218
rect 1694 3162 1697 3288
rect 1702 3262 1705 3428
rect 1710 3362 1713 3418
rect 1710 3292 1713 3318
rect 1718 3281 1721 3528
rect 1726 3471 1729 3668
rect 1758 3662 1761 3688
rect 1738 3658 1742 3661
rect 1750 3601 1753 3658
rect 1746 3598 1753 3601
rect 1726 3468 1734 3471
rect 1730 3458 1734 3461
rect 1726 3422 1729 3428
rect 1766 3421 1769 3718
rect 1782 3682 1785 3738
rect 1790 3662 1793 3718
rect 1798 3692 1801 3818
rect 1810 3748 1814 3751
rect 1822 3742 1825 3778
rect 1830 3752 1833 3818
rect 1838 3742 1841 3938
rect 1846 3872 1849 3878
rect 1854 3872 1857 3918
rect 1846 3812 1849 3858
rect 1854 3802 1857 3858
rect 1854 3752 1857 3788
rect 1862 3761 1865 3948
rect 1886 3932 1889 3948
rect 1874 3928 1878 3931
rect 1886 3882 1889 3928
rect 1874 3878 1878 3881
rect 1870 3862 1873 3868
rect 1886 3862 1889 3868
rect 1910 3862 1913 3998
rect 1934 3992 1937 4068
rect 1942 4032 1945 4058
rect 1950 4032 1953 4148
rect 1958 4052 1961 4058
rect 1966 4052 1969 4148
rect 1974 4092 1977 4248
rect 1982 4112 1985 4258
rect 2002 4168 2006 4171
rect 1994 4158 1998 4161
rect 1994 4148 1998 4151
rect 1990 4138 1998 4141
rect 1990 4112 1993 4138
rect 2022 4132 2025 4168
rect 2038 4122 2041 4258
rect 2046 4222 2049 4338
rect 2072 4303 2074 4307
rect 2078 4303 2081 4307
rect 2085 4303 2088 4307
rect 2062 4272 2065 4278
rect 2086 4242 2089 4258
rect 2062 4152 2065 4158
rect 2102 4142 2105 4408
rect 2114 4368 2118 4371
rect 2134 4362 2137 4368
rect 2114 4348 2118 4351
rect 2142 4342 2145 4378
rect 2134 4282 2137 4338
rect 2142 4332 2145 4338
rect 2150 4282 2153 4348
rect 2158 4342 2161 4348
rect 2166 4292 2169 4418
rect 2214 4372 2217 4418
rect 2190 4362 2193 4368
rect 2174 4332 2177 4338
rect 2150 4262 2153 4268
rect 2166 4252 2169 4278
rect 2174 4252 2177 4318
rect 2190 4302 2193 4318
rect 2198 4272 2201 4318
rect 2214 4282 2217 4288
rect 2222 4282 2225 4448
rect 2262 4431 2265 4438
rect 2270 4431 2273 4538
rect 2278 4512 2281 4548
rect 2294 4472 2297 4618
rect 2390 4552 2393 4558
rect 2354 4538 2358 4541
rect 2342 4532 2345 4538
rect 2358 4522 2361 4528
rect 2278 4462 2281 4468
rect 2298 4458 2302 4461
rect 2326 4442 2329 4448
rect 2334 4442 2337 4518
rect 2262 4428 2273 4431
rect 2302 4432 2305 4438
rect 2262 4342 2265 4428
rect 2270 4302 2273 4418
rect 2278 4322 2281 4347
rect 2222 4272 2225 4278
rect 2198 4262 2201 4268
rect 2238 4262 2241 4268
rect 2186 4258 2190 4261
rect 2246 4252 2249 4298
rect 2302 4292 2305 4318
rect 2334 4292 2337 4347
rect 2342 4322 2345 4468
rect 2350 4452 2353 4498
rect 2374 4472 2377 4538
rect 2398 4481 2401 4638
rect 2526 4622 2529 4668
rect 2534 4662 2537 4668
rect 2394 4478 2401 4481
rect 2414 4472 2417 4618
rect 2542 4602 2545 4738
rect 2582 4672 2585 4748
rect 2626 4747 2630 4750
rect 2654 4672 2657 4748
rect 2686 4722 2689 4728
rect 2694 4722 2697 4738
rect 2694 4692 2697 4718
rect 2562 4668 2566 4671
rect 2550 4652 2553 4658
rect 2574 4642 2577 4658
rect 2582 4632 2585 4668
rect 2630 4663 2633 4668
rect 2654 4662 2657 4668
rect 2694 4642 2697 4658
rect 2702 4631 2705 4748
rect 2710 4682 2713 4758
rect 2718 4662 2721 4738
rect 2726 4702 2729 4858
rect 2738 4828 2742 4831
rect 2726 4662 2729 4668
rect 2718 4632 2721 4658
rect 2702 4628 2713 4631
rect 2584 4603 2586 4607
rect 2590 4603 2593 4607
rect 2597 4603 2600 4607
rect 2526 4578 2534 4581
rect 2702 4581 2705 4618
rect 2698 4578 2705 4581
rect 2710 4582 2713 4628
rect 2726 4592 2729 4658
rect 2526 4562 2529 4578
rect 2466 4558 2470 4561
rect 2422 4551 2425 4558
rect 2486 4552 2489 4558
rect 2522 4548 2526 4551
rect 2454 4542 2457 4548
rect 2430 4492 2433 4508
rect 2418 4468 2422 4471
rect 2446 4462 2449 4508
rect 2454 4472 2457 4518
rect 2462 4502 2465 4548
rect 2534 4542 2537 4548
rect 2502 4532 2505 4538
rect 2362 4458 2366 4461
rect 2418 4458 2422 4461
rect 2418 4448 2430 4451
rect 2390 4442 2393 4448
rect 2270 4272 2273 4288
rect 2366 4282 2369 4418
rect 2382 4292 2385 4418
rect 2446 4382 2449 4458
rect 2394 4368 2398 4371
rect 2414 4352 2417 4368
rect 2442 4348 2446 4351
rect 2454 4351 2457 4468
rect 2486 4462 2489 4468
rect 2470 4458 2478 4461
rect 2462 4392 2465 4448
rect 2470 4362 2473 4458
rect 2478 4432 2481 4438
rect 2494 4402 2497 4458
rect 2510 4452 2513 4538
rect 2518 4492 2521 4518
rect 2566 4492 2569 4558
rect 2574 4542 2577 4548
rect 2590 4542 2593 4568
rect 2702 4562 2705 4568
rect 2710 4552 2713 4578
rect 2718 4562 2721 4568
rect 2610 4547 2614 4550
rect 2698 4548 2702 4551
rect 2674 4538 2678 4541
rect 2534 4482 2537 4488
rect 2530 4468 2534 4471
rect 2518 4462 2521 4468
rect 2542 4422 2545 4468
rect 2550 4462 2553 4468
rect 2574 4442 2577 4518
rect 2614 4482 2617 4538
rect 2686 4532 2689 4548
rect 2666 4518 2670 4521
rect 2674 4488 2678 4491
rect 2690 4468 2694 4471
rect 2614 4442 2617 4459
rect 2466 4358 2470 4361
rect 2482 4358 2486 4361
rect 2510 4352 2513 4378
rect 2530 4358 2534 4361
rect 2574 4361 2577 4438
rect 2694 4432 2697 4458
rect 2710 4422 2713 4538
rect 2718 4452 2721 4508
rect 2734 4482 2737 4828
rect 2754 4768 2758 4771
rect 2746 4758 2750 4761
rect 2814 4752 2817 4758
rect 2742 4702 2745 4748
rect 2838 4742 2841 4818
rect 2754 4738 2758 4741
rect 2854 4732 2857 4818
rect 2894 4802 2897 4868
rect 2982 4862 2985 4868
rect 2962 4858 2966 4861
rect 3010 4858 3014 4861
rect 3090 4858 3094 4861
rect 3050 4838 3054 4841
rect 3062 4762 3065 4818
rect 2862 4692 2865 4718
rect 2746 4658 2750 4661
rect 2742 4642 2745 4648
rect 2766 4642 2769 4678
rect 2878 4672 2881 4738
rect 2902 4712 2905 4748
rect 2974 4732 2977 4738
rect 2998 4722 3001 4748
rect 2782 4662 2785 4668
rect 2878 4662 2881 4668
rect 2798 4652 2801 4659
rect 2902 4642 2905 4658
rect 2858 4638 2862 4641
rect 2794 4548 2798 4551
rect 2846 4542 2849 4638
rect 2862 4562 2865 4638
rect 2958 4602 2961 4718
rect 3014 4672 3017 4688
rect 2986 4658 2990 4661
rect 3002 4648 3006 4651
rect 2862 4542 2865 4547
rect 2742 4492 2745 4518
rect 2798 4492 2801 4538
rect 2790 4472 2793 4488
rect 2806 4472 2809 4528
rect 2734 4461 2737 4468
rect 2730 4458 2737 4461
rect 2584 4403 2586 4407
rect 2590 4403 2593 4407
rect 2597 4403 2600 4407
rect 2574 4358 2582 4361
rect 2542 4352 2545 4358
rect 2662 4352 2665 4388
rect 2694 4372 2697 4418
rect 2710 4372 2713 4418
rect 2718 4362 2721 4368
rect 2454 4348 2465 4351
rect 2474 4348 2478 4351
rect 2406 4302 2409 4348
rect 2454 4332 2457 4338
rect 2462 4332 2465 4348
rect 2306 4268 2310 4271
rect 2278 4262 2281 4268
rect 2350 4262 2353 4278
rect 2374 4262 2377 4268
rect 2398 4262 2401 4298
rect 2422 4262 2425 4308
rect 2314 4258 2318 4261
rect 2386 4258 2390 4261
rect 2110 4162 2113 4248
rect 2122 4138 2126 4141
rect 2072 4103 2074 4107
rect 2078 4103 2081 4107
rect 2085 4103 2088 4107
rect 1990 4072 1993 4088
rect 1942 3952 1945 4028
rect 1958 4012 1961 4038
rect 1966 3992 1969 4048
rect 1982 4022 1985 4068
rect 1998 4062 2001 4088
rect 2102 4072 2105 4138
rect 2134 4132 2137 4138
rect 2142 4132 2145 4218
rect 2158 4152 2161 4218
rect 2170 4148 2174 4151
rect 2154 4118 2161 4121
rect 2142 4092 2145 4118
rect 2158 4102 2161 4118
rect 2018 4058 2025 4061
rect 2022 4052 2025 4058
rect 2078 4052 2081 4058
rect 2010 4048 2014 4051
rect 2022 4012 2025 4018
rect 1958 3951 1961 3958
rect 1974 3942 1977 3978
rect 2086 3972 2089 3978
rect 2022 3962 2025 3968
rect 1990 3952 1993 3958
rect 1998 3952 2001 3958
rect 2018 3948 2022 3951
rect 2042 3948 2046 3951
rect 2006 3942 2009 3948
rect 2018 3938 2022 3941
rect 2050 3938 2054 3941
rect 1930 3888 1934 3891
rect 1974 3872 1977 3938
rect 2074 3918 2078 3921
rect 2072 3903 2074 3907
rect 2078 3903 2081 3907
rect 2085 3903 2088 3907
rect 2022 3882 2025 3888
rect 2102 3872 2105 3898
rect 2110 3882 2113 3918
rect 2058 3868 2062 3871
rect 1990 3863 1993 3868
rect 2042 3858 2046 3861
rect 1878 3852 1881 3858
rect 2086 3852 2089 3858
rect 2110 3832 2113 3878
rect 1894 3762 1897 3768
rect 1862 3758 1873 3761
rect 1862 3742 1865 3748
rect 1870 3742 1873 3758
rect 1878 3752 1881 3758
rect 1870 3722 1873 3738
rect 1782 3652 1785 3658
rect 1774 3602 1777 3618
rect 1774 3551 1777 3558
rect 1790 3542 1793 3548
rect 1806 3542 1809 3698
rect 1846 3692 1849 3718
rect 1818 3678 1822 3681
rect 1846 3662 1849 3668
rect 1854 3662 1857 3678
rect 1886 3662 1889 3688
rect 1902 3682 1905 3818
rect 1910 3752 1913 3758
rect 1902 3662 1905 3668
rect 1826 3658 1830 3661
rect 1838 3652 1841 3658
rect 1814 3562 1817 3568
rect 1790 3462 1793 3538
rect 1814 3522 1817 3548
rect 1758 3418 1769 3421
rect 1750 3362 1753 3378
rect 1758 3342 1761 3418
rect 1774 3402 1777 3458
rect 1822 3391 1825 3618
rect 1838 3571 1841 3598
rect 1846 3592 1849 3658
rect 1870 3572 1873 3618
rect 1894 3602 1897 3658
rect 1918 3622 1921 3748
rect 1926 3742 1929 3818
rect 2018 3768 2022 3771
rect 2030 3761 2033 3818
rect 2070 3762 2073 3828
rect 2030 3758 2038 3761
rect 2050 3758 2054 3761
rect 1958 3751 1961 3758
rect 2118 3752 2121 4068
rect 2134 4042 2137 4058
rect 2150 4032 2153 4078
rect 2158 4072 2161 4098
rect 2182 4092 2185 4238
rect 2190 4092 2193 4218
rect 2206 4202 2209 4218
rect 2230 4152 2233 4158
rect 2162 4058 2166 4061
rect 2126 3872 2129 3928
rect 2134 3911 2137 3947
rect 2134 3908 2145 3911
rect 2142 3892 2145 3908
rect 2146 3868 2150 3871
rect 2126 3862 2129 3868
rect 2158 3852 2161 3858
rect 2166 3802 2169 3868
rect 2174 3862 2177 4088
rect 2214 4072 2217 4098
rect 2190 4052 2193 4058
rect 2190 3802 2193 4048
rect 2206 4011 2209 4068
rect 2222 4062 2225 4088
rect 2226 4018 2230 4021
rect 2202 4008 2209 4011
rect 2222 3952 2225 3978
rect 2198 3942 2201 3948
rect 2222 3872 2225 3948
rect 2238 3882 2241 4248
rect 2262 4172 2265 4218
rect 2270 4192 2273 4258
rect 2286 4252 2289 4258
rect 2342 4252 2345 4258
rect 2302 4242 2305 4248
rect 2334 4241 2337 4248
rect 2334 4238 2345 4241
rect 2342 4192 2345 4238
rect 2358 4212 2361 4218
rect 2414 4212 2417 4218
rect 2310 4172 2313 4178
rect 2358 4172 2361 4198
rect 2282 4158 2286 4161
rect 2270 4142 2273 4148
rect 2246 4072 2249 4078
rect 2254 3982 2257 4138
rect 2262 4052 2265 4118
rect 2270 4072 2273 4108
rect 2270 4032 2273 4068
rect 2278 4062 2281 4148
rect 2294 4132 2297 4158
rect 2306 4148 2310 4151
rect 2318 4141 2321 4158
rect 2306 4138 2321 4141
rect 2326 4142 2329 4158
rect 2366 4152 2369 4158
rect 2398 4152 2401 4178
rect 2430 4161 2433 4318
rect 2438 4282 2441 4288
rect 2458 4218 2465 4221
rect 2430 4158 2438 4161
rect 2418 4148 2422 4151
rect 2434 4148 2438 4151
rect 2334 4142 2337 4148
rect 2342 4112 2345 4148
rect 2386 4138 2390 4141
rect 2366 4132 2369 4138
rect 2446 4132 2449 4218
rect 2454 4152 2457 4168
rect 2438 4122 2441 4128
rect 2294 4062 2297 4098
rect 2302 4092 2305 4098
rect 2302 4052 2305 4058
rect 2302 3992 2305 4048
rect 2274 3958 2278 3961
rect 2302 3952 2305 3958
rect 2282 3938 2286 3941
rect 2254 3922 2257 3928
rect 2262 3902 2265 3938
rect 2198 3862 2201 3868
rect 2246 3862 2249 3868
rect 2206 3762 2209 3858
rect 2254 3792 2257 3808
rect 2246 3762 2249 3768
rect 2170 3758 2174 3761
rect 2262 3752 2265 3898
rect 2270 3772 2273 3778
rect 1986 3748 1990 3751
rect 2130 3748 2134 3751
rect 2234 3748 2238 3751
rect 2118 3742 2121 3748
rect 2030 3732 2033 3738
rect 2054 3732 2057 3738
rect 1926 3662 1929 3668
rect 1934 3662 1937 3668
rect 1942 3612 1945 3658
rect 1950 3652 1953 3658
rect 1958 3592 1961 3728
rect 2030 3722 2033 3728
rect 2206 3722 2209 3748
rect 2214 3742 2217 3748
rect 2230 3722 2233 3738
rect 2262 3732 2265 3738
rect 2274 3718 2278 3721
rect 2026 3678 2030 3681
rect 1982 3662 1985 3668
rect 2006 3662 2009 3668
rect 1974 3652 1977 3658
rect 1994 3648 1998 3651
rect 1966 3592 1969 3618
rect 1838 3568 1849 3571
rect 1838 3532 1841 3558
rect 1846 3462 1849 3568
rect 1902 3552 1905 3558
rect 1926 3552 1929 3588
rect 1962 3568 1966 3571
rect 1974 3552 1977 3628
rect 1998 3562 2001 3568
rect 1982 3552 1985 3558
rect 1854 3512 1857 3548
rect 1862 3532 1865 3538
rect 1838 3452 1841 3458
rect 1878 3452 1881 3458
rect 1886 3452 1889 3488
rect 1926 3462 1929 3548
rect 1958 3532 1961 3548
rect 1966 3532 1969 3538
rect 1974 3522 1977 3548
rect 1998 3522 2001 3558
rect 1950 3463 1953 3488
rect 1986 3468 1990 3471
rect 1998 3462 2001 3468
rect 1986 3458 1990 3461
rect 1886 3442 1889 3448
rect 1834 3418 1838 3421
rect 1814 3388 1825 3391
rect 1782 3372 1785 3378
rect 1738 3338 1742 3341
rect 1754 3338 1758 3341
rect 1726 3312 1729 3338
rect 1766 3332 1769 3348
rect 1714 3278 1721 3281
rect 1730 3258 1734 3261
rect 1702 3202 1705 3258
rect 1750 3252 1753 3318
rect 1734 3162 1737 3218
rect 1630 3158 1641 3161
rect 1674 3158 1678 3161
rect 1638 3152 1641 3158
rect 1626 3148 1630 3151
rect 1666 3148 1670 3151
rect 1698 3148 1702 3151
rect 1722 3148 1726 3151
rect 1690 3138 1694 3141
rect 1622 3082 1625 3138
rect 1654 3092 1657 3118
rect 1630 3082 1633 3088
rect 1638 3082 1641 3088
rect 1658 3078 1662 3081
rect 1590 3042 1593 3048
rect 1560 3003 1562 3007
rect 1566 3003 1569 3007
rect 1573 3003 1576 3007
rect 1598 3002 1601 3058
rect 1622 3032 1625 3068
rect 1646 3052 1649 3078
rect 1666 3068 1670 3071
rect 1674 3058 1678 3061
rect 1662 3032 1665 3058
rect 1686 3051 1689 3118
rect 1726 3112 1729 3138
rect 1694 3062 1697 3068
rect 1686 3048 1694 3051
rect 1586 2968 1590 2971
rect 1478 2952 1481 2968
rect 1538 2948 1542 2951
rect 1478 2932 1481 2948
rect 1606 2942 1609 3018
rect 1702 3012 1705 3068
rect 1710 3062 1713 3078
rect 1734 3062 1737 3148
rect 1734 3052 1737 3058
rect 1722 3048 1726 3051
rect 1710 3022 1713 3028
rect 1658 2968 1662 2971
rect 1682 2958 1686 2961
rect 1690 2958 1694 2961
rect 1618 2948 1622 2951
rect 1706 2948 1710 2951
rect 1742 2951 1745 3248
rect 1750 3122 1753 3128
rect 1750 3082 1753 3088
rect 1738 2948 1745 2951
rect 1638 2942 1641 2948
rect 1486 2852 1489 2878
rect 1518 2872 1521 2928
rect 1678 2922 1681 2948
rect 1694 2942 1697 2948
rect 1726 2942 1729 2948
rect 1714 2938 1718 2941
rect 1630 2912 1633 2918
rect 1534 2872 1537 2878
rect 1542 2872 1545 2888
rect 1506 2868 1510 2871
rect 1550 2862 1553 2888
rect 1578 2868 1582 2871
rect 1598 2862 1601 2908
rect 1622 2862 1625 2878
rect 1638 2862 1641 2868
rect 1646 2862 1649 2868
rect 1670 2862 1673 2888
rect 1678 2862 1681 2918
rect 1686 2872 1689 2938
rect 1466 2848 1470 2851
rect 1490 2848 1494 2851
rect 1502 2842 1505 2858
rect 1534 2852 1537 2858
rect 1514 2848 1518 2851
rect 1502 2792 1505 2798
rect 1466 2758 1470 2761
rect 1490 2758 1494 2761
rect 1438 2712 1441 2748
rect 1470 2742 1473 2758
rect 1486 2742 1489 2748
rect 1450 2738 1454 2741
rect 1406 2672 1409 2678
rect 1418 2668 1422 2671
rect 1378 2648 1382 2651
rect 1390 2562 1393 2608
rect 1370 2558 1374 2561
rect 1366 2532 1369 2548
rect 1382 2492 1385 2558
rect 1390 2532 1393 2558
rect 1406 2542 1409 2658
rect 1414 2542 1417 2548
rect 1406 2492 1409 2538
rect 1358 2462 1361 2488
rect 1422 2482 1425 2598
rect 1430 2592 1433 2648
rect 1438 2622 1441 2708
rect 1494 2682 1497 2698
rect 1446 2662 1449 2668
rect 1470 2662 1473 2678
rect 1506 2668 1513 2671
rect 1510 2662 1513 2668
rect 1478 2652 1481 2658
rect 1470 2632 1473 2638
rect 1446 2602 1449 2618
rect 1430 2542 1433 2548
rect 1462 2542 1465 2558
rect 1450 2538 1454 2541
rect 1470 2532 1473 2628
rect 1518 2592 1521 2828
rect 1550 2812 1553 2858
rect 1562 2848 1566 2851
rect 1560 2803 1562 2807
rect 1566 2803 1569 2807
rect 1573 2803 1576 2807
rect 1570 2748 1574 2751
rect 1526 2652 1529 2678
rect 1534 2662 1537 2718
rect 1550 2672 1553 2678
rect 1490 2558 1494 2561
rect 1510 2552 1513 2558
rect 1482 2548 1486 2551
rect 1494 2542 1497 2548
rect 1502 2542 1505 2548
rect 1430 2462 1433 2498
rect 1478 2492 1481 2538
rect 1482 2488 1486 2491
rect 1470 2452 1473 2488
rect 1494 2462 1497 2528
rect 1510 2492 1513 2498
rect 1526 2482 1529 2488
rect 1502 2462 1505 2468
rect 1534 2451 1537 2548
rect 1542 2502 1545 2658
rect 1550 2482 1553 2648
rect 1566 2622 1569 2668
rect 1582 2622 1585 2858
rect 1590 2851 1593 2858
rect 1590 2848 1598 2851
rect 1678 2842 1681 2858
rect 1686 2852 1689 2868
rect 1734 2862 1737 2948
rect 1742 2892 1745 2918
rect 1746 2868 1750 2871
rect 1734 2852 1737 2858
rect 1686 2832 1689 2848
rect 1710 2842 1713 2848
rect 1614 2802 1617 2818
rect 1662 2762 1665 2818
rect 1718 2792 1721 2828
rect 1678 2758 1686 2761
rect 1590 2752 1593 2758
rect 1666 2748 1670 2751
rect 1614 2682 1617 2738
rect 1630 2732 1633 2748
rect 1638 2742 1641 2748
rect 1678 2732 1681 2758
rect 1706 2738 1710 2741
rect 1646 2681 1649 2718
rect 1678 2692 1681 2728
rect 1638 2678 1649 2681
rect 1638 2662 1641 2678
rect 1694 2672 1697 2718
rect 1710 2692 1713 2728
rect 1682 2668 1686 2671
rect 1662 2612 1665 2638
rect 1560 2603 1562 2607
rect 1566 2603 1569 2607
rect 1573 2603 1576 2607
rect 1598 2552 1601 2598
rect 1686 2582 1689 2658
rect 1710 2652 1713 2668
rect 1718 2662 1721 2688
rect 1726 2672 1729 2798
rect 1734 2792 1737 2818
rect 1742 2772 1745 2868
rect 1750 2832 1753 2838
rect 1750 2762 1753 2828
rect 1734 2742 1737 2748
rect 1742 2682 1745 2748
rect 1750 2732 1753 2748
rect 1758 2732 1761 3268
rect 1766 3192 1769 3308
rect 1774 3242 1777 3248
rect 1766 3152 1769 3168
rect 1782 3102 1785 3358
rect 1814 3352 1817 3388
rect 1826 3378 1830 3381
rect 1834 3368 1838 3371
rect 1802 3348 1806 3351
rect 1814 3312 1817 3338
rect 1802 3268 1806 3271
rect 1794 3258 1798 3261
rect 1806 3252 1809 3258
rect 1782 3092 1785 3098
rect 1806 3062 1809 3078
rect 1766 3052 1769 3058
rect 1766 2992 1769 3038
rect 1822 3032 1825 3308
rect 1854 3272 1857 3338
rect 1838 3252 1841 3259
rect 1862 3162 1865 3418
rect 1918 3352 1921 3408
rect 1934 3392 1937 3458
rect 1874 3348 1878 3351
rect 1902 3342 1905 3348
rect 1934 3292 1937 3338
rect 1914 3268 1918 3271
rect 1830 3122 1833 3147
rect 1846 3132 1849 3138
rect 1862 3102 1865 3138
rect 1886 3132 1889 3148
rect 1902 3142 1905 3148
rect 1910 3122 1913 3138
rect 1878 3081 1881 3118
rect 1878 3078 1889 3081
rect 1830 3062 1833 3078
rect 1846 3072 1849 3078
rect 1886 3071 1889 3078
rect 1918 3072 1921 3218
rect 1942 3152 1945 3438
rect 1998 3422 2001 3448
rect 1974 3392 1977 3398
rect 1998 3372 2001 3418
rect 1950 3352 1953 3368
rect 2006 3362 2009 3658
rect 2038 3652 2041 3718
rect 2062 3552 2065 3718
rect 2072 3703 2074 3707
rect 2078 3703 2081 3707
rect 2085 3703 2088 3707
rect 2134 3672 2137 3698
rect 2150 3672 2153 3678
rect 2198 3672 2201 3708
rect 2114 3659 2118 3662
rect 2166 3662 2169 3668
rect 2158 3652 2161 3658
rect 2186 3648 2190 3651
rect 2114 3568 2118 3571
rect 2050 3548 2054 3551
rect 2014 3512 2017 3548
rect 2030 3542 2033 3548
rect 2030 3522 2033 3528
rect 2014 3472 2017 3508
rect 2062 3492 2065 3538
rect 2094 3522 2097 3538
rect 2072 3503 2074 3507
rect 2078 3503 2081 3507
rect 2085 3503 2088 3507
rect 2034 3488 2038 3491
rect 2126 3482 2129 3608
rect 2138 3558 2142 3561
rect 2146 3558 2150 3561
rect 2166 3552 2169 3618
rect 2178 3568 2182 3571
rect 2154 3548 2158 3551
rect 2082 3468 2086 3471
rect 2014 3442 2017 3458
rect 2022 3352 2025 3468
rect 2062 3462 2065 3468
rect 2094 3458 2102 3461
rect 2038 3452 2041 3458
rect 2030 3442 2033 3448
rect 2038 3372 2041 3378
rect 2046 3351 2049 3458
rect 2054 3442 2057 3448
rect 2062 3442 2065 3458
rect 2082 3448 2086 3451
rect 2094 3432 2097 3458
rect 2106 3448 2110 3451
rect 2134 3442 2137 3548
rect 2146 3538 2153 3541
rect 2142 3452 2145 3458
rect 2058 3358 2062 3361
rect 2046 3348 2057 3351
rect 1958 3282 1961 3348
rect 1954 3258 1958 3261
rect 1950 3192 1953 3248
rect 1958 3242 1961 3248
rect 1966 3162 1969 3338
rect 1974 3212 1977 3348
rect 2006 3272 2009 3348
rect 2030 3342 2033 3348
rect 2018 3338 2022 3341
rect 2038 3302 2041 3348
rect 2038 3282 2041 3298
rect 2054 3272 2057 3348
rect 2066 3338 2070 3341
rect 2014 3262 2017 3268
rect 2054 3251 2057 3268
rect 2062 3262 2065 3308
rect 2072 3303 2074 3307
rect 2078 3303 2081 3307
rect 2085 3303 2088 3307
rect 2074 3268 2078 3271
rect 2066 3258 2070 3261
rect 2054 3248 2065 3251
rect 1962 3148 1966 3151
rect 1930 3138 1934 3141
rect 1942 3122 1945 3148
rect 1958 3082 1961 3088
rect 1886 3068 1897 3071
rect 1906 3068 1910 3071
rect 1838 3052 1841 3058
rect 1782 3002 1785 3018
rect 1766 2751 1769 2978
rect 1774 2972 1777 2998
rect 1782 2942 1785 2948
rect 1790 2942 1793 3028
rect 1854 3022 1857 3058
rect 1870 3032 1873 3068
rect 1878 3062 1881 3068
rect 1822 2992 1825 3018
rect 1798 2982 1801 2988
rect 1818 2958 1822 2961
rect 1834 2958 1838 2961
rect 1846 2952 1849 2958
rect 1802 2948 1806 2951
rect 1878 2951 1881 2978
rect 1822 2942 1825 2948
rect 1766 2748 1774 2751
rect 1766 2682 1769 2738
rect 1750 2662 1753 2668
rect 1782 2662 1785 2888
rect 1790 2872 1793 2938
rect 1822 2932 1825 2938
rect 1830 2932 1833 2948
rect 1830 2888 1838 2891
rect 1878 2891 1881 2928
rect 1870 2888 1881 2891
rect 1830 2872 1833 2888
rect 1790 2782 1793 2868
rect 1854 2862 1857 2868
rect 1798 2792 1801 2858
rect 1846 2852 1849 2858
rect 1870 2832 1873 2888
rect 1878 2852 1881 2858
rect 1790 2762 1793 2768
rect 1862 2762 1865 2818
rect 1886 2792 1889 3058
rect 1894 3052 1897 3068
rect 1942 3062 1945 3068
rect 1914 3058 1918 3061
rect 1918 2992 1921 3058
rect 1926 3052 1929 3058
rect 1942 3042 1945 3048
rect 1910 2892 1913 2928
rect 1894 2862 1897 2868
rect 1902 2858 1918 2861
rect 1902 2852 1905 2858
rect 1926 2852 1929 2898
rect 1934 2892 1937 3008
rect 1942 2962 1945 2968
rect 1950 2872 1953 3018
rect 1966 2942 1969 3108
rect 1974 3092 1977 3118
rect 1982 2992 1985 3218
rect 2010 3148 2014 3151
rect 2014 3132 2017 3138
rect 1990 3012 1993 3058
rect 1998 3052 2001 3058
rect 2006 3032 2009 3058
rect 2014 3052 2017 3128
rect 2062 3122 2065 3248
rect 2094 3242 2097 3248
rect 2078 3162 2081 3168
rect 2090 3138 2094 3141
rect 2072 3103 2074 3107
rect 2078 3103 2081 3107
rect 2085 3103 2088 3107
rect 2070 3072 2073 3078
rect 2078 3062 2081 3068
rect 2034 3058 2038 3061
rect 2046 3042 2049 3048
rect 2054 3042 2057 3058
rect 2062 3022 2065 3058
rect 2094 3052 2097 3118
rect 2102 3082 2105 3338
rect 2134 3312 2137 3438
rect 2118 3262 2121 3308
rect 2150 3292 2153 3538
rect 2166 3522 2169 3548
rect 2190 3542 2193 3558
rect 2214 3542 2217 3618
rect 2230 3602 2233 3718
rect 2234 3548 2238 3551
rect 2262 3542 2265 3698
rect 2274 3668 2278 3671
rect 2286 3662 2289 3898
rect 2302 3862 2305 3888
rect 2310 3872 2313 4088
rect 2318 4062 2321 4068
rect 2326 3992 2329 4068
rect 2334 4032 2337 4058
rect 2342 4022 2345 4108
rect 2354 4068 2369 4071
rect 2366 4062 2369 4068
rect 2414 4062 2417 4118
rect 2446 4062 2449 4068
rect 2394 4058 2398 4061
rect 2434 4058 2438 4061
rect 2358 4052 2361 4058
rect 2350 4042 2353 4048
rect 2462 4042 2465 4218
rect 2486 4182 2489 4328
rect 2494 4282 2497 4348
rect 2502 4342 2505 4348
rect 2542 4342 2545 4348
rect 2630 4342 2633 4347
rect 2514 4338 2518 4341
rect 2566 4332 2569 4338
rect 2558 4322 2561 4328
rect 2494 4242 2497 4278
rect 2518 4242 2521 4259
rect 2470 4152 2473 4158
rect 2478 4152 2481 4168
rect 2486 4152 2489 4178
rect 2478 4142 2481 4148
rect 2374 4002 2377 4018
rect 2354 3968 2358 3971
rect 2342 3952 2345 3968
rect 2390 3952 2393 3968
rect 2414 3952 2417 3968
rect 2366 3932 2369 3948
rect 2374 3942 2377 3948
rect 2318 3922 2321 3928
rect 2342 3872 2345 3878
rect 2330 3868 2334 3871
rect 2310 3822 2313 3868
rect 2374 3862 2377 3878
rect 2318 3812 2321 3858
rect 2330 3848 2334 3851
rect 2342 3842 2345 3858
rect 2374 3852 2377 3858
rect 2354 3848 2358 3851
rect 2318 3702 2321 3738
rect 2330 3668 2334 3671
rect 2310 3662 2313 3668
rect 2322 3658 2326 3661
rect 2334 3642 2337 3658
rect 2294 3602 2297 3618
rect 2342 3592 2345 3838
rect 2382 3812 2385 3948
rect 2402 3918 2406 3921
rect 2422 3912 2425 4018
rect 2462 3982 2465 4018
rect 2462 3952 2465 3978
rect 2470 3931 2473 4108
rect 2486 4031 2489 4148
rect 2498 4118 2502 4121
rect 2518 4072 2521 4088
rect 2526 4082 2529 4198
rect 2534 4152 2537 4158
rect 2542 4092 2545 4238
rect 2574 4162 2577 4318
rect 2590 4282 2593 4338
rect 2690 4318 2694 4321
rect 2658 4288 2662 4291
rect 2662 4262 2665 4268
rect 2598 4232 2601 4258
rect 2678 4252 2681 4318
rect 2702 4302 2705 4338
rect 2710 4291 2713 4318
rect 2718 4312 2721 4338
rect 2734 4312 2737 4348
rect 2710 4288 2718 4291
rect 2686 4282 2689 4288
rect 2702 4262 2705 4268
rect 2710 4262 2713 4268
rect 2742 4262 2745 4468
rect 2774 4462 2777 4468
rect 2750 4412 2753 4428
rect 2758 4422 2761 4448
rect 2766 4351 2769 4428
rect 2782 4392 2785 4438
rect 2790 4422 2793 4458
rect 2798 4442 2801 4448
rect 2806 4392 2809 4468
rect 2814 4462 2817 4498
rect 2822 4472 2825 4508
rect 2870 4501 2873 4568
rect 2946 4558 2950 4561
rect 2974 4561 2977 4618
rect 2982 4592 2985 4648
rect 2990 4632 2993 4638
rect 3014 4622 3017 4658
rect 3022 4572 3025 4618
rect 3030 4592 3033 4708
rect 2974 4558 2982 4561
rect 3018 4558 3022 4561
rect 2990 4552 2993 4558
rect 3030 4552 3033 4558
rect 3026 4548 3030 4551
rect 2978 4538 2982 4541
rect 2966 4532 2969 4538
rect 2862 4498 2873 4501
rect 2834 4488 2838 4491
rect 2790 4362 2793 4368
rect 2762 4348 2769 4351
rect 2778 4348 2782 4351
rect 2794 4348 2798 4351
rect 2766 4338 2774 4341
rect 2730 4258 2734 4261
rect 2584 4203 2586 4207
rect 2590 4203 2593 4207
rect 2597 4203 2600 4207
rect 2670 4162 2673 4218
rect 2626 4158 2630 4161
rect 2682 4158 2686 4161
rect 2614 4142 2617 4148
rect 2566 4072 2569 4098
rect 2542 4052 2545 4068
rect 2462 3928 2473 3931
rect 2478 4028 2489 4031
rect 2430 3922 2433 3928
rect 2434 3918 2438 3921
rect 2418 3878 2422 3881
rect 2462 3862 2465 3928
rect 2470 3882 2473 3918
rect 2418 3858 2422 3861
rect 2434 3858 2438 3861
rect 2398 3822 2401 3858
rect 2410 3848 2414 3851
rect 2442 3828 2446 3831
rect 2350 3751 2353 3768
rect 2382 3752 2385 3788
rect 2390 3772 2393 3778
rect 2414 3752 2417 3758
rect 2426 3738 2430 3741
rect 2366 3732 2369 3738
rect 2382 3722 2385 3738
rect 2438 3722 2441 3758
rect 2478 3752 2481 4028
rect 2538 4018 2542 4021
rect 2486 3882 2489 3958
rect 2494 3911 2497 3947
rect 2510 3932 2513 3938
rect 2526 3932 2529 4018
rect 2558 4012 2561 4058
rect 2538 3988 2542 3991
rect 2494 3908 2505 3911
rect 2502 3892 2505 3908
rect 2486 3862 2489 3878
rect 2510 3872 2513 3878
rect 2518 3872 2521 3898
rect 2534 3862 2537 3878
rect 2518 3762 2521 3858
rect 2542 3822 2545 3948
rect 2574 3942 2577 4138
rect 2606 4132 2609 4138
rect 2670 4132 2673 4148
rect 2654 4112 2657 4118
rect 2582 4072 2585 4078
rect 2614 4072 2617 4098
rect 2650 4068 2654 4071
rect 2586 4038 2590 4041
rect 2584 4003 2586 4007
rect 2590 4003 2593 4007
rect 2597 4003 2600 4007
rect 2598 3952 2601 3978
rect 2598 3942 2601 3948
rect 2606 3932 2609 4058
rect 2638 4052 2641 4068
rect 2678 4062 2681 4148
rect 2694 4132 2697 4218
rect 2702 4212 2705 4258
rect 2710 4152 2713 4258
rect 2726 4242 2729 4248
rect 2750 4232 2753 4278
rect 2726 4192 2729 4228
rect 2750 4162 2753 4168
rect 2750 4152 2753 4158
rect 2722 4148 2726 4151
rect 2686 4122 2689 4128
rect 2702 4122 2705 4148
rect 2766 4142 2769 4338
rect 2806 4321 2809 4388
rect 2814 4372 2817 4458
rect 2822 4392 2825 4398
rect 2846 4352 2849 4388
rect 2814 4332 2817 4348
rect 2834 4338 2838 4341
rect 2806 4318 2817 4321
rect 2814 4262 2817 4318
rect 2854 4292 2857 4338
rect 2782 4252 2785 4259
rect 2782 4192 2785 4208
rect 2806 4162 2809 4228
rect 2794 4148 2798 4151
rect 2710 4132 2713 4138
rect 2766 4132 2769 4138
rect 2774 4102 2777 4128
rect 2758 4072 2761 4088
rect 2774 4072 2777 4098
rect 2622 4042 2625 4048
rect 2570 3918 2577 3921
rect 2558 3862 2561 3898
rect 2566 3852 2569 3858
rect 2458 3748 2462 3751
rect 2446 3742 2449 3748
rect 2374 3672 2377 3698
rect 2398 3692 2401 3718
rect 2358 3662 2361 3668
rect 2366 3652 2369 3658
rect 2310 3552 2313 3568
rect 2286 3542 2289 3548
rect 2174 3532 2177 3538
rect 2158 3462 2161 3498
rect 2166 3462 2169 3488
rect 2174 3452 2177 3458
rect 2158 3402 2161 3418
rect 2158 3351 2161 3368
rect 2190 3362 2193 3538
rect 2222 3472 2225 3538
rect 2218 3458 2222 3461
rect 2202 3368 2206 3371
rect 2218 3358 2222 3361
rect 2190 3352 2193 3358
rect 2174 3342 2177 3348
rect 2194 3338 2198 3341
rect 2214 3312 2217 3338
rect 2130 3268 2134 3271
rect 2166 3262 2169 3298
rect 2182 3262 2185 3268
rect 2134 3252 2137 3258
rect 2150 3232 2153 3238
rect 2110 3152 2113 3158
rect 2126 3152 2129 3168
rect 2110 3132 2113 3148
rect 2134 3142 2137 3148
rect 2150 3142 2153 3168
rect 2158 3152 2161 3188
rect 2222 3182 2225 3358
rect 2230 3352 2233 3538
rect 2278 3472 2281 3498
rect 2326 3462 2329 3588
rect 2374 3552 2377 3668
rect 2382 3592 2385 3658
rect 2398 3652 2401 3678
rect 2462 3672 2465 3738
rect 2474 3718 2478 3721
rect 2442 3658 2446 3661
rect 2398 3612 2401 3648
rect 2454 3592 2457 3638
rect 2462 3572 2465 3658
rect 2390 3552 2393 3558
rect 2334 3472 2337 3548
rect 2398 3542 2401 3568
rect 2414 3542 2417 3548
rect 2370 3538 2374 3541
rect 2370 3518 2374 3521
rect 2346 3488 2350 3491
rect 2422 3472 2425 3568
rect 2450 3548 2454 3551
rect 2474 3538 2478 3541
rect 2486 3532 2489 3748
rect 2518 3742 2521 3748
rect 2502 3732 2505 3738
rect 2514 3668 2518 3671
rect 2534 3662 2537 3798
rect 2550 3742 2553 3778
rect 2574 3762 2577 3918
rect 2594 3858 2598 3861
rect 2606 3842 2609 3928
rect 2614 3882 2617 4018
rect 2630 3962 2633 4018
rect 2638 3992 2641 4008
rect 2630 3922 2633 3947
rect 2646 3942 2649 4058
rect 2742 4052 2745 4059
rect 2674 4048 2678 4051
rect 2682 4018 2686 4021
rect 2654 3992 2657 4018
rect 2662 3962 2665 3968
rect 2674 3948 2678 3951
rect 2622 3862 2625 3878
rect 2630 3862 2633 3868
rect 2646 3862 2649 3868
rect 2584 3803 2586 3807
rect 2590 3803 2593 3807
rect 2597 3803 2600 3807
rect 2606 3792 2609 3818
rect 2630 3812 2633 3858
rect 2630 3792 2633 3798
rect 2594 3758 2598 3761
rect 2570 3738 2574 3741
rect 2610 3738 2614 3741
rect 2542 3662 2545 3668
rect 2550 3662 2553 3688
rect 2566 3672 2569 3698
rect 2574 3682 2577 3688
rect 2522 3658 2526 3661
rect 2430 3522 2433 3528
rect 2298 3458 2302 3461
rect 2402 3459 2406 3462
rect 2270 3442 2273 3448
rect 2286 3442 2289 3458
rect 2314 3448 2318 3451
rect 2254 3421 2257 3438
rect 2246 3418 2257 3421
rect 2230 3312 2233 3348
rect 2230 3272 2233 3308
rect 2238 3302 2241 3338
rect 2238 3262 2241 3278
rect 2214 3152 2217 3158
rect 2246 3152 2249 3418
rect 2302 3362 2305 3368
rect 2270 3352 2273 3358
rect 2258 3338 2262 3341
rect 2270 3202 2273 3348
rect 2286 3342 2289 3348
rect 2278 3332 2281 3338
rect 2278 3212 2281 3288
rect 2318 3282 2321 3448
rect 2438 3442 2441 3468
rect 2446 3462 2449 3498
rect 2454 3462 2457 3468
rect 2446 3452 2449 3458
rect 2470 3452 2473 3488
rect 2426 3368 2430 3371
rect 2330 3358 2334 3361
rect 2366 3351 2369 3358
rect 2326 3292 2329 3348
rect 2334 3342 2337 3348
rect 2310 3272 2313 3278
rect 2290 3268 2294 3271
rect 2306 3258 2310 3261
rect 2326 3242 2329 3248
rect 2290 3238 2294 3241
rect 2170 3148 2174 3151
rect 2206 3142 2209 3148
rect 2246 3142 2249 3148
rect 2254 3142 2257 3148
rect 2194 3138 2198 3141
rect 2182 3122 2185 3128
rect 2126 3092 2129 3118
rect 2130 3068 2134 3071
rect 2154 3068 2158 3071
rect 2266 3068 2270 3071
rect 2022 2992 2025 3018
rect 2006 2952 2009 2968
rect 1998 2942 2001 2948
rect 2014 2942 2017 2978
rect 2030 2952 2033 2958
rect 2038 2952 2041 2978
rect 2102 2951 2105 2958
rect 1958 2902 1961 2918
rect 1966 2892 1969 2938
rect 1998 2932 2001 2938
rect 2070 2932 2073 2948
rect 2014 2892 2017 2928
rect 2072 2903 2074 2907
rect 2078 2903 2081 2907
rect 2085 2903 2088 2907
rect 1942 2862 1945 2868
rect 1958 2862 1961 2888
rect 1910 2842 1913 2848
rect 1854 2752 1857 2758
rect 1842 2748 1846 2751
rect 1790 2742 1793 2748
rect 1726 2652 1729 2658
rect 1734 2612 1737 2648
rect 1702 2592 1705 2598
rect 1686 2572 1689 2578
rect 1674 2558 1678 2561
rect 1742 2561 1745 2618
rect 1742 2558 1753 2561
rect 1702 2552 1705 2558
rect 1574 2542 1577 2548
rect 1662 2542 1665 2548
rect 1742 2542 1745 2548
rect 1654 2512 1657 2518
rect 1574 2492 1577 2508
rect 1598 2482 1601 2488
rect 1546 2458 1550 2461
rect 1534 2448 1545 2451
rect 1382 2382 1385 2418
rect 1422 2392 1425 2428
rect 1358 2352 1361 2368
rect 1322 2348 1326 2351
rect 1302 2342 1305 2348
rect 1294 2281 1297 2338
rect 1334 2281 1337 2348
rect 1346 2338 1350 2341
rect 1294 2278 1305 2281
rect 1334 2278 1342 2281
rect 1262 2252 1265 2278
rect 1302 2272 1305 2278
rect 1366 2272 1369 2378
rect 1398 2352 1401 2368
rect 1406 2352 1409 2388
rect 1450 2368 1454 2371
rect 1446 2352 1449 2368
rect 1374 2348 1382 2351
rect 1374 2312 1377 2348
rect 1390 2342 1393 2348
rect 1430 2332 1433 2348
rect 1290 2268 1294 2271
rect 1306 2258 1310 2261
rect 1282 2248 1286 2251
rect 1294 2242 1297 2258
rect 1278 2152 1281 2158
rect 1286 2152 1289 2178
rect 1294 2142 1297 2228
rect 1302 2192 1305 2238
rect 1314 2218 1318 2221
rect 1314 2148 1318 2151
rect 1270 2132 1273 2138
rect 1326 2122 1329 2268
rect 1430 2262 1433 2308
rect 1334 2242 1337 2258
rect 1342 2192 1345 2258
rect 1350 2172 1353 2188
rect 1366 2182 1369 2218
rect 1358 2152 1361 2168
rect 1366 2152 1369 2158
rect 1246 2092 1249 2118
rect 1226 2088 1230 2091
rect 1154 2058 1158 2061
rect 1190 2032 1193 2058
rect 1206 2042 1209 2058
rect 1182 1992 1185 2008
rect 1158 1952 1161 1958
rect 1098 1948 1102 1951
rect 1058 1938 1062 1941
rect 1022 1888 1033 1891
rect 1022 1872 1025 1878
rect 982 1862 985 1868
rect 1030 1862 1033 1888
rect 1010 1858 1014 1861
rect 1038 1852 1041 1918
rect 1048 1903 1050 1907
rect 1054 1903 1057 1907
rect 1061 1903 1064 1907
rect 1062 1852 1065 1888
rect 974 1848 982 1851
rect 994 1848 998 1851
rect 950 1712 953 1748
rect 958 1742 961 1748
rect 958 1692 961 1718
rect 966 1692 969 1758
rect 982 1732 985 1738
rect 998 1711 1001 1747
rect 990 1708 1001 1711
rect 926 1682 929 1688
rect 930 1668 934 1671
rect 942 1662 945 1688
rect 862 1652 865 1659
rect 966 1652 969 1678
rect 982 1672 985 1698
rect 990 1692 993 1708
rect 1006 1662 1009 1818
rect 1070 1752 1073 1948
rect 1142 1942 1145 1948
rect 1090 1918 1094 1921
rect 1158 1881 1161 1948
rect 1166 1942 1169 1948
rect 1190 1942 1193 1948
rect 1154 1878 1161 1881
rect 1078 1852 1081 1858
rect 1086 1822 1089 1858
rect 1026 1738 1030 1741
rect 1086 1732 1089 1758
rect 1094 1732 1097 1868
rect 1126 1852 1129 1859
rect 1126 1828 1134 1831
rect 1102 1752 1105 1818
rect 1118 1792 1121 1808
rect 1118 1752 1121 1788
rect 1114 1738 1118 1741
rect 1030 1692 1033 1728
rect 1048 1703 1050 1707
rect 1054 1703 1057 1707
rect 1061 1703 1064 1707
rect 1070 1691 1073 1718
rect 1062 1688 1073 1691
rect 1054 1672 1057 1688
rect 1062 1682 1065 1688
rect 1102 1682 1105 1738
rect 1018 1668 1022 1671
rect 1050 1668 1054 1671
rect 1038 1662 1041 1668
rect 954 1648 958 1651
rect 934 1592 937 1648
rect 870 1552 873 1568
rect 898 1548 902 1551
rect 838 1542 841 1547
rect 878 1542 881 1548
rect 890 1538 894 1541
rect 790 1472 793 1528
rect 830 1472 833 1538
rect 878 1482 881 1538
rect 754 1468 758 1471
rect 770 1468 774 1471
rect 718 1462 721 1468
rect 790 1462 793 1468
rect 810 1458 814 1461
rect 850 1459 854 1462
rect 742 1422 745 1448
rect 734 1352 737 1388
rect 758 1362 761 1388
rect 726 1342 729 1348
rect 774 1342 777 1348
rect 782 1342 785 1448
rect 798 1432 801 1458
rect 878 1452 881 1458
rect 806 1448 814 1451
rect 806 1392 809 1448
rect 906 1418 910 1421
rect 830 1372 833 1418
rect 846 1362 849 1368
rect 854 1362 857 1398
rect 870 1362 873 1368
rect 906 1358 910 1361
rect 806 1352 809 1358
rect 830 1342 833 1358
rect 918 1352 921 1548
rect 926 1542 929 1558
rect 982 1552 985 1658
rect 994 1648 998 1651
rect 1006 1592 1009 1648
rect 1002 1558 1006 1561
rect 1014 1561 1017 1658
rect 1022 1582 1025 1648
rect 1038 1572 1041 1658
rect 1046 1592 1049 1648
rect 1102 1592 1105 1668
rect 1110 1662 1113 1708
rect 1110 1632 1113 1648
rect 1010 1558 1017 1561
rect 1022 1552 1025 1558
rect 954 1548 958 1551
rect 994 1548 998 1551
rect 1050 1548 1054 1551
rect 1030 1542 1033 1548
rect 946 1538 958 1541
rect 974 1532 977 1538
rect 1014 1522 1017 1538
rect 934 1472 937 1498
rect 966 1492 969 1508
rect 1048 1503 1050 1507
rect 1054 1503 1057 1507
rect 1061 1503 1064 1507
rect 942 1462 945 1468
rect 954 1458 958 1461
rect 982 1452 985 1468
rect 1010 1458 1014 1461
rect 1070 1452 1073 1578
rect 1082 1548 1086 1551
rect 1118 1542 1121 1728
rect 1126 1562 1129 1828
rect 1134 1682 1137 1718
rect 1150 1642 1153 1858
rect 1174 1792 1177 1938
rect 1206 1932 1209 1948
rect 1186 1888 1190 1891
rect 1214 1872 1217 2078
rect 1234 2068 1238 2071
rect 1238 2052 1241 2058
rect 1230 1952 1233 2028
rect 1230 1912 1233 1948
rect 1202 1868 1206 1871
rect 1226 1868 1230 1871
rect 1202 1858 1206 1861
rect 1214 1812 1217 1868
rect 1238 1862 1241 2048
rect 1254 1961 1257 2118
rect 1270 2082 1273 2088
rect 1294 2062 1297 2068
rect 1302 2062 1305 2118
rect 1310 2072 1313 2078
rect 1326 2072 1329 2118
rect 1266 2058 1270 2061
rect 1286 2052 1289 2058
rect 1270 2042 1273 2048
rect 1310 2042 1313 2058
rect 1250 1958 1257 1961
rect 1278 1942 1281 2018
rect 1302 1968 1310 1971
rect 1286 1952 1289 1958
rect 1294 1952 1297 1958
rect 1302 1952 1305 1968
rect 1310 1952 1313 1958
rect 1298 1938 1302 1941
rect 1278 1912 1281 1918
rect 1226 1858 1230 1861
rect 1226 1848 1230 1851
rect 1238 1842 1241 1848
rect 1254 1842 1257 1848
rect 1218 1788 1222 1791
rect 1158 1752 1161 1758
rect 1238 1752 1241 1798
rect 1246 1752 1249 1808
rect 1262 1782 1265 1868
rect 1178 1748 1182 1751
rect 1222 1748 1230 1751
rect 1198 1702 1201 1748
rect 1206 1742 1209 1748
rect 1170 1678 1174 1681
rect 1190 1672 1193 1688
rect 1206 1662 1209 1688
rect 1182 1652 1185 1658
rect 1170 1638 1174 1641
rect 1142 1542 1145 1548
rect 1150 1542 1153 1638
rect 1174 1592 1177 1628
rect 1190 1582 1193 1658
rect 1206 1602 1209 1658
rect 1214 1642 1217 1738
rect 1222 1692 1225 1748
rect 1254 1742 1257 1748
rect 1266 1738 1270 1741
rect 1278 1741 1281 1818
rect 1290 1748 1294 1751
rect 1278 1738 1286 1741
rect 1234 1668 1238 1671
rect 1246 1652 1249 1688
rect 1254 1671 1257 1738
rect 1274 1728 1278 1731
rect 1290 1728 1294 1731
rect 1262 1712 1265 1718
rect 1270 1692 1273 1718
rect 1302 1692 1305 1718
rect 1310 1692 1313 1948
rect 1318 1772 1321 2038
rect 1334 2022 1337 2148
rect 1374 2102 1377 2258
rect 1406 2252 1409 2259
rect 1394 2168 1398 2171
rect 1382 2142 1385 2148
rect 1342 2072 1345 2078
rect 1350 2062 1353 2098
rect 1366 2042 1369 2068
rect 1386 2059 1390 2062
rect 1346 2018 1350 2021
rect 1382 1982 1385 1988
rect 1334 1962 1337 1978
rect 1358 1952 1361 1958
rect 1386 1948 1390 1951
rect 1354 1938 1358 1941
rect 1366 1902 1369 1948
rect 1398 1942 1401 2158
rect 1414 2152 1417 2168
rect 1422 2162 1425 2198
rect 1406 2142 1409 2148
rect 1430 2042 1433 2258
rect 1438 2142 1441 2198
rect 1454 2172 1457 2238
rect 1462 2152 1465 2238
rect 1446 2142 1449 2148
rect 1446 2042 1449 2048
rect 1414 1932 1417 1998
rect 1454 1962 1457 2148
rect 1462 2082 1465 2088
rect 1430 1952 1433 1958
rect 1454 1942 1457 1948
rect 1470 1942 1473 2448
rect 1494 2312 1497 2348
rect 1518 2342 1521 2348
rect 1506 2288 1510 2291
rect 1478 2272 1481 2278
rect 1494 2272 1497 2288
rect 1486 2262 1489 2268
rect 1502 2152 1505 2278
rect 1514 2268 1518 2271
rect 1526 2262 1529 2418
rect 1542 2382 1545 2448
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1573 2403 1576 2407
rect 1582 2372 1585 2478
rect 1654 2472 1657 2478
rect 1662 2472 1665 2538
rect 1670 2482 1673 2488
rect 1678 2482 1681 2508
rect 1686 2492 1689 2498
rect 1702 2492 1705 2528
rect 1710 2502 1713 2538
rect 1726 2512 1729 2518
rect 1742 2492 1745 2508
rect 1674 2468 1678 2471
rect 1694 2462 1697 2488
rect 1706 2478 1710 2481
rect 1730 2478 1734 2481
rect 1750 2462 1753 2558
rect 1758 2492 1761 2518
rect 1758 2472 1761 2478
rect 1766 2472 1769 2628
rect 1774 2492 1777 2658
rect 1798 2651 1801 2718
rect 1806 2682 1809 2738
rect 1814 2722 1817 2748
rect 1822 2742 1825 2748
rect 1870 2742 1873 2758
rect 1882 2748 1886 2751
rect 1922 2747 1926 2750
rect 1822 2672 1825 2728
rect 1822 2652 1825 2668
rect 1854 2662 1857 2708
rect 1862 2672 1865 2738
rect 1886 2732 1889 2738
rect 1918 2722 1921 2728
rect 1894 2682 1897 2718
rect 1942 2692 1945 2708
rect 1950 2691 1953 2778
rect 1950 2688 1961 2691
rect 1950 2672 1953 2678
rect 1798 2648 1806 2651
rect 1790 2552 1793 2618
rect 1802 2578 1806 2581
rect 1822 2552 1825 2558
rect 1830 2552 1833 2618
rect 1838 2552 1841 2578
rect 1862 2552 1865 2588
rect 1894 2562 1897 2668
rect 1950 2662 1953 2668
rect 1958 2662 1961 2688
rect 1966 2662 1969 2798
rect 1974 2662 1977 2818
rect 1990 2812 1993 2858
rect 1998 2852 2001 2858
rect 1990 2752 1993 2758
rect 1990 2732 1993 2738
rect 2006 2732 2009 2748
rect 1982 2722 1985 2728
rect 2022 2682 2025 2898
rect 2074 2888 2078 2891
rect 2038 2872 2041 2888
rect 2094 2882 2097 2888
rect 2106 2858 2110 2861
rect 2030 2802 2033 2858
rect 2046 2852 2049 2858
rect 2046 2812 2049 2818
rect 2054 2792 2057 2798
rect 2030 2762 2033 2768
rect 2034 2748 2038 2751
rect 2034 2738 2038 2741
rect 2022 2672 2025 2678
rect 2062 2672 2065 2848
rect 2118 2832 2121 3058
rect 2126 3032 2129 3048
rect 2134 2972 2137 3048
rect 2142 3012 2145 3068
rect 2230 3052 2233 3059
rect 2134 2952 2137 2968
rect 2166 2952 2169 2968
rect 2182 2952 2185 2988
rect 2222 2952 2225 2978
rect 2230 2952 2233 3038
rect 2246 2972 2249 3068
rect 2262 2982 2265 3058
rect 2270 3042 2273 3048
rect 2174 2942 2177 2948
rect 2206 2942 2209 2948
rect 2158 2902 2161 2938
rect 2238 2932 2241 2938
rect 2246 2921 2249 2968
rect 2270 2962 2273 3008
rect 2278 2992 2281 3208
rect 2326 3182 2329 3238
rect 2318 3172 2321 3178
rect 2318 3162 2321 3168
rect 2334 3162 2337 3338
rect 2350 3281 2353 3348
rect 2366 3312 2369 3328
rect 2438 3302 2441 3318
rect 2342 3278 2353 3281
rect 2342 3262 2345 3278
rect 2358 3272 2361 3278
rect 2350 3232 2353 3268
rect 2378 3258 2382 3261
rect 2398 3252 2401 3298
rect 2438 3262 2441 3278
rect 2446 3262 2449 3418
rect 2462 3352 2465 3358
rect 2454 3332 2457 3338
rect 2478 3292 2481 3508
rect 2486 3342 2489 3528
rect 2494 3472 2497 3618
rect 2518 3612 2521 3648
rect 2514 3538 2518 3541
rect 2494 3452 2497 3458
rect 2502 3452 2505 3458
rect 2494 3342 2497 3438
rect 2502 3352 2505 3418
rect 2494 3292 2497 3338
rect 2502 3272 2505 3348
rect 2490 3258 2494 3261
rect 2430 3202 2433 3218
rect 2446 3172 2449 3258
rect 2502 3242 2505 3258
rect 2354 3158 2358 3161
rect 2366 3152 2369 3168
rect 2454 3162 2457 3188
rect 2446 3152 2449 3158
rect 2486 3152 2489 3198
rect 2502 3152 2505 3238
rect 2426 3148 2430 3151
rect 2338 3138 2342 3141
rect 2374 3122 2377 3128
rect 2306 3118 2310 3121
rect 2286 3052 2289 3058
rect 2294 3052 2297 3118
rect 2310 3072 2313 3078
rect 2350 3062 2353 3078
rect 2418 3068 2422 3071
rect 2310 3052 2313 3058
rect 2238 2918 2249 2921
rect 2154 2888 2158 2891
rect 2130 2868 2134 2871
rect 2134 2852 2137 2858
rect 2150 2822 2153 2868
rect 2134 2762 2137 2768
rect 2094 2752 2097 2758
rect 2086 2742 2089 2748
rect 2114 2738 2118 2741
rect 2072 2703 2074 2707
rect 2078 2703 2081 2707
rect 2085 2703 2088 2707
rect 2110 2682 2113 2688
rect 2038 2662 2041 2668
rect 2046 2662 2049 2668
rect 1930 2658 1934 2661
rect 2010 2658 2014 2661
rect 1958 2632 1961 2658
rect 1998 2652 2001 2658
rect 2078 2652 2081 2678
rect 2102 2662 2105 2668
rect 1898 2548 1902 2551
rect 1782 2542 1785 2548
rect 1814 2501 1817 2548
rect 1918 2542 1921 2588
rect 1934 2552 1937 2598
rect 1982 2561 1985 2618
rect 1974 2558 1985 2561
rect 1974 2552 1977 2558
rect 2022 2552 2025 2558
rect 1946 2548 1950 2551
rect 1986 2548 1990 2551
rect 2010 2548 2014 2551
rect 1926 2542 1929 2548
rect 1998 2542 2001 2548
rect 1882 2538 1886 2541
rect 1946 2538 1950 2541
rect 1814 2498 1825 2501
rect 1822 2492 1825 2498
rect 1810 2488 1814 2491
rect 1798 2472 1801 2488
rect 1830 2482 1833 2508
rect 1862 2492 1865 2518
rect 1830 2472 1833 2478
rect 1854 2472 1857 2478
rect 1618 2458 1622 2461
rect 1714 2458 1718 2461
rect 1794 2458 1798 2461
rect 1590 2442 1593 2458
rect 1622 2412 1625 2448
rect 1558 2342 1561 2368
rect 1582 2352 1585 2368
rect 1606 2362 1609 2368
rect 1622 2352 1625 2408
rect 1642 2368 1646 2371
rect 1626 2348 1630 2351
rect 1574 2292 1577 2328
rect 1582 2282 1585 2348
rect 1594 2338 1598 2341
rect 1622 2312 1625 2338
rect 1546 2268 1550 2271
rect 1590 2262 1593 2308
rect 1622 2262 1625 2268
rect 1486 2122 1489 2128
rect 1486 2062 1489 2068
rect 1494 2062 1497 2098
rect 1510 2092 1513 2248
rect 1526 2202 1529 2258
rect 1550 2252 1553 2258
rect 1598 2252 1601 2258
rect 1534 2248 1542 2251
rect 1526 2152 1529 2158
rect 1522 2138 1526 2141
rect 1534 2092 1537 2248
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1573 2203 1576 2207
rect 1542 2142 1545 2158
rect 1554 2118 1558 2121
rect 1502 2072 1505 2078
rect 1518 2072 1521 2088
rect 1550 2072 1553 2078
rect 1574 2062 1577 2098
rect 1582 2092 1585 2248
rect 1598 2152 1601 2168
rect 1598 2072 1601 2088
rect 1614 2081 1617 2218
rect 1630 2172 1633 2338
rect 1638 2332 1641 2338
rect 1646 2292 1649 2348
rect 1654 2342 1657 2418
rect 1702 2392 1705 2438
rect 1706 2388 1710 2391
rect 1718 2382 1721 2418
rect 1670 2362 1673 2368
rect 1666 2348 1670 2351
rect 1654 2312 1657 2338
rect 1686 2332 1689 2338
rect 1694 2322 1697 2328
rect 1670 2302 1673 2318
rect 1702 2292 1705 2378
rect 1710 2352 1713 2358
rect 1722 2348 1726 2351
rect 1734 2341 1737 2458
rect 1746 2448 1753 2451
rect 1750 2352 1753 2448
rect 1814 2442 1817 2448
rect 1822 2431 1825 2458
rect 1814 2428 1825 2431
rect 1734 2338 1742 2341
rect 1658 2268 1662 2271
rect 1682 2268 1686 2271
rect 1638 2222 1641 2248
rect 1662 2232 1665 2258
rect 1670 2252 1673 2268
rect 1694 2262 1697 2278
rect 1686 2212 1689 2218
rect 1694 2172 1697 2258
rect 1710 2252 1713 2338
rect 1722 2268 1726 2271
rect 1722 2258 1726 2261
rect 1734 2252 1737 2298
rect 1742 2292 1745 2318
rect 1750 2282 1753 2348
rect 1758 2302 1761 2318
rect 1750 2262 1753 2268
rect 1702 2242 1705 2248
rect 1746 2238 1750 2241
rect 1662 2162 1665 2168
rect 1622 2142 1625 2148
rect 1670 2112 1673 2128
rect 1614 2078 1625 2081
rect 1634 2078 1638 2081
rect 1586 2068 1590 2071
rect 1614 2062 1617 2068
rect 1622 2062 1625 2078
rect 1662 2072 1665 2108
rect 1678 2092 1681 2138
rect 1686 2101 1689 2158
rect 1710 2152 1713 2228
rect 1698 2118 1702 2121
rect 1686 2098 1697 2101
rect 1694 2092 1697 2098
rect 1710 2072 1713 2138
rect 1718 2092 1721 2118
rect 1726 2082 1729 2168
rect 1734 2152 1737 2168
rect 1742 2152 1745 2208
rect 1746 2138 1750 2141
rect 1750 2081 1753 2118
rect 1742 2078 1753 2081
rect 1758 2102 1761 2268
rect 1782 2262 1785 2268
rect 1790 2262 1793 2348
rect 1798 2342 1801 2348
rect 1798 2292 1801 2308
rect 1806 2282 1809 2298
rect 1814 2292 1817 2428
rect 1830 2392 1833 2468
rect 1870 2461 1873 2538
rect 1878 2472 1881 2478
rect 1866 2458 1873 2461
rect 1846 2442 1849 2448
rect 1854 2442 1857 2458
rect 1886 2452 1889 2518
rect 1894 2472 1897 2488
rect 1902 2471 1905 2498
rect 1910 2492 1913 2538
rect 1926 2482 1929 2518
rect 1934 2472 1937 2498
rect 1942 2472 1945 2518
rect 1902 2468 1910 2471
rect 1906 2458 1910 2461
rect 1866 2448 1870 2451
rect 1910 2448 1918 2451
rect 1854 2422 1857 2438
rect 1858 2368 1862 2371
rect 1822 2351 1825 2368
rect 1878 2352 1881 2448
rect 1890 2348 1894 2351
rect 1870 2332 1873 2338
rect 1854 2312 1857 2328
rect 1838 2272 1841 2278
rect 1846 2272 1849 2298
rect 1858 2278 1862 2281
rect 1870 2272 1873 2318
rect 1886 2312 1889 2328
rect 1774 2152 1777 2158
rect 1766 2102 1769 2138
rect 1782 2132 1785 2248
rect 1742 2072 1745 2078
rect 1538 2058 1545 2061
rect 1690 2058 1694 2061
rect 1738 2058 1742 2061
rect 1530 2048 1534 2051
rect 1542 2042 1545 2058
rect 1606 2052 1609 2058
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1573 2003 1576 2007
rect 1510 1992 1513 1998
rect 1502 1952 1505 1978
rect 1410 1918 1414 1921
rect 1430 1882 1433 1888
rect 1446 1872 1449 1878
rect 1470 1871 1473 1938
rect 1486 1932 1489 1938
rect 1486 1892 1489 1918
rect 1494 1872 1497 1888
rect 1470 1868 1478 1871
rect 1326 1862 1329 1868
rect 1342 1862 1345 1868
rect 1358 1852 1361 1859
rect 1366 1772 1369 1868
rect 1422 1842 1425 1868
rect 1502 1862 1505 1878
rect 1526 1862 1529 1898
rect 1534 1862 1537 1868
rect 1514 1858 1518 1861
rect 1418 1838 1422 1841
rect 1438 1832 1441 1838
rect 1470 1822 1473 1858
rect 1490 1848 1497 1851
rect 1318 1692 1321 1738
rect 1302 1682 1305 1688
rect 1334 1672 1337 1748
rect 1358 1722 1361 1748
rect 1366 1682 1369 1768
rect 1422 1752 1425 1758
rect 1398 1742 1401 1748
rect 1406 1742 1409 1748
rect 1430 1742 1433 1748
rect 1478 1741 1481 1838
rect 1474 1738 1481 1741
rect 1254 1668 1262 1671
rect 1262 1662 1265 1668
rect 1282 1658 1286 1661
rect 1190 1552 1193 1558
rect 1178 1548 1182 1551
rect 1118 1532 1121 1538
rect 1158 1522 1161 1548
rect 1198 1542 1201 1588
rect 1214 1572 1217 1638
rect 1230 1542 1233 1548
rect 1150 1472 1153 1488
rect 1166 1472 1169 1498
rect 1174 1492 1177 1498
rect 1174 1468 1198 1471
rect 934 1442 937 1448
rect 966 1442 969 1448
rect 966 1392 969 1398
rect 950 1352 953 1358
rect 974 1352 977 1358
rect 906 1348 910 1351
rect 938 1348 942 1351
rect 870 1342 873 1348
rect 746 1338 750 1341
rect 882 1338 886 1341
rect 798 1332 801 1338
rect 726 1292 729 1298
rect 678 1282 681 1288
rect 702 1282 705 1288
rect 638 1272 641 1278
rect 646 1262 649 1268
rect 654 1262 657 1268
rect 698 1258 702 1261
rect 562 1148 566 1151
rect 554 1138 558 1141
rect 574 1141 577 1148
rect 566 1138 577 1141
rect 510 1132 513 1138
rect 446 1128 454 1131
rect 426 1068 430 1071
rect 334 1042 337 1058
rect 342 942 345 1068
rect 350 1062 353 1068
rect 374 1052 377 1058
rect 398 1052 401 1058
rect 366 1042 369 1048
rect 382 1042 385 1048
rect 350 1032 353 1038
rect 370 988 374 991
rect 390 972 393 998
rect 406 992 409 1068
rect 414 1042 417 1058
rect 430 1052 433 1058
rect 414 1012 417 1038
rect 446 1022 449 1128
rect 462 1082 465 1128
rect 502 1122 505 1128
rect 486 1092 489 1118
rect 462 1063 465 1068
rect 358 942 361 958
rect 370 948 374 951
rect 342 882 345 908
rect 306 868 310 871
rect 318 862 321 868
rect 326 862 329 868
rect 278 762 281 818
rect 246 748 254 751
rect 238 742 241 748
rect 222 738 230 741
rect 206 732 209 738
rect 214 682 217 718
rect 222 692 225 738
rect 230 692 233 728
rect 202 678 206 681
rect 190 662 193 668
rect 206 652 209 668
rect 214 662 217 668
rect 174 592 177 648
rect 238 582 241 648
rect 230 572 233 578
rect 150 482 153 548
rect 158 521 161 538
rect 166 532 169 538
rect 182 532 185 558
rect 206 552 209 558
rect 194 548 198 551
rect 218 538 222 541
rect 198 522 201 538
rect 158 518 169 521
rect 70 392 73 438
rect 90 388 94 391
rect 102 342 105 348
rect 38 252 41 258
rect 38 152 41 158
rect 14 92 17 138
rect 62 132 65 138
rect 78 72 81 338
rect 102 272 105 278
rect 110 262 113 448
rect 118 352 121 418
rect 126 342 129 468
rect 150 462 153 468
rect 158 462 161 478
rect 166 472 169 518
rect 246 512 249 748
rect 286 742 289 858
rect 294 852 297 858
rect 350 792 353 838
rect 298 738 302 741
rect 254 672 257 678
rect 262 672 265 718
rect 294 712 297 738
rect 294 672 297 698
rect 358 672 361 938
rect 406 922 409 948
rect 414 942 417 978
rect 438 952 441 1008
rect 518 1002 521 1128
rect 566 1062 569 1138
rect 582 1122 585 1138
rect 630 1132 633 1158
rect 678 1152 681 1168
rect 686 1152 689 1248
rect 718 1182 721 1258
rect 758 1252 761 1258
rect 746 1168 750 1171
rect 726 1162 729 1168
rect 758 1162 761 1168
rect 766 1152 769 1158
rect 574 1102 577 1118
rect 582 1091 585 1118
rect 574 1088 585 1091
rect 574 1072 577 1088
rect 590 1072 593 1078
rect 534 1052 537 1058
rect 546 1048 550 1051
rect 536 1003 538 1007
rect 542 1003 545 1007
rect 549 1003 552 1007
rect 454 952 457 988
rect 502 972 505 988
rect 470 952 473 958
rect 498 948 502 951
rect 450 938 457 941
rect 474 938 478 941
rect 422 902 425 928
rect 430 872 433 918
rect 438 892 441 898
rect 374 842 377 868
rect 386 858 390 861
rect 402 858 406 861
rect 454 842 457 938
rect 486 922 489 948
rect 470 863 473 918
rect 510 902 513 958
rect 526 932 529 938
rect 478 862 481 868
rect 518 862 521 918
rect 518 772 521 838
rect 458 768 462 771
rect 494 762 497 768
rect 474 758 478 761
rect 398 752 401 758
rect 526 752 529 918
rect 534 892 537 988
rect 566 922 569 1058
rect 606 942 609 1068
rect 614 1062 617 1098
rect 630 1002 633 1118
rect 646 962 649 998
rect 662 961 665 1138
rect 670 1092 673 1148
rect 686 1082 689 1148
rect 734 1142 737 1148
rect 742 1102 745 1148
rect 686 1072 689 1078
rect 710 1062 713 1078
rect 730 1058 734 1061
rect 654 958 665 961
rect 614 942 617 947
rect 646 942 649 948
rect 550 882 553 918
rect 598 892 601 908
rect 570 888 574 891
rect 598 872 601 888
rect 590 862 593 868
rect 606 862 609 868
rect 614 862 617 918
rect 574 852 577 858
rect 630 852 633 878
rect 654 862 657 958
rect 666 948 670 951
rect 670 912 673 938
rect 678 932 681 988
rect 694 942 697 948
rect 702 942 705 948
rect 702 922 705 938
rect 642 858 646 861
rect 654 852 657 858
rect 662 842 665 868
rect 590 812 593 818
rect 536 803 538 807
rect 542 803 545 807
rect 549 803 552 807
rect 566 772 569 798
rect 586 758 590 761
rect 474 748 478 751
rect 462 742 465 748
rect 382 672 385 678
rect 398 672 401 738
rect 330 668 334 671
rect 330 658 334 661
rect 270 632 273 658
rect 286 642 289 648
rect 294 622 297 658
rect 322 648 326 651
rect 302 642 305 648
rect 258 578 262 581
rect 254 552 257 568
rect 270 552 273 618
rect 342 562 345 658
rect 350 642 353 648
rect 370 638 374 641
rect 358 592 361 638
rect 382 572 385 658
rect 422 642 425 658
rect 430 572 433 668
rect 446 652 449 708
rect 470 662 473 748
rect 590 742 593 748
rect 598 742 601 788
rect 678 772 681 868
rect 694 852 697 859
rect 694 792 697 798
rect 710 792 713 1028
rect 718 952 721 968
rect 718 872 721 948
rect 730 938 734 941
rect 742 792 745 848
rect 614 742 617 768
rect 630 751 633 758
rect 486 672 489 698
rect 518 682 521 738
rect 574 692 577 698
rect 598 692 601 728
rect 630 682 633 728
rect 582 672 585 678
rect 490 668 494 671
rect 518 662 521 668
rect 446 592 449 648
rect 478 642 481 648
rect 494 642 497 658
rect 514 648 518 651
rect 550 642 553 648
rect 262 541 265 548
rect 258 538 265 541
rect 310 542 313 548
rect 386 547 390 550
rect 462 542 465 638
rect 494 622 497 638
rect 536 603 538 607
rect 542 603 545 607
rect 549 603 552 607
rect 538 588 542 591
rect 478 551 481 558
rect 302 492 305 508
rect 342 472 345 538
rect 410 468 414 471
rect 426 468 430 471
rect 142 452 145 458
rect 158 442 161 448
rect 158 392 161 418
rect 166 392 169 468
rect 190 452 193 458
rect 174 432 177 438
rect 206 422 209 468
rect 222 442 225 459
rect 270 442 273 468
rect 318 462 321 468
rect 350 462 353 468
rect 410 458 414 461
rect 286 442 289 458
rect 178 348 182 351
rect 150 262 153 348
rect 174 332 177 338
rect 158 272 161 298
rect 94 242 97 258
rect 134 252 137 258
rect 110 242 113 248
rect 98 188 102 191
rect 134 152 137 168
rect 110 142 113 148
rect 142 72 145 258
rect 166 242 169 318
rect 182 302 185 348
rect 182 262 185 298
rect 190 272 193 328
rect 198 312 201 358
rect 218 348 222 351
rect 270 342 273 438
rect 278 352 281 378
rect 226 338 230 341
rect 230 322 233 338
rect 206 252 209 318
rect 286 312 289 428
rect 326 362 329 368
rect 334 342 337 458
rect 438 452 441 528
rect 502 522 505 538
rect 478 492 481 498
rect 502 472 505 518
rect 558 492 561 668
rect 566 632 569 658
rect 566 582 569 628
rect 590 602 593 678
rect 638 662 641 668
rect 654 662 657 768
rect 722 758 726 761
rect 686 702 689 758
rect 714 748 718 751
rect 702 732 705 738
rect 694 692 697 698
rect 702 672 705 718
rect 734 712 737 758
rect 750 742 753 1128
rect 774 1082 777 1328
rect 782 1302 785 1328
rect 790 1282 793 1318
rect 822 1262 825 1268
rect 790 1252 793 1259
rect 834 1258 838 1261
rect 830 1242 833 1248
rect 838 1222 841 1258
rect 846 1252 849 1318
rect 878 1292 881 1328
rect 894 1282 897 1288
rect 854 1272 857 1278
rect 866 1258 870 1261
rect 878 1212 881 1248
rect 878 1192 881 1198
rect 786 1168 790 1171
rect 794 1158 798 1161
rect 842 1148 846 1151
rect 790 1112 793 1138
rect 790 1062 793 1068
rect 782 992 785 998
rect 798 952 801 1148
rect 810 1138 814 1141
rect 806 1112 809 1118
rect 806 1082 809 1088
rect 810 1068 814 1071
rect 822 1062 825 1138
rect 806 992 809 1038
rect 822 972 825 1058
rect 830 1042 833 1068
rect 838 1062 841 1098
rect 846 1051 849 1108
rect 854 1092 857 1148
rect 870 1092 873 1168
rect 898 1148 902 1151
rect 886 1132 889 1148
rect 910 1141 913 1328
rect 926 1302 929 1348
rect 934 1312 937 1338
rect 950 1272 953 1318
rect 982 1282 985 1448
rect 1014 1392 1017 1448
rect 1030 1352 1033 1358
rect 1054 1352 1057 1448
rect 1066 1438 1070 1441
rect 1086 1382 1089 1468
rect 1118 1462 1121 1468
rect 1138 1458 1142 1461
rect 1094 1422 1097 1458
rect 1146 1448 1150 1451
rect 1110 1442 1113 1448
rect 1094 1372 1097 1378
rect 1078 1362 1081 1368
rect 1110 1362 1113 1368
rect 1018 1348 1022 1351
rect 1098 1348 1102 1351
rect 998 1332 1001 1348
rect 966 1272 969 1278
rect 990 1262 993 1268
rect 974 1192 977 1198
rect 1006 1192 1009 1208
rect 934 1152 937 1158
rect 946 1148 950 1151
rect 1010 1148 1014 1151
rect 902 1138 913 1141
rect 902 1092 905 1138
rect 942 1132 945 1138
rect 910 1122 913 1128
rect 858 1078 862 1081
rect 874 1068 878 1071
rect 886 1062 889 1068
rect 918 1062 921 1068
rect 934 1062 937 1128
rect 958 1112 961 1148
rect 946 1058 950 1061
rect 846 1048 854 1051
rect 902 1042 905 1048
rect 838 972 841 988
rect 818 948 822 951
rect 818 938 822 941
rect 758 882 761 888
rect 766 792 769 868
rect 774 862 777 928
rect 790 892 793 908
rect 798 882 801 928
rect 822 872 825 878
rect 830 872 833 948
rect 854 942 857 948
rect 838 892 841 928
rect 862 922 865 948
rect 870 942 873 1018
rect 918 972 921 1058
rect 962 988 966 991
rect 902 942 905 947
rect 918 942 921 968
rect 838 872 841 888
rect 870 881 873 938
rect 878 892 881 898
rect 894 892 897 898
rect 918 892 921 918
rect 974 892 977 958
rect 982 952 985 1148
rect 994 1138 998 1141
rect 1022 1141 1025 1158
rect 1014 1138 1025 1141
rect 1014 1092 1017 1138
rect 1030 1092 1033 1158
rect 1038 1152 1041 1348
rect 1078 1342 1081 1348
rect 1142 1342 1145 1347
rect 1050 1338 1054 1341
rect 1048 1303 1050 1307
rect 1054 1303 1057 1307
rect 1061 1303 1064 1307
rect 1050 1288 1054 1291
rect 1086 1272 1089 1338
rect 1074 1268 1078 1271
rect 1098 1268 1102 1271
rect 1110 1262 1113 1268
rect 1094 1222 1097 1258
rect 1110 1242 1113 1248
rect 1118 1192 1121 1308
rect 1126 1272 1129 1288
rect 1142 1282 1145 1328
rect 1158 1272 1161 1408
rect 1174 1312 1177 1468
rect 1198 1442 1201 1458
rect 1206 1452 1209 1458
rect 1202 1368 1206 1371
rect 1214 1362 1217 1518
rect 1254 1492 1257 1658
rect 1262 1542 1265 1548
rect 1226 1488 1230 1491
rect 1302 1472 1305 1668
rect 1374 1662 1377 1668
rect 1334 1652 1337 1658
rect 1318 1612 1321 1618
rect 1330 1588 1334 1591
rect 1314 1578 1318 1581
rect 1334 1572 1337 1578
rect 1362 1558 1366 1561
rect 1370 1558 1374 1561
rect 1318 1542 1321 1548
rect 1358 1501 1361 1548
rect 1374 1542 1377 1548
rect 1366 1532 1369 1538
rect 1358 1498 1369 1501
rect 1258 1468 1262 1471
rect 1302 1462 1305 1468
rect 1338 1458 1342 1461
rect 1238 1432 1241 1438
rect 1230 1362 1233 1388
rect 1246 1382 1249 1418
rect 1270 1412 1273 1418
rect 1266 1358 1270 1361
rect 1234 1348 1238 1351
rect 1218 1338 1222 1341
rect 1270 1332 1273 1338
rect 1254 1322 1257 1328
rect 1190 1292 1193 1308
rect 1166 1272 1169 1278
rect 1198 1272 1201 1278
rect 1206 1272 1209 1298
rect 1126 1252 1129 1268
rect 1138 1258 1142 1261
rect 1134 1242 1137 1248
rect 1078 1152 1081 1158
rect 1150 1152 1153 1158
rect 1158 1152 1161 1268
rect 1182 1262 1185 1268
rect 1214 1262 1217 1268
rect 1222 1262 1225 1268
rect 1170 1258 1177 1261
rect 1050 1148 1054 1151
rect 1054 1132 1057 1138
rect 1102 1128 1110 1131
rect 1048 1103 1050 1107
rect 1054 1103 1057 1107
rect 1061 1103 1064 1107
rect 1002 1088 1006 1091
rect 1070 1072 1073 1078
rect 1026 1068 1030 1071
rect 1046 1062 1049 1068
rect 1066 1058 1070 1061
rect 1002 1048 1006 1051
rect 1022 992 1025 1048
rect 994 938 998 941
rect 990 892 993 918
rect 862 878 873 881
rect 778 858 782 861
rect 786 848 790 851
rect 802 848 806 851
rect 806 822 809 828
rect 782 752 785 808
rect 802 758 806 761
rect 770 748 774 751
rect 758 702 761 728
rect 766 682 769 708
rect 762 678 766 681
rect 722 668 726 671
rect 714 658 718 661
rect 770 658 774 661
rect 590 572 593 598
rect 606 572 609 638
rect 574 552 577 568
rect 618 558 622 561
rect 630 552 633 558
rect 646 552 649 568
rect 618 548 622 551
rect 570 538 574 541
rect 606 538 614 541
rect 618 538 622 541
rect 598 492 601 498
rect 606 472 609 538
rect 630 502 633 548
rect 654 542 657 658
rect 726 642 729 648
rect 750 592 753 598
rect 814 592 817 748
rect 822 742 825 788
rect 846 762 849 818
rect 862 792 865 878
rect 982 872 985 888
rect 1006 882 1009 948
rect 1030 942 1033 968
rect 1062 952 1065 968
rect 1048 903 1050 907
rect 1054 903 1057 907
rect 1061 903 1064 907
rect 930 868 934 871
rect 870 862 873 868
rect 886 852 889 858
rect 910 852 913 868
rect 870 822 873 838
rect 894 802 897 848
rect 918 831 921 848
rect 914 828 921 831
rect 926 832 929 868
rect 966 852 969 858
rect 958 842 961 848
rect 938 838 942 841
rect 942 792 945 818
rect 838 752 841 758
rect 878 751 881 758
rect 830 732 833 748
rect 862 712 865 738
rect 822 661 825 698
rect 830 672 833 678
rect 886 672 889 768
rect 902 692 905 758
rect 910 672 913 678
rect 846 662 849 668
rect 918 662 921 668
rect 926 662 929 788
rect 950 762 953 798
rect 966 772 969 828
rect 966 742 969 768
rect 974 752 977 758
rect 950 732 953 738
rect 942 692 945 708
rect 966 672 969 718
rect 982 692 985 848
rect 990 792 993 878
rect 1006 862 1009 868
rect 1014 792 1017 868
rect 1030 772 1033 868
rect 1070 862 1073 868
rect 1078 792 1081 1128
rect 1094 1102 1097 1118
rect 1102 1092 1105 1128
rect 1090 1068 1094 1071
rect 1102 1052 1105 1088
rect 1118 1032 1121 1058
rect 1110 992 1113 998
rect 1126 981 1129 1148
rect 1162 1138 1166 1141
rect 1134 1082 1137 1118
rect 1134 1052 1137 1068
rect 1142 1042 1145 1048
rect 1150 1002 1153 1128
rect 1158 1052 1161 1058
rect 1166 1042 1169 1048
rect 1118 978 1129 981
rect 1118 962 1121 978
rect 1130 968 1134 971
rect 1118 942 1121 958
rect 1142 952 1145 988
rect 1150 972 1153 998
rect 1166 952 1169 1028
rect 1174 1022 1177 1258
rect 1230 1252 1233 1318
rect 1262 1263 1265 1268
rect 1278 1252 1281 1458
rect 1286 1452 1289 1458
rect 1366 1452 1369 1498
rect 1382 1481 1385 1738
rect 1446 1732 1449 1738
rect 1454 1692 1457 1728
rect 1434 1688 1438 1691
rect 1422 1552 1425 1688
rect 1462 1672 1465 1718
rect 1470 1712 1473 1738
rect 1486 1732 1489 1738
rect 1494 1732 1497 1848
rect 1502 1812 1505 1858
rect 1522 1848 1526 1851
rect 1542 1792 1545 1968
rect 1550 1892 1553 1968
rect 1562 1948 1566 1951
rect 1590 1942 1593 1948
rect 1614 1932 1617 2058
rect 1646 2012 1649 2058
rect 1670 2022 1673 2038
rect 1678 2002 1681 2048
rect 1686 1951 1689 1958
rect 1594 1888 1598 1891
rect 1598 1872 1601 1878
rect 1614 1872 1617 1918
rect 1638 1862 1641 1868
rect 1662 1862 1665 1948
rect 1562 1858 1566 1861
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1573 1803 1576 1807
rect 1526 1752 1529 1768
rect 1478 1662 1481 1668
rect 1442 1658 1446 1661
rect 1442 1648 1446 1651
rect 1434 1578 1438 1581
rect 1454 1562 1457 1658
rect 1486 1651 1489 1718
rect 1522 1688 1526 1691
rect 1542 1662 1545 1788
rect 1662 1772 1665 1858
rect 1550 1752 1553 1758
rect 1662 1752 1665 1768
rect 1658 1748 1662 1751
rect 1574 1742 1577 1748
rect 1610 1738 1614 1741
rect 1574 1672 1577 1738
rect 1498 1658 1502 1661
rect 1530 1658 1534 1661
rect 1486 1648 1494 1651
rect 1462 1592 1465 1648
rect 1510 1642 1513 1658
rect 1598 1652 1601 1658
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1573 1603 1576 1607
rect 1478 1562 1481 1588
rect 1438 1558 1446 1561
rect 1490 1558 1494 1561
rect 1402 1548 1406 1551
rect 1394 1538 1398 1541
rect 1406 1492 1409 1528
rect 1414 1492 1417 1498
rect 1382 1478 1393 1481
rect 1390 1472 1393 1478
rect 1422 1472 1425 1508
rect 1366 1422 1369 1448
rect 1386 1438 1390 1441
rect 1398 1412 1401 1458
rect 1414 1452 1417 1458
rect 1366 1392 1369 1398
rect 1346 1358 1350 1361
rect 1366 1352 1369 1358
rect 1406 1352 1409 1428
rect 1430 1402 1433 1498
rect 1438 1492 1441 1558
rect 1442 1458 1446 1461
rect 1442 1438 1446 1441
rect 1438 1362 1441 1398
rect 1454 1392 1457 1558
rect 1502 1552 1505 1588
rect 1534 1552 1537 1578
rect 1590 1552 1593 1558
rect 1554 1548 1558 1551
rect 1570 1548 1574 1551
rect 1470 1542 1473 1548
rect 1598 1542 1601 1548
rect 1494 1492 1497 1538
rect 1550 1532 1553 1538
rect 1522 1528 1526 1531
rect 1478 1472 1481 1488
rect 1502 1472 1505 1488
rect 1518 1481 1521 1508
rect 1510 1478 1521 1481
rect 1470 1462 1473 1468
rect 1510 1462 1513 1478
rect 1534 1462 1537 1488
rect 1462 1452 1465 1458
rect 1510 1452 1513 1458
rect 1486 1448 1494 1451
rect 1422 1352 1425 1358
rect 1434 1348 1438 1351
rect 1286 1312 1289 1348
rect 1294 1302 1297 1338
rect 1310 1292 1313 1348
rect 1334 1332 1337 1348
rect 1322 1318 1326 1321
rect 1342 1312 1345 1348
rect 1470 1342 1473 1347
rect 1366 1338 1374 1341
rect 1410 1338 1414 1341
rect 1334 1292 1337 1298
rect 1326 1282 1329 1288
rect 1342 1282 1345 1288
rect 1346 1268 1350 1271
rect 1358 1262 1361 1268
rect 1182 1132 1185 1248
rect 1190 1072 1193 1188
rect 1182 1032 1185 1038
rect 1130 948 1134 951
rect 1126 882 1129 888
rect 1022 762 1025 768
rect 990 752 993 758
rect 990 742 993 748
rect 998 732 1001 738
rect 986 668 990 671
rect 822 658 833 661
rect 822 642 825 648
rect 830 562 833 658
rect 778 558 782 561
rect 794 558 798 561
rect 686 551 689 558
rect 758 552 761 558
rect 770 538 774 541
rect 786 538 790 541
rect 818 538 822 541
rect 490 468 494 471
rect 454 462 457 468
rect 438 442 441 448
rect 402 438 406 441
rect 346 378 350 381
rect 358 352 361 358
rect 346 348 350 351
rect 366 342 369 388
rect 390 362 393 368
rect 378 358 382 361
rect 450 358 454 361
rect 334 332 337 338
rect 286 292 289 308
rect 222 282 225 288
rect 310 262 313 298
rect 366 292 369 338
rect 374 302 377 348
rect 390 301 393 348
rect 398 312 401 358
rect 382 298 393 301
rect 318 272 321 288
rect 222 252 225 259
rect 166 192 169 238
rect 182 162 185 218
rect 194 178 198 181
rect 194 158 198 161
rect 214 152 217 158
rect 202 148 206 151
rect 222 151 225 188
rect 294 182 297 238
rect 358 232 361 268
rect 382 261 385 298
rect 406 292 409 358
rect 414 352 417 358
rect 450 348 454 351
rect 462 342 465 468
rect 542 452 545 458
rect 470 432 473 448
rect 536 403 538 407
rect 542 403 545 407
rect 549 403 552 407
rect 598 382 601 418
rect 594 378 598 381
rect 502 372 505 378
rect 474 358 478 361
rect 434 338 438 341
rect 458 338 462 341
rect 422 322 425 338
rect 438 312 441 338
rect 422 292 425 308
rect 378 258 385 261
rect 430 261 433 298
rect 462 292 465 318
rect 470 302 473 348
rect 538 347 542 350
rect 606 341 609 468
rect 638 462 641 538
rect 646 492 649 538
rect 670 522 673 538
rect 654 472 657 478
rect 618 458 622 461
rect 634 448 638 451
rect 614 442 617 448
rect 614 392 617 398
rect 630 392 633 428
rect 654 362 657 468
rect 662 392 665 438
rect 622 352 625 358
rect 598 338 609 341
rect 618 338 622 341
rect 454 272 457 278
rect 442 268 446 271
rect 430 258 438 261
rect 422 252 425 258
rect 478 232 481 268
rect 502 262 505 268
rect 542 262 545 338
rect 566 262 569 298
rect 558 242 561 248
rect 230 152 233 158
rect 278 152 281 168
rect 286 162 289 168
rect 222 148 230 151
rect 258 148 262 151
rect 222 142 225 148
rect 238 142 241 148
rect 150 72 153 78
rect 158 72 161 138
rect 294 132 297 178
rect 310 172 313 218
rect 326 192 329 218
rect 306 148 310 151
rect 230 72 233 78
rect 246 63 249 118
rect 278 92 281 128
rect 310 122 313 138
rect 318 132 321 138
rect 358 132 361 228
rect 426 188 430 191
rect 370 148 374 151
rect 306 88 310 91
rect 326 72 329 78
rect 358 72 361 128
rect 406 92 409 168
rect 462 162 465 188
rect 494 172 497 218
rect 536 203 538 207
rect 542 203 545 207
rect 549 203 552 207
rect 494 162 497 168
rect 430 142 433 158
rect 510 152 513 178
rect 566 162 569 198
rect 450 148 454 151
rect 482 148 486 151
rect 438 132 441 148
rect 490 138 494 141
rect 522 138 526 141
rect 414 72 417 118
rect 210 58 214 61
rect 422 62 425 128
rect 454 72 457 78
rect 430 62 433 68
rect 478 62 481 78
rect 362 58 366 61
rect 438 52 441 58
rect 494 52 497 118
rect 542 112 545 138
rect 550 132 553 148
rect 574 142 577 298
rect 582 272 585 318
rect 598 302 601 338
rect 606 292 609 328
rect 646 292 649 358
rect 678 352 681 378
rect 686 352 689 518
rect 782 512 785 528
rect 750 482 753 488
rect 758 472 761 488
rect 830 482 833 548
rect 838 522 841 658
rect 866 648 870 651
rect 886 642 889 658
rect 894 652 897 658
rect 870 638 878 641
rect 846 592 849 638
rect 870 592 873 638
rect 886 572 889 638
rect 902 592 905 658
rect 950 592 953 648
rect 966 592 969 658
rect 978 648 982 651
rect 1006 632 1009 728
rect 1022 712 1025 718
rect 1030 701 1033 768
rect 1126 762 1129 858
rect 1134 812 1137 868
rect 1142 862 1145 948
rect 1166 922 1169 948
rect 1174 942 1177 948
rect 1190 932 1193 1058
rect 1206 992 1209 1218
rect 1214 1192 1217 1248
rect 1238 1192 1241 1238
rect 1242 1148 1246 1151
rect 1222 1042 1225 1059
rect 1230 1031 1233 1138
rect 1254 1132 1257 1158
rect 1286 1132 1289 1258
rect 1294 1142 1297 1148
rect 1250 1058 1254 1061
rect 1286 1061 1289 1128
rect 1294 1092 1297 1128
rect 1342 1082 1345 1198
rect 1366 1192 1369 1338
rect 1390 1332 1393 1338
rect 1382 1272 1385 1278
rect 1382 1252 1385 1258
rect 1374 1132 1377 1208
rect 1390 1192 1393 1328
rect 1402 1258 1406 1261
rect 1414 1252 1417 1258
rect 1422 1252 1425 1338
rect 1430 1292 1433 1298
rect 1486 1292 1489 1448
rect 1590 1442 1593 1468
rect 1494 1352 1497 1438
rect 1510 1402 1513 1418
rect 1526 1391 1529 1438
rect 1526 1388 1534 1391
rect 1482 1288 1486 1291
rect 1458 1278 1462 1281
rect 1470 1272 1473 1278
rect 1470 1262 1473 1268
rect 1398 1242 1401 1248
rect 1438 1242 1441 1258
rect 1494 1242 1497 1348
rect 1550 1342 1553 1418
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1573 1403 1576 1407
rect 1606 1392 1609 1698
rect 1614 1592 1617 1728
rect 1678 1672 1681 1778
rect 1686 1751 1689 1758
rect 1702 1732 1705 2048
rect 1726 2042 1729 2048
rect 1750 1992 1753 2068
rect 1758 2062 1761 2098
rect 1782 2072 1785 2128
rect 1790 2122 1793 2138
rect 1790 2062 1793 2078
rect 1798 2072 1801 2108
rect 1806 2092 1809 2218
rect 1814 2182 1817 2248
rect 1838 2222 1841 2258
rect 1830 2142 1833 2148
rect 1846 2142 1849 2268
rect 1862 2202 1865 2268
rect 1878 2262 1881 2298
rect 1886 2262 1889 2298
rect 1894 2292 1897 2318
rect 1902 2272 1905 2388
rect 1910 2322 1913 2448
rect 1930 2438 1934 2441
rect 1942 2432 1945 2448
rect 1946 2428 1950 2431
rect 1922 2368 1926 2371
rect 1958 2362 1961 2518
rect 1966 2492 1969 2538
rect 1990 2532 1993 2538
rect 1990 2472 1993 2508
rect 2006 2492 2009 2518
rect 2014 2492 2017 2538
rect 2006 2472 2009 2478
rect 1966 2392 1969 2428
rect 1974 2381 1977 2458
rect 1966 2378 1977 2381
rect 1926 2332 1929 2358
rect 1954 2348 1958 2351
rect 1918 2322 1921 2328
rect 1926 2312 1929 2328
rect 1934 2271 1937 2348
rect 1942 2342 1945 2348
rect 1942 2322 1945 2328
rect 1950 2302 1953 2318
rect 1950 2282 1953 2288
rect 1966 2282 1969 2378
rect 1990 2352 1993 2388
rect 2014 2372 2017 2458
rect 2022 2452 2025 2518
rect 2030 2492 2033 2638
rect 2054 2582 2057 2628
rect 2046 2542 2049 2548
rect 2054 2532 2057 2538
rect 2038 2472 2041 2518
rect 2062 2512 2065 2618
rect 2070 2562 2073 2598
rect 2126 2552 2129 2758
rect 2154 2748 2158 2751
rect 2174 2742 2177 2838
rect 2190 2782 2193 2918
rect 2238 2872 2241 2918
rect 2214 2862 2217 2868
rect 2238 2782 2241 2868
rect 2254 2862 2257 2918
rect 2262 2912 2265 2948
rect 2230 2762 2233 2768
rect 2226 2758 2230 2761
rect 2206 2752 2209 2758
rect 2230 2742 2233 2748
rect 2254 2742 2257 2768
rect 2158 2732 2161 2738
rect 2182 2732 2185 2738
rect 2190 2732 2193 2738
rect 2246 2732 2249 2738
rect 2166 2662 2169 2718
rect 2206 2692 2209 2698
rect 2242 2678 2246 2681
rect 2258 2678 2262 2681
rect 2190 2672 2193 2678
rect 2270 2672 2273 2958
rect 2294 2952 2297 2958
rect 2334 2952 2337 3008
rect 2314 2938 2318 2941
rect 2286 2932 2289 2938
rect 2278 2892 2281 2918
rect 2286 2812 2289 2858
rect 2294 2692 2297 2938
rect 2318 2912 2321 2918
rect 2314 2888 2318 2891
rect 2302 2882 2305 2888
rect 2314 2868 2318 2871
rect 2302 2852 2305 2858
rect 2334 2812 2337 2948
rect 2374 2942 2377 3058
rect 2430 3052 2433 3068
rect 2454 3062 2457 3098
rect 2470 3072 2473 3078
rect 2486 3072 2489 3098
rect 2502 3072 2505 3118
rect 2510 3112 2513 3528
rect 2534 3522 2537 3658
rect 2550 3642 2553 3658
rect 2582 3652 2585 3718
rect 2590 3712 2593 3738
rect 2610 3718 2614 3721
rect 2630 3692 2633 3718
rect 2638 3712 2641 3858
rect 2654 3792 2657 3918
rect 2670 3862 2673 3938
rect 2694 3862 2697 3988
rect 2702 3962 2705 4018
rect 2702 3932 2705 3958
rect 2718 3862 2721 4018
rect 2758 3992 2761 4058
rect 2726 3962 2729 3968
rect 2742 3962 2745 3968
rect 2774 3962 2777 4058
rect 2798 4042 2801 4048
rect 2786 3968 2790 3971
rect 2806 3961 2809 4118
rect 2814 4092 2817 4258
rect 2822 4142 2825 4208
rect 2838 4192 2841 4268
rect 2862 4262 2865 4498
rect 2878 4362 2881 4488
rect 2890 4468 2894 4471
rect 2898 4458 2902 4461
rect 2878 4332 2881 4338
rect 2846 4222 2849 4228
rect 2854 4202 2857 4258
rect 2870 4231 2873 4318
rect 2886 4262 2889 4378
rect 2910 4372 2913 4518
rect 2942 4512 2945 4518
rect 2942 4472 2945 4508
rect 2950 4452 2953 4458
rect 2958 4451 2961 4518
rect 2978 4468 2982 4471
rect 2998 4462 3001 4538
rect 2982 4452 2985 4458
rect 2958 4448 2966 4451
rect 3006 4451 3009 4518
rect 3022 4512 3025 4538
rect 3002 4448 3009 4451
rect 3038 4462 3041 4728
rect 3054 4652 3057 4718
rect 3070 4682 3073 4858
rect 3094 4792 3097 4848
rect 3126 4842 3129 4868
rect 3190 4862 3193 4928
rect 4112 4903 4114 4907
rect 4118 4903 4121 4907
rect 4125 4903 4128 4907
rect 3618 4888 3622 4891
rect 3986 4888 3990 4891
rect 5002 4888 5006 4891
rect 3830 4882 3833 4888
rect 4078 4882 4081 4888
rect 5166 4882 5169 4888
rect 3214 4872 3217 4878
rect 3342 4872 3345 4878
rect 3346 4868 3350 4871
rect 3226 4858 3230 4861
rect 3150 4842 3153 4858
rect 3254 4852 3257 4868
rect 3282 4858 3286 4861
rect 3362 4858 3366 4861
rect 3190 4842 3193 4848
rect 3222 4832 3225 4838
rect 3206 4782 3209 4818
rect 3222 4752 3225 4818
rect 3238 4772 3241 4848
rect 3318 4752 3321 4838
rect 3334 4802 3337 4818
rect 3110 4732 3113 4748
rect 3234 4748 3238 4751
rect 3338 4748 3342 4751
rect 3078 4692 3081 4718
rect 3096 4703 3098 4707
rect 3102 4703 3105 4707
rect 3109 4703 3112 4707
rect 3118 4692 3121 4718
rect 3142 4702 3145 4747
rect 3174 4742 3177 4748
rect 3210 4738 3214 4741
rect 3150 4682 3153 4688
rect 3158 4682 3161 4738
rect 3190 4732 3193 4738
rect 3062 4662 3065 4668
rect 3050 4648 3054 4651
rect 3062 4642 3065 4648
rect 3054 4572 3057 4598
rect 3058 4568 3062 4571
rect 2950 4432 2953 4438
rect 2894 4362 2897 4368
rect 2906 4318 2910 4321
rect 2894 4262 2897 4318
rect 2918 4262 2921 4328
rect 2934 4282 2937 4318
rect 2958 4262 2961 4418
rect 2966 4272 2969 4347
rect 2982 4302 2985 4418
rect 3006 4352 3009 4418
rect 2922 4258 2926 4261
rect 2962 4258 2966 4261
rect 2990 4252 2993 4258
rect 2918 4242 2921 4248
rect 2862 4228 2873 4231
rect 2846 4152 2849 4188
rect 2862 4162 2865 4228
rect 2850 4148 2854 4151
rect 2862 4142 2865 4148
rect 2822 4102 2825 4138
rect 2870 4102 2873 4218
rect 2878 4152 2881 4198
rect 2918 4152 2921 4168
rect 2834 4068 2838 4071
rect 2818 4058 2822 4061
rect 2826 4048 2830 4051
rect 2834 4038 2838 4041
rect 2830 3972 2833 3988
rect 2838 3962 2841 4038
rect 2802 3958 2809 3961
rect 2734 3951 2737 3958
rect 2814 3952 2817 3958
rect 2730 3948 2737 3951
rect 2726 3932 2729 3948
rect 2758 3942 2761 3948
rect 2734 3932 2737 3938
rect 2766 3922 2769 3938
rect 2774 3912 2777 3938
rect 2734 3872 2737 3878
rect 2758 3872 2761 3878
rect 2770 3868 2774 3871
rect 2782 3862 2785 3948
rect 2830 3942 2833 3958
rect 2854 3952 2857 4068
rect 2878 4002 2881 4148
rect 2902 4122 2905 4128
rect 2902 4082 2905 4088
rect 2894 4052 2897 4058
rect 2918 4052 2921 4148
rect 2926 4132 2929 4138
rect 2934 4092 2937 4158
rect 2946 4118 2950 4121
rect 2974 4092 2977 4248
rect 2998 4192 3001 4218
rect 2998 4142 3001 4148
rect 2982 4092 2985 4138
rect 3006 4102 3009 4348
rect 3022 4271 3025 4368
rect 3038 4342 3041 4458
rect 3054 4392 3057 4438
rect 3062 4402 3065 4458
rect 3046 4292 3049 4348
rect 3014 4268 3025 4271
rect 3042 4268 3046 4271
rect 3014 4262 3017 4268
rect 3022 4252 3025 4258
rect 3030 4222 3033 4258
rect 3054 4192 3057 4388
rect 3062 4262 3065 4268
rect 3038 4152 3041 4158
rect 3062 4142 3065 4258
rect 3070 4222 3073 4678
rect 3174 4672 3177 4718
rect 3182 4712 3185 4718
rect 3198 4712 3201 4728
rect 3182 4692 3185 4698
rect 3206 4691 3209 4718
rect 3214 4702 3217 4738
rect 3222 4722 3225 4748
rect 3254 4742 3257 4748
rect 3262 4742 3265 4748
rect 3206 4688 3217 4691
rect 3214 4672 3217 4688
rect 3230 4682 3233 4688
rect 3238 4672 3241 4738
rect 3294 4692 3297 4728
rect 3146 4668 3150 4671
rect 3078 4658 3086 4661
rect 3078 4582 3081 4658
rect 3086 4642 3089 4648
rect 3078 4552 3081 4578
rect 3086 4562 3089 4568
rect 3082 4538 3086 4541
rect 3094 4541 3097 4668
rect 3114 4648 3118 4651
rect 3134 4562 3137 4658
rect 3090 4538 3097 4541
rect 3154 4548 3158 4551
rect 3102 4542 3105 4548
rect 3142 4542 3145 4548
rect 3166 4542 3169 4658
rect 3174 4552 3177 4668
rect 3190 4662 3193 4668
rect 3230 4663 3233 4668
rect 3162 4538 3166 4541
rect 3086 4452 3089 4518
rect 3126 4512 3129 4528
rect 3096 4503 3098 4507
rect 3102 4503 3105 4507
rect 3109 4503 3112 4507
rect 3126 4492 3129 4508
rect 3134 4452 3137 4458
rect 3114 4448 3118 4451
rect 3078 4282 3081 4338
rect 3086 4291 3089 4348
rect 3126 4342 3129 4408
rect 3134 4372 3137 4418
rect 3142 4362 3145 4538
rect 3154 4478 3158 4481
rect 3174 4442 3177 4548
rect 3182 4512 3185 4518
rect 3190 4462 3193 4638
rect 3198 4632 3201 4658
rect 3238 4592 3241 4668
rect 3234 4548 3238 4551
rect 3262 4542 3265 4658
rect 3278 4562 3281 4648
rect 3294 4542 3297 4638
rect 3302 4562 3305 4728
rect 3318 4632 3321 4658
rect 3262 4482 3265 4538
rect 3202 4468 3206 4471
rect 3250 4468 3254 4471
rect 3278 4462 3281 4468
rect 3234 4458 3238 4461
rect 3258 4458 3262 4461
rect 3174 4402 3177 4418
rect 3190 4402 3193 4458
rect 3214 4452 3217 4458
rect 3242 4448 3246 4451
rect 3214 4422 3217 4448
rect 3150 4362 3153 4368
rect 3174 4361 3177 4398
rect 3190 4362 3193 4368
rect 3174 4358 3185 4361
rect 3134 4352 3137 4358
rect 3146 4348 3150 4351
rect 3170 4348 3174 4351
rect 3162 4338 3166 4341
rect 3096 4303 3098 4307
rect 3102 4303 3105 4307
rect 3109 4303 3112 4307
rect 3086 4288 3094 4291
rect 3086 4192 3089 4268
rect 3102 4252 3105 4268
rect 3118 4252 3121 4318
rect 3142 4262 3145 4338
rect 3150 4272 3153 4278
rect 3158 4262 3161 4268
rect 3182 4262 3185 4358
rect 3194 4338 3198 4341
rect 3194 4318 3198 4321
rect 3238 4262 3241 4278
rect 3246 4272 3249 4338
rect 3146 4258 3150 4261
rect 3194 4258 3198 4261
rect 3166 4251 3169 4258
rect 3146 4248 3169 4251
rect 3074 4148 3078 4151
rect 3082 4138 3086 4141
rect 3022 4122 3025 4138
rect 3102 4132 3105 4248
rect 3174 4172 3177 4218
rect 3246 4172 3249 4268
rect 3254 4212 3257 4458
rect 3286 4451 3289 4518
rect 3294 4492 3297 4538
rect 3282 4448 3289 4451
rect 3262 4382 3265 4418
rect 3302 4372 3305 4518
rect 3310 4362 3313 4618
rect 3318 4552 3321 4628
rect 3334 4552 3337 4698
rect 3350 4632 3353 4858
rect 3366 4832 3369 4848
rect 3374 4822 3377 4858
rect 3382 4842 3385 4868
rect 3398 4862 3401 4868
rect 3558 4862 3561 4878
rect 3482 4858 3486 4861
rect 3406 4842 3409 4858
rect 3582 4832 3585 4858
rect 3430 4792 3433 4818
rect 3402 4788 3406 4791
rect 3414 4762 3417 4778
rect 3430 4772 3433 4778
rect 3446 4762 3449 4798
rect 3462 4792 3465 4828
rect 3608 4803 3610 4807
rect 3614 4803 3617 4807
rect 3621 4803 3624 4807
rect 3670 4782 3673 4858
rect 3694 4832 3697 4858
rect 3730 4818 3734 4821
rect 3766 4812 3769 4858
rect 3782 4832 3785 4858
rect 3790 4842 3793 4858
rect 3582 4762 3585 4768
rect 3418 4758 3425 4761
rect 3450 4758 3457 4761
rect 3366 4732 3369 4738
rect 3382 4702 3385 4758
rect 3402 4748 3406 4751
rect 3410 4738 3414 4741
rect 3422 4741 3425 4758
rect 3434 4748 3438 4751
rect 3422 4738 3433 4741
rect 3442 4738 3446 4741
rect 3430 4682 3433 4738
rect 3366 4672 3369 4678
rect 3378 4668 3382 4671
rect 3398 4662 3401 4668
rect 3406 4662 3409 4668
rect 3370 4658 3374 4661
rect 3350 4562 3353 4568
rect 3354 4548 3358 4551
rect 3334 4542 3337 4548
rect 3318 4532 3321 4538
rect 3334 4462 3337 4478
rect 3366 4472 3369 4658
rect 3406 4572 3409 4658
rect 3406 4551 3409 4558
rect 3374 4522 3377 4528
rect 3390 4521 3393 4538
rect 3382 4518 3393 4521
rect 3382 4472 3385 4518
rect 3398 4482 3401 4508
rect 3414 4472 3417 4678
rect 3422 4672 3425 4678
rect 3438 4542 3441 4618
rect 3454 4502 3457 4758
rect 3510 4752 3513 4758
rect 3466 4748 3470 4751
rect 3470 4692 3473 4738
rect 3486 4732 3489 4738
rect 3574 4732 3577 4738
rect 3486 4672 3489 4728
rect 3562 4718 3566 4721
rect 3534 4682 3537 4688
rect 3550 4682 3553 4718
rect 3574 4682 3577 4688
rect 3582 4672 3585 4748
rect 3606 4662 3609 4748
rect 3622 4722 3625 4758
rect 3790 4752 3793 4838
rect 3806 4772 3809 4788
rect 3822 4772 3825 4818
rect 3830 4792 3833 4878
rect 3862 4872 3865 4878
rect 3874 4868 3878 4871
rect 3870 4862 3873 4868
rect 3850 4858 3854 4861
rect 3878 4852 3881 4858
rect 3910 4832 3913 4868
rect 3918 4842 3921 4858
rect 4046 4852 4049 4859
rect 4062 4832 4065 4868
rect 4206 4862 4209 4868
rect 4210 4858 4214 4861
rect 4142 4842 4145 4858
rect 4166 4832 4169 4858
rect 3910 4772 3913 4828
rect 3974 4802 3977 4818
rect 3894 4762 3897 4768
rect 3850 4758 3854 4761
rect 3770 4748 3774 4751
rect 3638 4712 3641 4748
rect 3710 4742 3713 4748
rect 3790 4742 3793 4748
rect 3770 4738 3774 4741
rect 3646 4682 3649 4738
rect 3614 4672 3617 4678
rect 3470 4652 3473 4659
rect 3554 4658 3558 4661
rect 3646 4652 3649 4658
rect 3586 4648 3590 4651
rect 3490 4548 3494 4551
rect 3474 4538 3478 4541
rect 3466 4518 3470 4521
rect 3486 4472 3489 4478
rect 3358 4452 3361 4458
rect 3406 4392 3409 4418
rect 3346 4358 3350 4361
rect 3270 4352 3273 4358
rect 3134 4142 3137 4148
rect 2934 4052 2937 4058
rect 2950 4052 2953 4068
rect 2958 4062 2961 4068
rect 2990 4062 2993 4098
rect 3014 4062 3017 4068
rect 3022 4062 3025 4078
rect 3030 4062 3033 4108
rect 3054 4092 3057 4118
rect 3070 4112 3073 4128
rect 3046 4062 3049 4078
rect 3070 4072 3073 4108
rect 3086 4092 3089 4118
rect 3096 4103 3098 4107
rect 3102 4103 3105 4107
rect 3109 4103 3112 4107
rect 3058 4068 3062 4071
rect 3078 4062 3081 4088
rect 2974 4012 2977 4048
rect 2994 4018 2998 4021
rect 2978 3988 2982 3991
rect 2870 3962 2873 3968
rect 2882 3958 2886 3961
rect 2806 3932 2809 3938
rect 2854 3932 2857 3938
rect 2790 3882 2793 3908
rect 2806 3862 2809 3928
rect 2838 3891 2841 3918
rect 2830 3888 2841 3891
rect 2814 3862 2817 3888
rect 2726 3852 2729 3858
rect 2738 3848 2742 3851
rect 2662 3792 2665 3818
rect 2674 3758 2678 3761
rect 2646 3732 2649 3738
rect 2654 3692 2657 3748
rect 2694 3732 2697 3748
rect 2702 3742 2705 3828
rect 2710 3752 2713 3818
rect 2742 3752 2745 3838
rect 2750 3832 2753 3858
rect 2766 3842 2769 3848
rect 2782 3782 2785 3848
rect 2618 3668 2622 3671
rect 2658 3668 2662 3671
rect 2610 3658 2614 3661
rect 2714 3658 2718 3661
rect 2646 3652 2649 3658
rect 2682 3648 2686 3651
rect 2550 3532 2553 3638
rect 2534 3482 2537 3488
rect 2526 3462 2529 3468
rect 2518 3362 2521 3368
rect 2526 3352 2529 3458
rect 2550 3452 2553 3518
rect 2558 3492 2561 3608
rect 2584 3603 2586 3607
rect 2590 3603 2593 3607
rect 2597 3603 2600 3607
rect 2566 3532 2569 3547
rect 2582 3542 2585 3568
rect 2598 3492 2601 3588
rect 2614 3552 2617 3608
rect 2694 3562 2697 3578
rect 2622 3542 2625 3548
rect 2662 3542 2665 3548
rect 2642 3538 2646 3541
rect 2642 3528 2646 3531
rect 2630 3522 2633 3528
rect 2654 3522 2657 3528
rect 2622 3472 2625 3488
rect 2630 3472 2633 3488
rect 2542 3372 2545 3418
rect 2550 3402 2553 3448
rect 2566 3442 2569 3468
rect 2630 3462 2633 3468
rect 2614 3452 2617 3458
rect 2646 3452 2649 3458
rect 2584 3403 2586 3407
rect 2590 3403 2593 3407
rect 2597 3403 2600 3407
rect 2534 3362 2537 3368
rect 2550 3352 2553 3358
rect 2534 3341 2537 3348
rect 2530 3338 2537 3341
rect 2558 3342 2561 3368
rect 2522 3328 2526 3331
rect 2534 3232 2537 3338
rect 2566 3332 2569 3348
rect 2606 3342 2609 3388
rect 2614 3372 2617 3448
rect 2630 3442 2633 3448
rect 2654 3442 2657 3448
rect 2618 3358 2622 3361
rect 2550 3272 2553 3288
rect 2542 3242 2545 3248
rect 2558 3192 2561 3258
rect 2518 3152 2521 3168
rect 2566 3152 2569 3288
rect 2582 3282 2585 3318
rect 2638 3278 2654 3281
rect 2574 3262 2577 3268
rect 2614 3262 2617 3268
rect 2630 3262 2633 3268
rect 2594 3248 2598 3251
rect 2626 3248 2630 3251
rect 2584 3203 2586 3207
rect 2590 3203 2593 3207
rect 2597 3203 2600 3207
rect 2638 3172 2641 3278
rect 2650 3268 2654 3271
rect 2650 3258 2654 3261
rect 2610 3168 2614 3171
rect 2642 3168 2646 3171
rect 2538 3148 2542 3151
rect 2518 3072 2521 3118
rect 2526 3082 2529 3148
rect 2566 3142 2569 3148
rect 2538 3138 2542 3141
rect 2542 3081 2545 3138
rect 2550 3132 2553 3138
rect 2558 3092 2561 3128
rect 2574 3092 2577 3148
rect 2606 3142 2609 3148
rect 2630 3142 2633 3148
rect 2638 3122 2641 3138
rect 2614 3082 2617 3088
rect 2542 3078 2553 3081
rect 2510 3062 2513 3068
rect 2550 3062 2553 3078
rect 2566 3072 2569 3078
rect 2578 3068 2582 3071
rect 2490 3058 2494 3061
rect 2430 3042 2433 3048
rect 2410 3038 2414 3041
rect 2422 3002 2425 3018
rect 2382 2952 2385 2958
rect 2406 2952 2409 2998
rect 2342 2932 2345 2938
rect 2382 2882 2385 2938
rect 2422 2872 2425 2978
rect 2462 2952 2465 3008
rect 2494 2982 2497 3048
rect 2506 3038 2510 3041
rect 2526 3032 2529 3058
rect 2470 2962 2473 2968
rect 2486 2962 2489 2968
rect 2494 2952 2497 2958
rect 2490 2948 2494 2951
rect 2522 2948 2526 2951
rect 2446 2942 2449 2948
rect 2502 2922 2505 2948
rect 2518 2912 2521 2918
rect 2486 2872 2489 2898
rect 2414 2862 2417 2868
rect 2422 2862 2425 2868
rect 2350 2782 2353 2858
rect 2382 2852 2385 2859
rect 2446 2852 2449 2868
rect 2462 2852 2465 2868
rect 2470 2852 2473 2868
rect 2510 2862 2513 2868
rect 2426 2848 2430 2851
rect 2302 2672 2305 2778
rect 2446 2772 2449 2848
rect 2470 2822 2473 2848
rect 2486 2762 2489 2858
rect 2518 2842 2521 2868
rect 2534 2862 2537 3058
rect 2542 3052 2545 3058
rect 2550 3032 2553 3058
rect 2542 2962 2545 2968
rect 2558 2962 2561 3068
rect 2654 3062 2657 3128
rect 2662 3102 2665 3538
rect 2670 3532 2673 3538
rect 2678 3502 2681 3548
rect 2694 3542 2697 3548
rect 2702 3542 2705 3618
rect 2726 3602 2729 3718
rect 2750 3682 2753 3748
rect 2762 3738 2766 3741
rect 2782 3672 2785 3728
rect 2790 3682 2793 3818
rect 2806 3702 2809 3858
rect 2830 3852 2833 3888
rect 2842 3878 2846 3881
rect 2814 3692 2817 3818
rect 2838 3792 2841 3808
rect 2822 3742 2825 3748
rect 2822 3702 2825 3738
rect 2790 3672 2793 3678
rect 2830 3671 2833 3788
rect 2854 3762 2857 3928
rect 2862 3922 2865 3938
rect 2854 3742 2857 3748
rect 2862 3742 2865 3748
rect 2870 3722 2873 3948
rect 2902 3942 2905 3978
rect 2918 3951 2921 3968
rect 2982 3892 2985 3898
rect 2950 3872 2953 3878
rect 2962 3868 2966 3871
rect 2918 3863 2921 3868
rect 2878 3752 2881 3778
rect 2934 3772 2937 3868
rect 2954 3858 2958 3861
rect 2974 3852 2977 3868
rect 2990 3862 2993 3958
rect 3014 3942 3017 4048
rect 3094 4042 3097 4058
rect 3118 4012 3121 4128
rect 3062 3972 3065 4008
rect 3074 3958 3081 3961
rect 3038 3952 3041 3958
rect 3066 3948 3070 3951
rect 2998 3872 3001 3918
rect 3006 3872 3009 3918
rect 3014 3912 3017 3938
rect 3046 3932 3049 3938
rect 3014 3872 3017 3878
rect 3002 3858 3006 3861
rect 2986 3848 2990 3851
rect 3014 3772 3017 3858
rect 3022 3832 3025 3918
rect 3042 3868 3046 3871
rect 3054 3852 3057 3918
rect 3078 3892 3081 3958
rect 3066 3868 3070 3871
rect 3086 3852 3089 3948
rect 3094 3922 3097 3938
rect 3134 3922 3137 4138
rect 3142 4112 3145 4118
rect 3182 4072 3185 4118
rect 3198 4082 3201 4108
rect 3206 4102 3209 4147
rect 3222 4142 3225 4168
rect 3250 4148 3254 4151
rect 3242 4138 3246 4141
rect 3270 4132 3273 4138
rect 3210 4088 3214 4091
rect 3246 4072 3249 4078
rect 3158 4062 3161 4068
rect 3182 4062 3185 4068
rect 3214 4012 3217 4018
rect 3186 3948 3190 3951
rect 3250 3948 3254 3951
rect 3096 3903 3098 3907
rect 3102 3903 3105 3907
rect 3109 3903 3112 3907
rect 3142 3862 3145 3898
rect 3166 3872 3169 3948
rect 3230 3921 3233 3928
rect 3254 3922 3257 3938
rect 3222 3918 3233 3921
rect 3222 3882 3225 3918
rect 3238 3902 3241 3918
rect 3254 3872 3257 3918
rect 3262 3871 3265 4118
rect 3278 4082 3281 4358
rect 3294 4342 3297 4348
rect 3310 4292 3313 4338
rect 3366 4332 3369 4338
rect 3314 4278 3318 4281
rect 3306 4268 3310 4271
rect 3326 4252 3329 4318
rect 3334 4262 3337 4298
rect 3374 4272 3377 4388
rect 3442 4368 3446 4371
rect 3434 4358 3438 4361
rect 3446 4352 3449 4358
rect 3398 4342 3401 4347
rect 3414 4342 3417 4348
rect 3454 4342 3457 4458
rect 3462 4362 3465 4368
rect 3470 4352 3473 4418
rect 3494 4382 3497 4538
rect 3502 4492 3505 4558
rect 3510 4552 3513 4558
rect 3518 4552 3521 4638
rect 3534 4562 3537 4618
rect 3530 4538 3534 4541
rect 3502 4452 3505 4458
rect 3510 4452 3513 4518
rect 3534 4512 3537 4518
rect 3542 4512 3545 4618
rect 3550 4562 3553 4648
rect 3610 4618 3614 4621
rect 3608 4603 3610 4607
rect 3614 4603 3617 4607
rect 3621 4603 3624 4607
rect 3646 4562 3649 4618
rect 3566 4552 3569 4558
rect 3594 4547 3598 4550
rect 3634 4548 3638 4551
rect 3654 4551 3657 4718
rect 3734 4672 3737 4738
rect 3750 4722 3753 4728
rect 3798 4672 3801 4748
rect 3806 4682 3809 4758
rect 3866 4748 3870 4751
rect 3838 4742 3841 4748
rect 3690 4668 3694 4671
rect 3726 4663 3729 4668
rect 3674 4658 3678 4661
rect 3662 4642 3665 4648
rect 3646 4548 3657 4551
rect 3670 4551 3673 4648
rect 3686 4592 3689 4658
rect 3666 4548 3673 4551
rect 3534 4472 3537 4488
rect 3606 4482 3609 4498
rect 3594 4468 3598 4471
rect 3542 4462 3545 4468
rect 3534 4442 3537 4458
rect 3542 4432 3545 4458
rect 3526 4402 3529 4418
rect 3550 4392 3553 4458
rect 3566 4452 3569 4458
rect 3598 4452 3601 4458
rect 3562 4448 3566 4451
rect 3590 4442 3593 4448
rect 3550 4362 3553 4388
rect 3546 4348 3550 4351
rect 3462 4342 3465 4348
rect 3478 4342 3481 4348
rect 3502 4342 3505 4348
rect 3414 4272 3417 4338
rect 3454 4282 3457 4338
rect 3486 4332 3489 4338
rect 3346 4268 3350 4271
rect 3346 4258 3350 4261
rect 3346 4248 3350 4251
rect 3286 4172 3289 4188
rect 3302 4142 3305 4168
rect 3318 4092 3321 4248
rect 3366 4242 3369 4258
rect 3398 4152 3401 4158
rect 3406 4152 3409 4259
rect 3422 4182 3425 4278
rect 3474 4268 3478 4271
rect 3482 4258 3486 4261
rect 3502 4252 3505 4318
rect 3510 4282 3513 4288
rect 3510 4262 3513 4268
rect 3526 4252 3529 4348
rect 3598 4342 3601 4448
rect 3608 4403 3610 4407
rect 3614 4403 3617 4407
rect 3621 4403 3624 4407
rect 3622 4372 3625 4378
rect 3630 4351 3633 4418
rect 3646 4372 3649 4548
rect 3662 4542 3665 4548
rect 3686 4542 3689 4558
rect 3714 4548 3718 4551
rect 3670 4532 3673 4538
rect 3662 4442 3665 4459
rect 3622 4348 3633 4351
rect 3670 4352 3673 4468
rect 3726 4462 3729 4488
rect 3734 4472 3737 4588
rect 3750 4572 3753 4658
rect 3798 4652 3801 4668
rect 3814 4642 3817 4718
rect 3822 4702 3825 4738
rect 3830 4702 3833 4738
rect 3838 4712 3841 4738
rect 3878 4722 3881 4748
rect 3886 4732 3889 4738
rect 3830 4682 3833 4698
rect 3878 4682 3881 4688
rect 3910 4682 3913 4768
rect 3946 4748 3950 4751
rect 3974 4742 3977 4758
rect 3878 4652 3881 4659
rect 3782 4621 3785 4638
rect 3782 4618 3790 4621
rect 3810 4618 3814 4621
rect 3758 4492 3761 4548
rect 3766 4512 3769 4518
rect 3782 4492 3785 4618
rect 3766 4482 3769 4488
rect 3678 4392 3681 4438
rect 3582 4282 3585 4318
rect 3590 4312 3593 4338
rect 3598 4272 3601 4318
rect 3606 4272 3609 4288
rect 3622 4272 3625 4348
rect 3534 4262 3537 4268
rect 3558 4262 3561 4268
rect 3574 4262 3577 4268
rect 3566 4252 3569 4258
rect 3582 4251 3585 4268
rect 3630 4262 3633 4338
rect 3642 4318 3646 4321
rect 3654 4262 3657 4338
rect 3594 4258 3598 4261
rect 3578 4248 3585 4251
rect 3630 4252 3633 4258
rect 3466 4218 3470 4221
rect 3414 4162 3417 4168
rect 3326 4142 3329 4148
rect 3422 4142 3425 4178
rect 3434 4168 3438 4171
rect 3446 4162 3449 4218
rect 3478 4192 3481 4248
rect 3434 4148 3438 4151
rect 3426 4138 3433 4141
rect 3390 4132 3393 4138
rect 3382 4101 3385 4118
rect 3390 4112 3393 4128
rect 3382 4098 3393 4101
rect 3358 4092 3361 4098
rect 3334 4072 3337 4088
rect 3390 4082 3393 4098
rect 3430 4092 3433 4138
rect 3446 4122 3449 4158
rect 3458 4148 3465 4151
rect 3462 4142 3465 4148
rect 3454 4092 3457 4138
rect 3402 4088 3406 4091
rect 3446 4082 3449 4088
rect 3390 4072 3393 4078
rect 3462 4072 3465 4138
rect 3470 4132 3473 4148
rect 3490 4138 3494 4141
rect 3458 4068 3462 4071
rect 3274 4058 3278 4061
rect 3310 4052 3313 4068
rect 3330 4048 3334 4051
rect 3342 4012 3345 4058
rect 3366 4012 3369 4048
rect 3270 3952 3273 3958
rect 3270 3882 3273 3948
rect 3262 3868 3270 3871
rect 3222 3862 3225 3868
rect 3246 3862 3249 3868
rect 3286 3862 3289 3998
rect 3374 3972 3377 4068
rect 3382 4062 3385 4068
rect 3406 4062 3409 4068
rect 3470 4062 3473 4108
rect 3390 3992 3393 4048
rect 3414 4022 3417 4058
rect 3470 4052 3473 4058
rect 3478 4052 3481 4118
rect 3502 4072 3505 4148
rect 3490 4068 3494 4071
rect 3342 3951 3345 3958
rect 3390 3952 3393 3988
rect 3406 3962 3409 3968
rect 3430 3962 3433 3988
rect 3510 3972 3513 4148
rect 3518 4071 3521 4218
rect 3526 4192 3529 4228
rect 3534 4072 3537 4098
rect 3518 4068 3526 4071
rect 3542 4062 3545 4138
rect 3550 4072 3553 4218
rect 3558 4172 3561 4218
rect 3566 4152 3569 4158
rect 3582 4142 3585 4208
rect 3608 4203 3610 4207
rect 3614 4203 3617 4207
rect 3621 4203 3624 4207
rect 3590 4122 3593 4148
rect 3606 4132 3609 4138
rect 3630 4122 3633 4208
rect 3638 4182 3641 4258
rect 3662 4252 3665 4318
rect 3650 4248 3654 4251
rect 3650 4218 3654 4221
rect 3642 4168 3646 4171
rect 3686 4141 3689 4388
rect 3718 4282 3721 4338
rect 3694 4152 3697 4158
rect 3702 4142 3705 4268
rect 3718 4263 3721 4268
rect 3734 4142 3737 4468
rect 3782 4462 3785 4468
rect 3742 4452 3745 4458
rect 3758 4452 3761 4458
rect 3790 4451 3793 4508
rect 3798 4472 3801 4618
rect 3870 4602 3873 4628
rect 3810 4548 3814 4551
rect 3786 4448 3793 4451
rect 3742 4351 3745 4398
rect 3758 4342 3761 4378
rect 3774 4352 3777 4418
rect 3790 4372 3793 4448
rect 3798 4372 3801 4458
rect 3806 4432 3809 4468
rect 3778 4338 3782 4341
rect 3790 4282 3793 4318
rect 3782 4272 3785 4278
rect 3754 4268 3758 4271
rect 3750 4252 3753 4258
rect 3766 4252 3769 4258
rect 3774 4202 3777 4268
rect 3790 4242 3793 4258
rect 3790 4182 3793 4218
rect 3786 4168 3790 4171
rect 3746 4158 3750 4161
rect 3742 4142 3745 4148
rect 3758 4142 3761 4158
rect 3766 4142 3769 4148
rect 3782 4142 3785 4148
rect 3686 4138 3697 4141
rect 3518 4042 3521 4058
rect 3558 4052 3561 4118
rect 3574 4092 3577 4118
rect 3566 4072 3569 4088
rect 3638 4072 3641 4098
rect 3662 4092 3665 4108
rect 3694 4092 3697 4138
rect 3734 4112 3737 4138
rect 3730 4068 3734 4071
rect 3574 4062 3577 4068
rect 3650 4058 3654 4061
rect 3674 4058 3678 4061
rect 3518 4022 3521 4028
rect 3542 4002 3545 4018
rect 3486 3952 3489 3958
rect 3070 3842 3073 3848
rect 3086 3832 3089 3848
rect 3022 3772 3025 3818
rect 2894 3752 2897 3758
rect 2910 3752 2913 3758
rect 2918 3752 2921 3768
rect 2878 3732 2881 3748
rect 2974 3742 2977 3748
rect 2998 3742 3001 3748
rect 3110 3742 3113 3748
rect 2898 3738 2902 3741
rect 3082 3738 3086 3741
rect 2826 3668 2833 3671
rect 2894 3672 2897 3698
rect 2998 3672 3001 3738
rect 3014 3702 3017 3738
rect 3096 3703 3098 3707
rect 3102 3703 3105 3707
rect 3109 3703 3112 3707
rect 3098 3688 3102 3691
rect 2906 3668 2910 3671
rect 2954 3668 2958 3671
rect 3090 3668 3094 3671
rect 2710 3582 2713 3588
rect 2726 3572 2729 3578
rect 2734 3572 2737 3668
rect 2782 3662 2785 3668
rect 2794 3658 2798 3661
rect 2942 3658 2950 3661
rect 2994 3659 2998 3662
rect 3066 3658 3070 3661
rect 2770 3648 2774 3651
rect 2786 3648 2798 3651
rect 2790 3552 2793 3568
rect 2710 3522 2713 3548
rect 2762 3547 2766 3550
rect 2710 3492 2713 3518
rect 2790 3482 2793 3548
rect 2814 3492 2817 3658
rect 2826 3578 2830 3581
rect 2838 3572 2841 3618
rect 2886 3572 2889 3578
rect 2858 3558 2870 3561
rect 2858 3548 2862 3551
rect 2830 3532 2833 3538
rect 2726 3472 2729 3478
rect 2790 3472 2793 3478
rect 2674 3468 2678 3471
rect 2674 3458 2678 3461
rect 2822 3462 2825 3498
rect 2710 3442 2713 3459
rect 2774 3442 2777 3448
rect 2670 3432 2673 3438
rect 2758 3352 2761 3358
rect 2682 3348 2686 3351
rect 2670 3242 2673 3348
rect 2678 3262 2681 3298
rect 2774 3292 2777 3438
rect 2750 3282 2753 3288
rect 2734 3262 2737 3268
rect 2782 3262 2785 3428
rect 2838 3422 2841 3548
rect 2862 3512 2865 3538
rect 2870 3522 2873 3548
rect 2886 3472 2889 3538
rect 2894 3492 2897 3498
rect 2874 3458 2878 3461
rect 2886 3452 2889 3468
rect 2874 3418 2878 3421
rect 2818 3368 2822 3371
rect 2854 3362 2857 3368
rect 2834 3358 2838 3361
rect 2858 3358 2862 3361
rect 2870 3352 2873 3408
rect 2886 3352 2889 3358
rect 2834 3348 2841 3351
rect 2818 3338 2822 3341
rect 2798 3272 2801 3318
rect 2822 3292 2825 3308
rect 2770 3258 2774 3261
rect 2802 3258 2806 3261
rect 2694 3252 2697 3258
rect 2742 3252 2745 3258
rect 2770 3248 2777 3251
rect 2754 3238 2758 3241
rect 2718 3202 2721 3218
rect 2750 3192 2753 3218
rect 2782 3212 2785 3258
rect 2826 3248 2830 3251
rect 2774 3192 2777 3198
rect 2698 3148 2702 3151
rect 2726 3142 2729 3188
rect 2806 3172 2809 3178
rect 2822 3172 2825 3178
rect 2838 3172 2841 3348
rect 2878 3332 2881 3338
rect 2846 3262 2849 3268
rect 2862 3262 2865 3298
rect 2886 3262 2889 3268
rect 2894 3262 2897 3468
rect 2902 3412 2905 3658
rect 2930 3648 2934 3651
rect 2922 3547 2926 3550
rect 2934 3542 2937 3568
rect 2942 3532 2945 3658
rect 2958 3651 2961 3658
rect 2954 3648 2961 3651
rect 3042 3648 3046 3651
rect 2978 3578 2982 3581
rect 2942 3482 2945 3518
rect 2974 3482 2977 3568
rect 2990 3532 2993 3588
rect 3006 3562 3009 3578
rect 3038 3552 3041 3588
rect 3054 3552 3057 3558
rect 3062 3552 3065 3638
rect 3078 3632 3081 3658
rect 3026 3548 3030 3551
rect 3090 3548 3094 3551
rect 3006 3542 3009 3548
rect 3034 3538 3038 3541
rect 3050 3538 3054 3541
rect 3022 3512 3025 3538
rect 2910 3422 2913 3478
rect 3046 3472 3049 3478
rect 3054 3462 3057 3468
rect 2986 3458 2990 3461
rect 2926 3452 2929 3458
rect 2926 3372 2929 3448
rect 3042 3438 3046 3441
rect 2934 3361 2937 3418
rect 2942 3372 2945 3418
rect 3054 3412 3057 3458
rect 2934 3358 2945 3361
rect 2930 3348 2934 3351
rect 2942 3342 2945 3358
rect 2958 3342 2961 3378
rect 2906 3338 2910 3341
rect 2910 3292 2913 3318
rect 2902 3262 2905 3268
rect 2934 3262 2937 3268
rect 2894 3252 2897 3258
rect 2910 3252 2913 3258
rect 2790 3162 2793 3168
rect 2574 3052 2577 3058
rect 2594 3048 2598 3051
rect 2614 3012 2617 3018
rect 2584 3003 2586 3007
rect 2590 3003 2593 3007
rect 2597 3003 2600 3007
rect 2574 2972 2577 2998
rect 2678 2971 2681 3128
rect 2742 3112 2745 3148
rect 2766 3142 2769 3158
rect 2854 3151 2857 3198
rect 2758 3132 2761 3138
rect 2774 3102 2777 3148
rect 2798 3142 2801 3148
rect 2806 3142 2809 3148
rect 2798 3122 2801 3138
rect 2710 3082 2713 3088
rect 2694 3062 2697 3068
rect 2710 3052 2713 3078
rect 2670 2968 2681 2971
rect 2702 2968 2710 2971
rect 2630 2962 2633 2968
rect 2670 2952 2673 2968
rect 2686 2962 2689 2968
rect 2702 2952 2705 2968
rect 2618 2948 2622 2951
rect 2558 2942 2561 2948
rect 2586 2938 2590 2941
rect 2542 2932 2545 2938
rect 2558 2862 2561 2868
rect 2502 2792 2505 2838
rect 2526 2812 2529 2858
rect 2522 2788 2526 2791
rect 2358 2752 2361 2758
rect 2430 2752 2433 2758
rect 2534 2752 2537 2758
rect 2542 2752 2545 2818
rect 2574 2761 2577 2918
rect 2598 2862 2601 2898
rect 2606 2842 2609 2938
rect 2584 2803 2586 2807
rect 2590 2803 2593 2807
rect 2597 2803 2600 2807
rect 2606 2772 2609 2818
rect 2574 2758 2582 2761
rect 2386 2748 2390 2751
rect 2562 2748 2566 2751
rect 2310 2742 2313 2748
rect 2334 2742 2337 2748
rect 2298 2668 2302 2671
rect 2222 2662 2225 2668
rect 2270 2662 2273 2668
rect 2154 2658 2158 2661
rect 2258 2648 2262 2651
rect 2298 2648 2302 2651
rect 2098 2548 2102 2551
rect 2138 2548 2142 2551
rect 2150 2541 2153 2558
rect 2158 2552 2161 2568
rect 2142 2538 2153 2541
rect 2072 2503 2074 2507
rect 2078 2503 2081 2507
rect 2085 2503 2088 2507
rect 2094 2482 2097 2538
rect 2102 2512 2105 2538
rect 2110 2522 2113 2528
rect 2118 2492 2121 2538
rect 2134 2532 2137 2538
rect 2142 2492 2145 2538
rect 2058 2478 2062 2481
rect 2158 2472 2161 2518
rect 2166 2472 2169 2508
rect 2198 2472 2201 2508
rect 2206 2502 2209 2638
rect 2246 2632 2249 2638
rect 2214 2532 2217 2548
rect 2214 2492 2217 2518
rect 2222 2492 2225 2528
rect 2238 2522 2241 2578
rect 2270 2562 2273 2598
rect 2294 2552 2297 2598
rect 2302 2551 2305 2588
rect 2334 2562 2337 2728
rect 2350 2722 2353 2748
rect 2386 2738 2390 2741
rect 2366 2702 2369 2718
rect 2430 2702 2433 2728
rect 2362 2668 2366 2671
rect 2374 2662 2377 2668
rect 2382 2662 2385 2668
rect 2414 2662 2417 2668
rect 2422 2662 2425 2698
rect 2430 2672 2433 2698
rect 2446 2672 2449 2748
rect 2478 2702 2481 2738
rect 2542 2702 2545 2728
rect 2526 2692 2529 2698
rect 2462 2663 2465 2668
rect 2350 2592 2353 2658
rect 2402 2648 2406 2651
rect 2314 2558 2318 2561
rect 2366 2552 2369 2588
rect 2302 2548 2313 2551
rect 2258 2538 2262 2541
rect 2238 2492 2241 2498
rect 2246 2472 2249 2478
rect 2030 2352 2033 2448
rect 2046 2362 2049 2468
rect 2070 2452 2073 2468
rect 2118 2462 2121 2468
rect 2126 2462 2129 2468
rect 2166 2462 2169 2468
rect 2070 2442 2073 2448
rect 2018 2348 2022 2351
rect 2002 2338 2006 2341
rect 1978 2328 1982 2331
rect 2022 2322 2025 2338
rect 2006 2312 2009 2318
rect 1990 2272 1993 2308
rect 1998 2282 2001 2288
rect 2014 2272 2017 2278
rect 1934 2268 1942 2271
rect 1942 2262 1945 2268
rect 1998 2262 2001 2268
rect 1870 2222 1873 2258
rect 1910 2212 1913 2258
rect 1966 2222 1969 2258
rect 1930 2218 1934 2221
rect 1862 2151 1865 2158
rect 1814 2072 1817 2128
rect 1846 2102 1849 2138
rect 1870 2062 1873 2088
rect 1878 2081 1881 2198
rect 1902 2162 1905 2168
rect 1926 2162 1929 2198
rect 1934 2192 1937 2208
rect 1886 2092 1889 2118
rect 1894 2112 1897 2138
rect 1902 2102 1905 2148
rect 1918 2142 1921 2158
rect 1950 2152 1953 2198
rect 1958 2182 1961 2218
rect 1926 2112 1929 2148
rect 1958 2142 1961 2158
rect 1974 2152 1977 2248
rect 1990 2172 1993 2188
rect 1990 2162 1993 2168
rect 1986 2148 1990 2151
rect 1998 2142 2001 2258
rect 2014 2252 2017 2258
rect 2006 2142 2009 2218
rect 2014 2182 2017 2218
rect 1970 2138 1974 2141
rect 1878 2078 1889 2081
rect 1826 2058 1830 2061
rect 1758 2002 1761 2018
rect 1774 1982 1777 2028
rect 1782 2002 1785 2058
rect 1838 2052 1841 2058
rect 1850 2048 1854 2051
rect 1790 1992 1793 2008
rect 1734 1952 1737 1958
rect 1718 1892 1721 1938
rect 1726 1862 1729 1948
rect 1738 1868 1742 1871
rect 1750 1862 1753 1958
rect 1774 1952 1777 1978
rect 1782 1942 1785 1948
rect 1762 1938 1766 1941
rect 1766 1872 1769 1908
rect 1806 1872 1809 2028
rect 1862 2022 1865 2058
rect 1826 1958 1833 1961
rect 1866 1958 1870 1961
rect 1830 1892 1833 1958
rect 1818 1868 1822 1871
rect 1730 1858 1734 1861
rect 1770 1858 1774 1861
rect 1810 1858 1814 1861
rect 1750 1852 1753 1858
rect 1782 1852 1785 1858
rect 1710 1781 1713 1818
rect 1710 1778 1718 1781
rect 1726 1752 1729 1778
rect 1750 1762 1753 1848
rect 1718 1742 1721 1748
rect 1726 1722 1729 1748
rect 1734 1742 1737 1748
rect 1742 1722 1745 1758
rect 1750 1742 1753 1748
rect 1674 1658 1678 1661
rect 1702 1652 1705 1668
rect 1726 1662 1729 1668
rect 1742 1662 1745 1698
rect 1758 1662 1761 1788
rect 1770 1758 1774 1761
rect 1790 1752 1793 1758
rect 1778 1748 1782 1751
rect 1770 1658 1774 1661
rect 1694 1632 1697 1648
rect 1718 1632 1721 1658
rect 1750 1652 1753 1658
rect 1726 1648 1734 1651
rect 1670 1552 1673 1558
rect 1678 1552 1681 1558
rect 1694 1552 1697 1598
rect 1726 1592 1729 1648
rect 1758 1602 1761 1648
rect 1790 1632 1793 1748
rect 1798 1712 1801 1738
rect 1806 1672 1809 1728
rect 1830 1692 1833 1868
rect 1838 1862 1841 1948
rect 1858 1938 1862 1941
rect 1846 1932 1849 1938
rect 1878 1912 1881 2058
rect 1862 1872 1865 1908
rect 1846 1851 1849 1868
rect 1854 1862 1857 1868
rect 1846 1848 1857 1851
rect 1838 1842 1841 1848
rect 1822 1662 1825 1688
rect 1810 1658 1814 1661
rect 1774 1592 1777 1598
rect 1702 1552 1705 1558
rect 1790 1552 1793 1578
rect 1798 1562 1801 1658
rect 1830 1552 1833 1588
rect 1846 1581 1849 1658
rect 1854 1592 1857 1848
rect 1870 1762 1873 1848
rect 1886 1802 1889 2078
rect 1926 2072 1929 2078
rect 1934 2072 1937 2138
rect 1942 2132 1945 2138
rect 1962 2128 1966 2131
rect 1990 2112 1993 2118
rect 2014 2092 2017 2128
rect 2022 2122 2025 2158
rect 1910 2022 1913 2058
rect 1902 1962 1905 1978
rect 1894 1952 1897 1958
rect 1902 1952 1905 1958
rect 1902 1932 1905 1938
rect 1910 1932 1913 1968
rect 1918 1932 1921 1968
rect 1902 1892 1905 1898
rect 1922 1858 1926 1861
rect 1910 1852 1913 1858
rect 1934 1851 1937 2068
rect 1974 2022 1977 2058
rect 1990 2002 1993 2018
rect 2014 2002 2017 2018
rect 2022 2012 2025 2118
rect 2030 2011 2033 2328
rect 2038 2272 2041 2338
rect 2054 2332 2057 2338
rect 2046 2262 2049 2318
rect 2054 2282 2057 2288
rect 2062 2271 2065 2358
rect 2070 2352 2073 2438
rect 2078 2332 2081 2448
rect 2110 2432 2113 2458
rect 2150 2442 2153 2458
rect 2110 2352 2113 2428
rect 2158 2422 2161 2458
rect 2090 2338 2094 2341
rect 2072 2303 2074 2307
rect 2078 2303 2081 2307
rect 2085 2303 2088 2307
rect 2062 2268 2073 2271
rect 2070 2262 2073 2268
rect 2058 2258 2065 2261
rect 2062 2252 2065 2258
rect 2054 2182 2057 2248
rect 2062 2192 2065 2218
rect 2046 2162 2049 2178
rect 2038 2062 2041 2148
rect 2046 2102 2049 2118
rect 2054 2072 2057 2138
rect 2062 2122 2065 2148
rect 2070 2142 2073 2198
rect 2078 2152 2081 2268
rect 2086 2152 2089 2158
rect 2094 2141 2097 2328
rect 2102 2292 2105 2328
rect 2110 2281 2113 2338
rect 2102 2278 2113 2281
rect 2102 2202 2105 2278
rect 2118 2271 2121 2368
rect 2110 2268 2121 2271
rect 2126 2272 2129 2318
rect 2134 2312 2137 2388
rect 2142 2352 2145 2368
rect 2150 2352 2153 2408
rect 2142 2338 2150 2341
rect 2110 2222 2113 2268
rect 2118 2252 2121 2258
rect 2102 2152 2105 2198
rect 2118 2142 2121 2168
rect 2126 2151 2129 2268
rect 2134 2232 2137 2238
rect 2142 2222 2145 2338
rect 2158 2272 2161 2398
rect 2166 2312 2169 2438
rect 2174 2392 2177 2458
rect 2182 2422 2185 2468
rect 2230 2462 2233 2468
rect 2190 2451 2193 2458
rect 2222 2452 2225 2458
rect 2190 2448 2201 2451
rect 2178 2358 2190 2361
rect 2174 2342 2177 2348
rect 2182 2332 2185 2348
rect 2198 2332 2201 2448
rect 2206 2352 2209 2448
rect 2214 2382 2217 2438
rect 2230 2342 2233 2348
rect 2246 2342 2249 2468
rect 2254 2462 2257 2468
rect 2262 2462 2265 2518
rect 2270 2472 2273 2548
rect 2278 2532 2281 2538
rect 2294 2532 2297 2548
rect 2278 2492 2281 2518
rect 2286 2482 2289 2518
rect 2302 2482 2305 2508
rect 2310 2492 2313 2548
rect 2334 2532 2337 2548
rect 2302 2472 2305 2478
rect 2342 2472 2345 2478
rect 2358 2472 2361 2548
rect 2374 2542 2377 2618
rect 2406 2592 2409 2628
rect 2382 2552 2385 2558
rect 2390 2542 2393 2588
rect 2398 2552 2401 2578
rect 2414 2562 2417 2568
rect 2462 2562 2465 2608
rect 2434 2558 2438 2561
rect 2450 2558 2454 2561
rect 2450 2548 2457 2551
rect 2366 2472 2369 2528
rect 2422 2482 2425 2548
rect 2438 2522 2441 2538
rect 2390 2472 2393 2478
rect 2430 2472 2433 2478
rect 2446 2472 2449 2498
rect 2274 2468 2278 2471
rect 2318 2462 2321 2468
rect 2406 2462 2409 2468
rect 2362 2458 2366 2461
rect 2434 2458 2438 2461
rect 2294 2442 2297 2458
rect 2278 2362 2281 2408
rect 2278 2352 2281 2358
rect 2286 2352 2289 2378
rect 2258 2348 2262 2351
rect 2294 2342 2297 2428
rect 2206 2332 2209 2338
rect 2194 2318 2198 2321
rect 2170 2268 2174 2271
rect 2198 2262 2201 2278
rect 2214 2262 2217 2338
rect 2290 2328 2294 2331
rect 2302 2312 2305 2438
rect 2310 2342 2313 2448
rect 2326 2442 2329 2458
rect 2334 2452 2337 2458
rect 2362 2438 2366 2441
rect 2334 2352 2337 2368
rect 2358 2362 2361 2368
rect 2322 2348 2326 2351
rect 2286 2292 2289 2308
rect 2310 2292 2313 2338
rect 2318 2292 2321 2338
rect 2326 2282 2329 2338
rect 2342 2282 2345 2358
rect 2374 2351 2377 2458
rect 2382 2432 2385 2458
rect 2434 2448 2438 2451
rect 2454 2441 2457 2548
rect 2462 2472 2465 2558
rect 2494 2532 2497 2658
rect 2526 2652 2529 2688
rect 2534 2682 2537 2688
rect 2558 2682 2561 2718
rect 2566 2692 2569 2728
rect 2534 2622 2537 2638
rect 2494 2492 2497 2528
rect 2478 2458 2486 2461
rect 2462 2452 2465 2458
rect 2454 2438 2465 2441
rect 2382 2362 2385 2368
rect 2374 2348 2385 2351
rect 2418 2348 2422 2351
rect 2358 2342 2361 2348
rect 2370 2338 2374 2341
rect 2234 2278 2238 2281
rect 2262 2272 2265 2278
rect 2326 2272 2329 2278
rect 2234 2268 2238 2271
rect 2270 2268 2278 2271
rect 2270 2262 2273 2268
rect 2302 2262 2305 2268
rect 2154 2258 2158 2261
rect 2142 2152 2145 2158
rect 2126 2148 2137 2151
rect 2134 2142 2137 2148
rect 2086 2138 2097 2141
rect 2146 2138 2150 2141
rect 2086 2121 2089 2138
rect 2098 2128 2102 2131
rect 2086 2118 2097 2121
rect 2062 2062 2065 2118
rect 2072 2103 2074 2107
rect 2078 2103 2081 2107
rect 2085 2103 2088 2107
rect 2094 2092 2097 2118
rect 2110 2112 2113 2138
rect 2126 2132 2129 2138
rect 2158 2131 2161 2248
rect 2206 2202 2209 2258
rect 2182 2182 2185 2188
rect 2170 2158 2174 2161
rect 2178 2148 2182 2151
rect 2198 2142 2201 2168
rect 2206 2142 2209 2148
rect 2150 2128 2161 2131
rect 2214 2132 2217 2248
rect 2254 2242 2257 2258
rect 2302 2232 2305 2258
rect 2350 2252 2353 2258
rect 2230 2152 2233 2208
rect 2318 2192 2321 2248
rect 2350 2192 2353 2218
rect 2294 2152 2297 2168
rect 2234 2148 2241 2151
rect 2098 2068 2105 2071
rect 2114 2068 2118 2071
rect 2038 2022 2041 2058
rect 2086 2052 2089 2068
rect 2030 2008 2041 2011
rect 1950 1951 1953 1958
rect 1974 1892 1977 1998
rect 2038 1992 2041 2008
rect 2054 1982 2057 2018
rect 2102 1992 2105 2068
rect 2118 2002 2121 2058
rect 2010 1968 2014 1971
rect 2022 1952 2025 1958
rect 2066 1948 2070 1951
rect 2090 1948 2094 1951
rect 1946 1858 1950 1861
rect 1926 1848 1937 1851
rect 1894 1812 1897 1828
rect 1902 1782 1905 1848
rect 1926 1832 1929 1848
rect 1934 1832 1937 1838
rect 1958 1802 1961 1858
rect 1934 1792 1937 1798
rect 1962 1778 1966 1781
rect 1862 1752 1865 1758
rect 1878 1742 1881 1768
rect 1862 1672 1865 1688
rect 1870 1662 1873 1688
rect 1902 1682 1905 1778
rect 1918 1752 1921 1758
rect 1918 1692 1921 1738
rect 1926 1732 1929 1748
rect 1950 1692 1953 1708
rect 1926 1662 1929 1668
rect 1890 1658 1894 1661
rect 1934 1652 1937 1658
rect 1878 1632 1881 1648
rect 1846 1578 1857 1581
rect 1738 1548 1742 1551
rect 1842 1548 1846 1551
rect 1622 1442 1625 1548
rect 1662 1542 1665 1548
rect 1638 1512 1641 1538
rect 1630 1391 1633 1458
rect 1638 1402 1641 1508
rect 1670 1492 1673 1508
rect 1686 1492 1689 1548
rect 1694 1532 1697 1538
rect 1682 1468 1686 1471
rect 1702 1462 1705 1488
rect 1710 1472 1713 1548
rect 1734 1462 1737 1488
rect 1630 1388 1638 1391
rect 1670 1382 1673 1418
rect 1678 1392 1681 1438
rect 1694 1372 1697 1448
rect 1658 1358 1662 1361
rect 1582 1352 1585 1358
rect 1702 1352 1705 1428
rect 1742 1402 1745 1458
rect 1750 1452 1753 1458
rect 1758 1442 1761 1548
rect 1782 1542 1785 1548
rect 1798 1542 1801 1548
rect 1806 1502 1809 1548
rect 1846 1512 1849 1528
rect 1810 1488 1814 1491
rect 1786 1468 1790 1471
rect 1766 1462 1769 1468
rect 1790 1432 1793 1458
rect 1810 1448 1814 1451
rect 1818 1438 1822 1441
rect 1710 1372 1713 1378
rect 1710 1352 1713 1358
rect 1726 1352 1729 1398
rect 1758 1352 1761 1408
rect 1838 1362 1841 1368
rect 1826 1358 1830 1361
rect 1594 1348 1598 1351
rect 1770 1348 1774 1351
rect 1834 1348 1838 1351
rect 1562 1338 1566 1341
rect 1550 1322 1553 1328
rect 1614 1302 1617 1348
rect 1630 1342 1633 1348
rect 1574 1282 1577 1288
rect 1630 1272 1633 1288
rect 1610 1268 1614 1271
rect 1422 1192 1425 1238
rect 1454 1212 1457 1238
rect 1494 1202 1497 1238
rect 1458 1158 1462 1161
rect 1422 1152 1425 1158
rect 1438 1152 1441 1158
rect 1386 1148 1390 1151
rect 1402 1128 1406 1131
rect 1350 1122 1353 1128
rect 1282 1058 1289 1061
rect 1310 1062 1313 1068
rect 1222 1028 1233 1031
rect 1222 992 1225 1028
rect 1214 942 1217 968
rect 1150 862 1153 868
rect 1166 862 1169 878
rect 1182 862 1185 918
rect 1166 852 1169 858
rect 1062 752 1065 758
rect 1126 752 1129 758
rect 1090 748 1094 751
rect 1042 738 1046 741
rect 1048 703 1050 707
rect 1054 703 1057 707
rect 1061 703 1064 707
rect 1026 698 1033 701
rect 1022 682 1025 698
rect 1030 662 1033 668
rect 926 572 929 578
rect 846 552 849 568
rect 906 558 910 561
rect 886 552 889 558
rect 926 552 929 558
rect 942 552 945 558
rect 990 552 993 558
rect 998 552 1001 618
rect 874 548 878 551
rect 862 542 865 548
rect 850 538 854 541
rect 890 528 894 531
rect 886 492 889 508
rect 918 492 921 548
rect 930 538 934 541
rect 950 502 953 548
rect 974 492 977 548
rect 1006 492 1009 608
rect 1038 592 1041 678
rect 1070 622 1073 748
rect 1094 592 1097 738
rect 1102 692 1105 748
rect 1150 742 1153 768
rect 1182 752 1185 768
rect 1130 738 1134 741
rect 1110 672 1113 718
rect 1110 652 1113 658
rect 1126 592 1129 728
rect 1150 692 1153 728
rect 1166 672 1169 708
rect 1138 668 1142 671
rect 1134 652 1137 658
rect 1142 652 1145 658
rect 1014 552 1017 558
rect 1014 532 1017 538
rect 1022 492 1025 558
rect 1078 552 1081 568
rect 1034 548 1038 551
rect 1066 548 1070 551
rect 1146 548 1150 551
rect 1042 538 1046 541
rect 694 452 697 458
rect 666 338 670 341
rect 638 272 641 278
rect 614 262 617 268
rect 598 242 601 258
rect 606 252 609 258
rect 614 242 617 248
rect 630 242 633 258
rect 642 248 646 251
rect 654 251 657 328
rect 694 321 697 358
rect 710 342 713 458
rect 758 412 761 468
rect 766 462 769 468
rect 766 442 769 448
rect 734 342 737 348
rect 694 318 705 321
rect 702 292 705 318
rect 666 268 670 271
rect 690 268 694 271
rect 710 262 713 338
rect 718 272 721 288
rect 726 272 729 308
rect 734 262 737 278
rect 774 262 777 458
rect 790 452 793 478
rect 902 472 905 488
rect 942 472 945 478
rect 930 468 934 471
rect 806 462 809 468
rect 782 442 785 448
rect 806 442 809 448
rect 790 392 793 418
rect 814 392 817 468
rect 838 462 841 468
rect 822 442 825 448
rect 822 422 825 438
rect 806 352 809 368
rect 830 362 833 458
rect 838 392 841 438
rect 846 412 849 468
rect 874 458 878 461
rect 854 422 857 458
rect 906 448 910 451
rect 886 441 889 448
rect 878 438 889 441
rect 854 392 857 408
rect 870 352 873 418
rect 782 272 785 348
rect 818 338 822 341
rect 866 338 870 341
rect 798 332 801 338
rect 654 248 662 251
rect 630 162 633 238
rect 582 152 585 158
rect 598 152 601 158
rect 638 152 641 168
rect 574 122 577 138
rect 534 92 537 98
rect 566 82 569 118
rect 502 72 505 78
rect 566 62 569 68
rect 598 62 601 118
rect 614 72 617 138
rect 646 92 649 158
rect 654 102 657 248
rect 670 202 673 258
rect 686 182 689 258
rect 694 192 697 218
rect 686 122 689 178
rect 702 172 705 248
rect 702 162 705 168
rect 706 148 710 151
rect 654 52 657 88
rect 718 82 721 248
rect 758 222 761 238
rect 734 172 737 218
rect 758 172 761 208
rect 774 162 777 258
rect 782 192 785 258
rect 798 252 801 268
rect 814 252 817 259
rect 790 161 793 198
rect 782 158 793 161
rect 774 152 777 158
rect 746 148 750 151
rect 738 138 742 141
rect 750 72 753 98
rect 714 59 718 62
rect 758 62 761 68
rect 766 62 769 68
rect 782 52 785 158
rect 798 152 801 238
rect 830 222 833 328
rect 846 192 849 328
rect 878 292 881 438
rect 926 432 929 458
rect 934 392 937 448
rect 950 442 953 468
rect 998 462 1001 468
rect 962 458 966 461
rect 886 292 889 358
rect 910 352 913 368
rect 894 252 897 318
rect 910 272 913 338
rect 918 282 921 338
rect 950 332 953 338
rect 914 268 918 271
rect 910 252 913 259
rect 878 212 881 218
rect 854 162 857 168
rect 822 152 825 158
rect 838 152 841 158
rect 918 152 921 268
rect 926 202 929 328
rect 974 312 977 348
rect 982 292 985 448
rect 1014 442 1017 478
rect 1014 372 1017 428
rect 1022 391 1025 438
rect 1030 412 1033 528
rect 1102 522 1105 548
rect 1154 538 1158 541
rect 1048 503 1050 507
rect 1054 503 1057 507
rect 1061 503 1064 507
rect 1070 491 1073 518
rect 1066 488 1073 491
rect 1086 472 1089 478
rect 1042 468 1046 471
rect 1078 462 1081 468
rect 1022 388 1030 391
rect 1054 332 1057 448
rect 1062 392 1065 418
rect 1078 392 1081 448
rect 1102 432 1105 468
rect 1166 462 1169 658
rect 1190 592 1193 908
rect 1198 872 1201 938
rect 1206 902 1209 918
rect 1214 872 1217 908
rect 1222 892 1225 978
rect 1258 958 1262 961
rect 1238 942 1241 958
rect 1258 948 1262 951
rect 1246 932 1249 948
rect 1278 942 1281 1058
rect 1286 1042 1289 1048
rect 1294 1042 1297 1048
rect 1298 947 1302 950
rect 1230 892 1233 928
rect 1258 888 1262 891
rect 1294 872 1297 928
rect 1250 868 1254 871
rect 1242 858 1246 861
rect 1198 852 1201 858
rect 1302 792 1305 868
rect 1310 852 1313 1058
rect 1326 1012 1329 1068
rect 1350 1052 1353 1058
rect 1358 992 1361 1128
rect 1374 1102 1377 1128
rect 1386 1118 1390 1121
rect 1406 1092 1409 1098
rect 1414 1082 1417 1118
rect 1430 1072 1433 1148
rect 1446 1132 1449 1158
rect 1454 1092 1457 1148
rect 1462 1132 1465 1148
rect 1470 1142 1473 1178
rect 1482 1158 1486 1161
rect 1498 1148 1502 1151
rect 1478 1142 1481 1148
rect 1510 1142 1513 1178
rect 1518 1152 1521 1188
rect 1502 1131 1505 1138
rect 1518 1132 1521 1148
rect 1502 1128 1513 1131
rect 1474 1088 1478 1091
rect 1450 1068 1454 1071
rect 1438 1052 1441 1058
rect 1418 1048 1422 1051
rect 1406 992 1409 1018
rect 1398 972 1401 978
rect 1462 972 1465 1048
rect 1502 1042 1505 1058
rect 1398 962 1401 968
rect 1442 958 1446 961
rect 1366 952 1369 958
rect 1442 948 1446 951
rect 1358 912 1361 928
rect 1382 922 1385 948
rect 1318 863 1321 898
rect 1350 872 1353 878
rect 1334 862 1337 868
rect 1358 862 1361 908
rect 1374 892 1377 898
rect 1234 778 1238 781
rect 1294 772 1297 778
rect 1250 768 1254 771
rect 1266 758 1270 761
rect 1282 758 1286 761
rect 1246 752 1249 758
rect 1238 742 1241 748
rect 1266 738 1270 741
rect 1230 662 1233 668
rect 1246 662 1249 668
rect 1270 662 1273 678
rect 1278 652 1281 748
rect 1302 732 1305 758
rect 1322 738 1326 741
rect 1310 682 1313 728
rect 1198 558 1206 561
rect 1178 548 1182 551
rect 1182 532 1185 538
rect 1190 532 1193 548
rect 1198 492 1201 558
rect 1206 472 1209 478
rect 1214 472 1217 538
rect 1118 452 1121 459
rect 1070 342 1073 368
rect 1094 362 1097 368
rect 1006 292 1009 308
rect 970 288 974 291
rect 982 272 985 278
rect 994 258 998 261
rect 1014 252 1017 328
rect 1030 252 1033 258
rect 946 168 950 171
rect 850 148 854 151
rect 994 148 998 151
rect 790 142 793 148
rect 894 142 897 148
rect 818 138 822 141
rect 798 132 801 138
rect 790 62 793 118
rect 798 112 801 128
rect 830 122 833 138
rect 806 72 809 88
rect 870 62 873 138
rect 906 88 910 91
rect 910 72 913 78
rect 918 62 921 98
rect 938 68 942 71
rect 794 58 798 61
rect 850 58 854 61
rect 930 58 934 61
rect 954 58 958 61
rect 966 52 969 88
rect 982 82 985 128
rect 982 72 985 78
rect 1006 62 1009 78
rect 1030 62 1033 248
rect 1038 201 1041 328
rect 1048 303 1050 307
rect 1054 303 1057 307
rect 1061 303 1064 307
rect 1070 292 1073 328
rect 1062 272 1065 288
rect 1078 281 1081 348
rect 1102 342 1105 398
rect 1182 392 1185 418
rect 1114 368 1118 371
rect 1126 362 1129 388
rect 1214 381 1217 468
rect 1222 462 1225 648
rect 1230 441 1233 608
rect 1270 592 1273 618
rect 1246 552 1249 558
rect 1238 512 1241 548
rect 1254 472 1257 548
rect 1262 462 1265 568
rect 1278 552 1281 578
rect 1294 552 1297 648
rect 1318 642 1321 738
rect 1334 672 1337 808
rect 1358 772 1361 858
rect 1382 852 1385 888
rect 1390 852 1393 938
rect 1398 862 1401 918
rect 1422 892 1425 938
rect 1430 912 1433 918
rect 1462 902 1465 918
rect 1426 878 1430 881
rect 1454 872 1457 878
rect 1406 852 1409 868
rect 1434 858 1438 861
rect 1390 792 1393 808
rect 1326 632 1329 638
rect 1334 602 1337 668
rect 1342 662 1345 768
rect 1406 762 1409 768
rect 1422 752 1425 758
rect 1430 752 1433 818
rect 1462 762 1465 768
rect 1470 762 1473 958
rect 1478 932 1481 938
rect 1486 872 1489 1038
rect 1510 992 1513 1128
rect 1526 1072 1529 1268
rect 1542 1263 1545 1268
rect 1638 1262 1641 1348
rect 1602 1258 1606 1261
rect 1634 1258 1638 1261
rect 1646 1252 1649 1328
rect 1654 1272 1657 1348
rect 1686 1272 1689 1278
rect 1662 1262 1665 1268
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1573 1203 1576 1207
rect 1586 1168 1590 1171
rect 1534 1162 1537 1168
rect 1562 1158 1566 1161
rect 1562 1148 1566 1151
rect 1562 1138 1566 1141
rect 1534 1063 1537 1068
rect 1566 1052 1569 1088
rect 1598 1062 1601 1188
rect 1638 1082 1641 1208
rect 1646 1152 1649 1158
rect 1654 1092 1657 1128
rect 1670 1102 1673 1268
rect 1678 1252 1681 1258
rect 1694 1192 1697 1348
rect 1702 1322 1705 1348
rect 1734 1332 1737 1338
rect 1742 1332 1745 1348
rect 1790 1342 1793 1348
rect 1798 1342 1801 1348
rect 1806 1342 1809 1348
rect 1834 1338 1841 1341
rect 1730 1288 1734 1291
rect 1710 1282 1713 1288
rect 1750 1282 1753 1318
rect 1726 1262 1729 1278
rect 1706 1258 1710 1261
rect 1786 1258 1790 1261
rect 1766 1242 1769 1258
rect 1758 1192 1761 1218
rect 1698 1148 1702 1151
rect 1722 1138 1726 1141
rect 1686 1132 1689 1138
rect 1734 1102 1737 1158
rect 1750 1152 1753 1168
rect 1790 1152 1793 1158
rect 1774 1131 1777 1148
rect 1782 1142 1785 1148
rect 1774 1128 1785 1131
rect 1638 1072 1641 1078
rect 1646 1072 1649 1078
rect 1662 1072 1665 1098
rect 1682 1068 1686 1071
rect 1598 1042 1601 1048
rect 1606 1032 1609 1068
rect 1614 1062 1617 1068
rect 1614 1042 1617 1048
rect 1622 1031 1625 1068
rect 1614 1028 1625 1031
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1573 1003 1576 1007
rect 1614 992 1617 1028
rect 1630 992 1633 1028
rect 1562 968 1566 971
rect 1618 968 1622 971
rect 1522 958 1526 961
rect 1594 958 1598 961
rect 1494 942 1497 948
rect 1502 942 1505 958
rect 1586 948 1590 951
rect 1522 938 1526 941
rect 1502 892 1505 938
rect 1502 872 1505 888
rect 1478 862 1481 868
rect 1354 748 1358 751
rect 1370 748 1374 751
rect 1350 732 1353 738
rect 1390 732 1393 748
rect 1410 738 1414 741
rect 1350 672 1353 678
rect 1366 661 1369 728
rect 1390 672 1393 718
rect 1438 712 1441 758
rect 1446 742 1449 748
rect 1450 738 1454 741
rect 1406 692 1409 708
rect 1414 672 1417 678
rect 1422 662 1425 668
rect 1430 662 1433 698
rect 1446 692 1449 728
rect 1454 702 1457 718
rect 1462 672 1465 678
rect 1358 658 1369 661
rect 1318 562 1321 568
rect 1342 552 1345 658
rect 1358 572 1361 658
rect 1382 652 1385 658
rect 1370 638 1374 641
rect 1354 568 1358 571
rect 1334 542 1337 548
rect 1290 538 1294 541
rect 1350 492 1353 538
rect 1398 532 1401 638
rect 1446 632 1449 648
rect 1478 642 1481 718
rect 1486 672 1489 868
rect 1518 772 1521 828
rect 1526 792 1529 928
rect 1534 922 1537 948
rect 1602 938 1606 941
rect 1534 902 1537 918
rect 1538 888 1542 891
rect 1542 852 1545 868
rect 1550 862 1553 898
rect 1566 852 1569 888
rect 1574 862 1577 868
rect 1598 861 1601 908
rect 1606 892 1609 928
rect 1630 892 1633 988
rect 1638 942 1641 1068
rect 1658 1058 1662 1061
rect 1646 1051 1649 1058
rect 1646 1048 1657 1051
rect 1654 1002 1657 1048
rect 1706 1038 1710 1041
rect 1654 892 1657 998
rect 1718 992 1721 1098
rect 1734 1062 1737 1088
rect 1766 1063 1769 1078
rect 1678 952 1681 958
rect 1702 942 1705 948
rect 1734 942 1737 1058
rect 1758 952 1761 1018
rect 1774 992 1777 1008
rect 1774 952 1777 958
rect 1730 928 1737 931
rect 1678 892 1681 898
rect 1614 872 1617 878
rect 1642 868 1646 871
rect 1706 868 1710 871
rect 1598 858 1606 861
rect 1534 742 1537 748
rect 1498 738 1502 741
rect 1510 728 1518 731
rect 1494 662 1497 668
rect 1502 662 1505 718
rect 1470 572 1473 578
rect 1410 548 1414 551
rect 1414 532 1417 538
rect 1278 472 1281 478
rect 1346 468 1350 471
rect 1230 438 1238 441
rect 1222 402 1225 418
rect 1230 391 1233 438
rect 1246 431 1249 448
rect 1226 388 1233 391
rect 1238 428 1249 431
rect 1206 378 1217 381
rect 1166 352 1169 368
rect 1110 342 1113 348
rect 1102 292 1105 338
rect 1070 278 1081 281
rect 1070 262 1073 278
rect 1110 272 1113 328
rect 1082 268 1086 271
rect 1150 262 1153 268
rect 1174 262 1177 338
rect 1206 332 1209 378
rect 1218 368 1225 371
rect 1222 351 1225 368
rect 1230 362 1233 368
rect 1222 348 1230 351
rect 1238 341 1241 428
rect 1270 422 1273 468
rect 1346 438 1350 441
rect 1246 352 1249 368
rect 1286 352 1289 368
rect 1326 352 1329 368
rect 1238 338 1249 341
rect 1206 292 1209 298
rect 1062 242 1065 248
rect 1078 202 1081 238
rect 1038 198 1046 201
rect 1046 192 1049 198
rect 1062 142 1065 158
rect 1070 152 1073 188
rect 1094 162 1097 258
rect 1102 252 1105 258
rect 1090 148 1094 151
rect 1062 132 1065 138
rect 1048 103 1050 107
rect 1054 103 1057 107
rect 1061 103 1064 107
rect 1070 92 1073 108
rect 1070 62 1073 68
rect 1110 62 1113 218
rect 1174 172 1177 258
rect 1214 232 1217 268
rect 1222 262 1225 318
rect 1246 292 1249 338
rect 1234 268 1238 271
rect 1238 252 1241 258
rect 1194 178 1198 181
rect 1206 152 1209 198
rect 1246 182 1249 248
rect 1254 232 1257 338
rect 1302 332 1305 338
rect 1262 272 1265 308
rect 1270 282 1273 318
rect 1342 292 1345 428
rect 1270 262 1273 268
rect 1278 262 1281 268
rect 1302 262 1305 268
rect 1326 262 1329 278
rect 1334 262 1337 278
rect 1354 268 1358 271
rect 1282 248 1286 251
rect 1298 248 1302 251
rect 1222 172 1225 178
rect 1138 148 1142 151
rect 1126 72 1129 128
rect 1198 122 1201 138
rect 1126 62 1129 68
rect 1150 62 1153 98
rect 1214 91 1217 168
rect 1254 162 1257 208
rect 1294 162 1297 238
rect 1326 222 1329 258
rect 1310 202 1313 218
rect 1230 142 1233 148
rect 1254 142 1257 158
rect 1270 152 1273 158
rect 1262 142 1265 148
rect 1278 101 1281 138
rect 1294 112 1297 158
rect 1310 152 1313 198
rect 1334 152 1337 178
rect 1350 152 1353 258
rect 1358 172 1361 258
rect 1330 138 1334 141
rect 1318 122 1321 138
rect 1270 98 1281 101
rect 1210 88 1217 91
rect 1222 62 1225 68
rect 1246 62 1249 88
rect 1270 82 1273 98
rect 1302 92 1305 108
rect 1342 102 1345 138
rect 1358 112 1361 128
rect 1326 82 1329 88
rect 1358 82 1361 108
rect 1366 72 1369 478
rect 1382 462 1385 468
rect 1398 392 1401 518
rect 1414 482 1417 528
rect 1454 492 1457 558
rect 1478 552 1481 618
rect 1494 592 1497 628
rect 1510 612 1513 728
rect 1542 722 1545 848
rect 1550 822 1553 838
rect 1550 772 1553 818
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1573 803 1576 807
rect 1558 742 1561 788
rect 1542 642 1545 658
rect 1486 552 1489 558
rect 1502 542 1505 588
rect 1478 522 1481 538
rect 1514 518 1518 521
rect 1462 472 1465 478
rect 1494 472 1497 478
rect 1526 472 1529 598
rect 1538 548 1542 551
rect 1534 512 1537 548
rect 1414 463 1417 468
rect 1502 462 1505 468
rect 1518 462 1521 468
rect 1426 388 1430 391
rect 1386 368 1390 371
rect 1398 282 1401 378
rect 1410 368 1414 371
rect 1438 362 1441 388
rect 1446 382 1449 448
rect 1470 442 1473 448
rect 1486 442 1489 448
rect 1458 368 1462 371
rect 1458 348 1462 351
rect 1422 342 1425 348
rect 1430 342 1433 348
rect 1374 252 1377 258
rect 1374 142 1377 148
rect 1382 142 1385 218
rect 1398 192 1401 268
rect 1414 262 1417 328
rect 1430 312 1433 338
rect 1462 332 1465 338
rect 1470 321 1473 348
rect 1494 342 1497 458
rect 1502 442 1505 448
rect 1502 352 1505 398
rect 1510 341 1513 378
rect 1506 338 1513 341
rect 1502 332 1505 338
rect 1470 318 1478 321
rect 1518 292 1521 448
rect 1526 392 1529 468
rect 1542 412 1545 418
rect 1550 382 1553 718
rect 1566 672 1569 688
rect 1574 662 1577 778
rect 1590 742 1593 758
rect 1590 702 1593 718
rect 1598 672 1601 838
rect 1606 682 1609 858
rect 1614 772 1617 848
rect 1622 792 1625 868
rect 1714 858 1718 861
rect 1694 852 1697 858
rect 1642 848 1646 851
rect 1638 752 1641 838
rect 1662 832 1665 848
rect 1654 782 1657 818
rect 1658 768 1662 771
rect 1694 762 1697 848
rect 1710 802 1713 818
rect 1706 778 1710 781
rect 1686 752 1689 758
rect 1718 752 1721 768
rect 1726 752 1729 908
rect 1734 852 1737 928
rect 1742 872 1745 918
rect 1766 902 1769 938
rect 1754 868 1758 871
rect 1734 792 1737 848
rect 1750 842 1753 858
rect 1766 851 1769 868
rect 1774 862 1777 918
rect 1782 872 1785 1128
rect 1798 1122 1801 1338
rect 1814 1262 1817 1338
rect 1830 1332 1833 1338
rect 1838 1202 1841 1338
rect 1846 1322 1849 1448
rect 1854 1412 1857 1578
rect 1870 1561 1873 1618
rect 1870 1558 1878 1561
rect 1894 1552 1897 1628
rect 1922 1588 1926 1591
rect 1918 1552 1921 1578
rect 1950 1562 1953 1618
rect 1902 1542 1905 1548
rect 1918 1542 1921 1548
rect 1874 1538 1878 1541
rect 1862 1442 1865 1528
rect 1870 1452 1873 1468
rect 1878 1463 1881 1518
rect 1918 1492 1921 1528
rect 1934 1492 1937 1558
rect 1946 1548 1950 1551
rect 1942 1532 1945 1538
rect 1958 1512 1961 1748
rect 1974 1702 1977 1818
rect 1982 1772 1985 1948
rect 2030 1932 2033 1948
rect 2054 1902 2057 1948
rect 2072 1903 2074 1907
rect 2078 1903 2081 1907
rect 2085 1903 2088 1907
rect 2110 1902 2113 1998
rect 2034 1878 2038 1881
rect 2018 1858 2022 1861
rect 2058 1858 2062 1861
rect 1998 1682 2001 1818
rect 2022 1742 2025 1748
rect 2046 1742 2049 1768
rect 2018 1688 2022 1691
rect 1978 1658 1982 1661
rect 1966 1552 1969 1558
rect 1974 1542 1977 1548
rect 1990 1522 1993 1558
rect 1982 1518 1990 1521
rect 1974 1492 1977 1518
rect 1982 1492 1985 1518
rect 1854 1292 1857 1358
rect 1870 1342 1873 1448
rect 1894 1332 1897 1348
rect 1886 1272 1889 1328
rect 1854 1263 1857 1268
rect 1838 1182 1841 1198
rect 1810 1168 1814 1171
rect 1874 1168 1878 1171
rect 1806 1152 1809 1158
rect 1830 1132 1833 1168
rect 1838 1122 1841 1138
rect 1830 1082 1833 1088
rect 1818 1068 1822 1071
rect 1838 1061 1841 1078
rect 1834 1058 1841 1061
rect 1826 1048 1830 1051
rect 1798 1042 1801 1048
rect 1814 1042 1817 1048
rect 1790 932 1793 958
rect 1806 952 1809 968
rect 1838 962 1841 968
rect 1826 958 1830 961
rect 1826 948 1830 951
rect 1798 912 1801 938
rect 1830 932 1833 938
rect 1790 861 1793 898
rect 1806 892 1809 928
rect 1802 868 1806 871
rect 1818 868 1822 871
rect 1782 858 1793 861
rect 1766 848 1777 851
rect 1774 792 1777 848
rect 1782 792 1785 858
rect 1802 848 1809 851
rect 1806 792 1809 848
rect 1814 832 1817 848
rect 1818 788 1822 791
rect 1758 752 1761 758
rect 1586 668 1590 671
rect 1590 642 1593 648
rect 1598 631 1601 668
rect 1606 652 1609 658
rect 1590 628 1601 631
rect 1606 632 1609 638
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1573 603 1576 607
rect 1566 532 1569 538
rect 1590 492 1593 628
rect 1598 542 1601 548
rect 1614 492 1617 718
rect 1622 662 1625 738
rect 1630 702 1633 738
rect 1646 732 1649 748
rect 1670 732 1673 748
rect 1678 741 1681 748
rect 1694 741 1697 748
rect 1678 738 1697 741
rect 1638 671 1641 708
rect 1654 692 1657 728
rect 1702 692 1705 748
rect 1798 742 1801 758
rect 1818 738 1822 741
rect 1770 728 1777 731
rect 1634 668 1641 671
rect 1674 668 1678 671
rect 1690 668 1694 671
rect 1622 652 1625 658
rect 1646 642 1649 648
rect 1630 482 1633 638
rect 1662 592 1665 668
rect 1674 658 1678 661
rect 1702 602 1705 648
rect 1650 588 1654 591
rect 1702 572 1705 588
rect 1674 558 1678 561
rect 1694 552 1697 558
rect 1682 548 1686 551
rect 1670 542 1673 548
rect 1558 462 1561 468
rect 1606 462 1609 468
rect 1646 462 1649 528
rect 1618 438 1622 441
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1573 403 1576 407
rect 1526 362 1529 368
rect 1542 362 1545 368
rect 1542 342 1545 348
rect 1526 322 1529 328
rect 1534 312 1537 338
rect 1542 322 1545 338
rect 1502 272 1505 278
rect 1526 272 1529 278
rect 1534 272 1537 278
rect 1482 268 1486 271
rect 1446 263 1449 268
rect 1430 172 1433 188
rect 1462 162 1465 268
rect 1498 258 1502 261
rect 1478 252 1481 258
rect 1454 152 1457 158
rect 1410 148 1414 151
rect 1446 142 1449 148
rect 1462 142 1465 148
rect 1478 142 1481 158
rect 1498 147 1502 150
rect 1410 138 1414 141
rect 1322 68 1326 71
rect 1342 62 1345 68
rect 1306 58 1310 61
rect 1390 52 1393 128
rect 1406 122 1409 138
rect 1510 132 1513 248
rect 1446 62 1449 68
rect 1470 62 1473 98
rect 1494 72 1497 78
rect 1426 58 1430 61
rect 1526 52 1529 88
rect 1542 72 1545 298
rect 1550 272 1553 378
rect 1654 372 1657 528
rect 1686 502 1689 548
rect 1698 538 1702 541
rect 1710 522 1713 668
rect 1742 662 1745 718
rect 1766 672 1769 688
rect 1722 658 1726 661
rect 1754 658 1758 661
rect 1718 652 1721 658
rect 1762 648 1766 651
rect 1734 642 1737 648
rect 1774 642 1777 728
rect 1770 638 1774 641
rect 1766 552 1769 558
rect 1722 548 1726 551
rect 1722 538 1726 541
rect 1678 463 1681 478
rect 1726 471 1729 538
rect 1742 532 1745 538
rect 1758 502 1761 528
rect 1742 482 1745 488
rect 1726 468 1734 471
rect 1758 462 1761 498
rect 1766 472 1769 478
rect 1774 462 1777 478
rect 1722 458 1726 461
rect 1738 448 1742 451
rect 1710 442 1713 448
rect 1726 442 1729 448
rect 1782 422 1785 458
rect 1694 392 1697 418
rect 1718 392 1721 408
rect 1790 392 1793 728
rect 1806 572 1809 658
rect 1822 652 1825 658
rect 1818 568 1822 571
rect 1806 552 1809 568
rect 1830 542 1833 928
rect 1838 892 1841 948
rect 1846 912 1849 1148
rect 1854 1121 1857 1148
rect 1894 1142 1897 1198
rect 1902 1192 1905 1348
rect 1910 1292 1913 1478
rect 1930 1468 1934 1471
rect 1950 1451 1953 1468
rect 1962 1458 1966 1461
rect 1950 1448 1961 1451
rect 1942 1342 1945 1448
rect 1958 1392 1961 1448
rect 1974 1362 1977 1448
rect 1990 1392 1993 1508
rect 1982 1352 1985 1368
rect 1942 1292 1945 1328
rect 1954 1318 1961 1321
rect 1914 1288 1918 1291
rect 1926 1272 1929 1278
rect 1926 1212 1929 1258
rect 1902 1152 1905 1188
rect 1930 1168 1934 1171
rect 1930 1148 1934 1151
rect 1866 1128 1870 1131
rect 1854 1118 1865 1121
rect 1862 1092 1865 1118
rect 1894 1092 1897 1138
rect 1870 1071 1873 1088
rect 1902 1082 1905 1148
rect 1910 1112 1913 1118
rect 1950 1072 1953 1298
rect 1958 1282 1961 1318
rect 1966 1251 1969 1328
rect 1990 1292 1993 1358
rect 1998 1282 2001 1668
rect 2030 1662 2033 1738
rect 2038 1662 2041 1678
rect 2046 1652 2049 1658
rect 2006 1532 2009 1548
rect 2014 1471 2017 1618
rect 2022 1592 2025 1648
rect 2054 1552 2057 1558
rect 2042 1548 2046 1551
rect 2030 1532 2033 1548
rect 2014 1468 2025 1471
rect 2014 1452 2017 1458
rect 2006 1352 2009 1358
rect 2014 1352 2017 1358
rect 2022 1292 2025 1468
rect 2038 1462 2041 1488
rect 2062 1412 2065 1818
rect 2082 1728 2086 1731
rect 2072 1703 2074 1707
rect 2078 1703 2081 1707
rect 2085 1703 2088 1707
rect 2086 1662 2089 1668
rect 2070 1592 2073 1658
rect 2078 1592 2081 1658
rect 2094 1642 2097 1898
rect 2102 1752 2105 1858
rect 2118 1842 2121 1848
rect 2126 1842 2129 1948
rect 2134 1862 2137 2008
rect 2142 1992 2145 2008
rect 2142 1882 2145 1918
rect 2142 1852 2145 1858
rect 2102 1742 2105 1748
rect 2134 1742 2137 1748
rect 2114 1728 2118 1731
rect 2110 1622 2113 1728
rect 2134 1672 2137 1678
rect 2126 1662 2129 1668
rect 2142 1631 2145 1748
rect 2150 1662 2153 2128
rect 2214 2092 2217 2128
rect 2222 2082 2225 2118
rect 2158 2062 2161 2078
rect 2230 2072 2233 2078
rect 2238 2072 2241 2148
rect 2246 2102 2249 2118
rect 2262 2092 2265 2098
rect 2270 2071 2273 2148
rect 2278 2142 2281 2148
rect 2270 2068 2278 2071
rect 2158 2002 2161 2018
rect 2158 1952 2161 1998
rect 2174 1992 2177 2038
rect 2182 2022 2185 2058
rect 2214 1982 2217 1988
rect 2198 1942 2201 1948
rect 2158 1892 2161 1928
rect 2166 1852 2169 1858
rect 2182 1812 2185 1868
rect 2190 1862 2193 1898
rect 2206 1892 2209 1958
rect 2214 1862 2217 1918
rect 2206 1762 2209 1778
rect 2162 1738 2166 1741
rect 2214 1732 2217 1848
rect 2222 1812 2225 2068
rect 2278 2062 2281 2068
rect 2246 2042 2249 2058
rect 2286 2002 2289 2148
rect 2302 2142 2305 2148
rect 2294 2092 2297 2118
rect 2318 2092 2321 2098
rect 2334 2092 2337 2158
rect 2350 2152 2353 2158
rect 2318 2072 2321 2088
rect 2358 2082 2361 2308
rect 2382 2302 2385 2348
rect 2382 2292 2385 2298
rect 2430 2292 2433 2428
rect 2370 2268 2374 2271
rect 2406 2262 2409 2268
rect 2370 2158 2374 2161
rect 2310 2062 2313 2068
rect 2342 2062 2345 2078
rect 2378 2068 2382 2071
rect 2350 2062 2353 2068
rect 2374 2052 2377 2058
rect 2230 1952 2233 1998
rect 2242 1978 2246 1981
rect 2286 1952 2289 1998
rect 2294 1992 2297 2018
rect 2310 1972 2313 2018
rect 2294 1942 2297 1968
rect 2334 1942 2337 2048
rect 2382 2022 2385 2058
rect 2390 2002 2393 2218
rect 2430 2182 2433 2218
rect 2438 2181 2441 2338
rect 2446 2272 2449 2398
rect 2446 2262 2449 2268
rect 2438 2178 2446 2181
rect 2438 2142 2441 2148
rect 2446 2142 2449 2178
rect 2462 2092 2465 2438
rect 2470 2392 2473 2458
rect 2478 2452 2481 2458
rect 2470 2382 2473 2388
rect 2482 2358 2486 2361
rect 2494 2342 2497 2488
rect 2502 2472 2505 2578
rect 2510 2522 2513 2548
rect 2534 2492 2537 2508
rect 2550 2492 2553 2668
rect 2590 2632 2593 2718
rect 2598 2662 2601 2668
rect 2558 2562 2561 2568
rect 2566 2552 2569 2618
rect 2584 2603 2586 2607
rect 2590 2603 2593 2607
rect 2597 2603 2600 2607
rect 2526 2472 2529 2478
rect 2534 2462 2537 2488
rect 2502 2412 2505 2458
rect 2510 2452 2513 2458
rect 2518 2361 2521 2418
rect 2534 2372 2537 2378
rect 2510 2358 2521 2361
rect 2510 2352 2513 2358
rect 2542 2352 2545 2468
rect 2558 2462 2561 2548
rect 2574 2532 2577 2538
rect 2598 2532 2601 2558
rect 2578 2518 2582 2521
rect 2578 2478 2582 2481
rect 2590 2472 2593 2518
rect 2586 2468 2590 2471
rect 2566 2462 2569 2468
rect 2574 2452 2577 2468
rect 2598 2462 2601 2468
rect 2584 2403 2586 2407
rect 2590 2403 2593 2407
rect 2597 2403 2600 2407
rect 2606 2382 2609 2748
rect 2614 2372 2617 2928
rect 2658 2918 2662 2921
rect 2622 2862 2625 2918
rect 2678 2912 2681 2948
rect 2706 2938 2710 2941
rect 2694 2932 2697 2938
rect 2622 2792 2625 2798
rect 2622 2762 2625 2788
rect 2630 2782 2633 2858
rect 2638 2852 2641 2888
rect 2682 2868 2686 2871
rect 2654 2862 2657 2868
rect 2662 2851 2665 2868
rect 2658 2848 2665 2851
rect 2634 2748 2638 2751
rect 2702 2742 2705 2838
rect 2710 2752 2713 2758
rect 2662 2662 2665 2738
rect 2686 2692 2689 2698
rect 2698 2658 2702 2661
rect 2718 2652 2721 3098
rect 2806 3072 2809 3078
rect 2826 3068 2830 3071
rect 2858 3068 2862 3071
rect 2766 3062 2769 3068
rect 2774 3062 2777 3068
rect 2750 2952 2753 2998
rect 2774 2971 2777 3058
rect 2822 3032 2825 3058
rect 2846 3032 2849 3068
rect 2774 2968 2782 2971
rect 2778 2958 2782 2961
rect 2738 2948 2742 2951
rect 2726 2932 2729 2948
rect 2758 2932 2761 2948
rect 2766 2922 2769 2938
rect 2766 2872 2769 2898
rect 2790 2872 2793 2958
rect 2814 2952 2817 2958
rect 2802 2948 2806 2951
rect 2830 2942 2833 2948
rect 2854 2922 2857 3058
rect 2870 3042 2873 3058
rect 2878 3052 2881 3218
rect 2886 3152 2889 3188
rect 2942 3182 2945 3258
rect 2950 3252 2953 3318
rect 2974 3272 2977 3338
rect 2990 3272 2993 3368
rect 3046 3351 3049 3368
rect 3046 3322 3049 3328
rect 3006 3272 3009 3298
rect 3038 3292 3041 3298
rect 3022 3288 3030 3291
rect 2982 3262 2985 3268
rect 2962 3258 2966 3261
rect 2994 3258 2998 3261
rect 2962 3248 2966 3251
rect 2974 3248 2982 3251
rect 2950 3192 2953 3198
rect 2974 3192 2977 3248
rect 3014 3232 3017 3258
rect 2914 3178 2918 3181
rect 2982 3172 2985 3178
rect 2938 3148 2942 3151
rect 2938 3138 2942 3141
rect 2986 3138 2990 3141
rect 2894 3072 2897 3078
rect 2886 3062 2889 3068
rect 2902 3062 2905 3138
rect 2958 3132 2961 3138
rect 2966 3132 2969 3138
rect 2998 3132 3001 3148
rect 3014 3131 3017 3158
rect 3022 3152 3025 3288
rect 3030 3282 3033 3288
rect 3046 3282 3049 3298
rect 3062 3292 3065 3548
rect 3070 3542 3073 3548
rect 3102 3542 3105 3678
rect 3126 3672 3129 3748
rect 3134 3692 3137 3748
rect 3158 3742 3161 3858
rect 3254 3852 3257 3858
rect 3230 3842 3233 3848
rect 3246 3842 3249 3848
rect 3202 3838 3206 3841
rect 3262 3812 3265 3858
rect 3142 3682 3145 3708
rect 3126 3662 3129 3668
rect 3078 3462 3081 3468
rect 3070 3442 3073 3448
rect 3086 3382 3089 3518
rect 3096 3503 3098 3507
rect 3102 3503 3105 3507
rect 3109 3503 3112 3507
rect 3102 3472 3105 3478
rect 3094 3432 3097 3458
rect 3090 3368 3094 3371
rect 3078 3342 3081 3348
rect 3030 3262 3033 3268
rect 3086 3202 3089 3348
rect 3096 3303 3098 3307
rect 3102 3303 3105 3307
rect 3109 3303 3112 3307
rect 3118 3282 3121 3628
rect 3126 3532 3129 3538
rect 3134 3492 3137 3548
rect 3126 3362 3129 3478
rect 3134 3472 3137 3488
rect 3126 3352 3129 3358
rect 3098 3268 3102 3271
rect 3118 3262 3121 3278
rect 3134 3272 3137 3438
rect 3142 3402 3145 3678
rect 3158 3672 3161 3738
rect 3198 3722 3201 3748
rect 3206 3742 3209 3748
rect 3214 3722 3217 3728
rect 3230 3722 3233 3748
rect 3246 3732 3249 3758
rect 3262 3742 3265 3748
rect 3278 3732 3281 3747
rect 3310 3742 3313 3948
rect 3398 3942 3401 3948
rect 3510 3942 3513 3948
rect 3390 3931 3393 3938
rect 3390 3928 3398 3931
rect 3374 3911 3377 3918
rect 3374 3908 3382 3911
rect 3374 3872 3377 3898
rect 3382 3862 3385 3868
rect 3370 3858 3374 3861
rect 3334 3852 3337 3858
rect 3326 3772 3329 3818
rect 3330 3758 3334 3761
rect 3190 3712 3193 3718
rect 3310 3672 3313 3738
rect 3238 3668 3246 3671
rect 3274 3668 3278 3671
rect 3238 3662 3241 3668
rect 3250 3658 3254 3661
rect 3182 3652 3185 3658
rect 3238 3592 3241 3618
rect 3150 3552 3153 3558
rect 3190 3552 3193 3568
rect 3222 3551 3225 3568
rect 3254 3532 3257 3588
rect 3262 3532 3265 3658
rect 3294 3652 3297 3668
rect 3334 3662 3337 3708
rect 3310 3592 3313 3628
rect 3286 3562 3289 3568
rect 3270 3552 3273 3558
rect 3154 3518 3158 3521
rect 3166 3471 3169 3518
rect 3262 3512 3265 3518
rect 3262 3502 3265 3508
rect 3162 3468 3169 3471
rect 3206 3472 3209 3498
rect 3286 3492 3289 3548
rect 3302 3542 3305 3588
rect 3326 3552 3329 3558
rect 3334 3542 3337 3548
rect 3342 3542 3345 3858
rect 3398 3852 3401 3908
rect 3414 3862 3417 3868
rect 3422 3862 3425 3938
rect 3446 3932 3449 3938
rect 3430 3872 3433 3878
rect 3446 3862 3449 3868
rect 3470 3862 3473 3868
rect 3486 3862 3489 3918
rect 3502 3882 3505 3908
rect 3510 3862 3513 3928
rect 3526 3862 3529 3868
rect 3490 3858 3494 3861
rect 3350 3842 3353 3848
rect 3358 3792 3361 3818
rect 3366 3792 3369 3818
rect 3374 3762 3377 3768
rect 3382 3752 3385 3808
rect 3414 3792 3417 3828
rect 3390 3752 3393 3778
rect 3402 3748 3406 3751
rect 3362 3738 3366 3741
rect 3398 3702 3401 3738
rect 3374 3612 3377 3698
rect 3394 3688 3398 3691
rect 3406 3672 3409 3718
rect 3414 3692 3417 3708
rect 3422 3702 3425 3728
rect 3430 3712 3433 3718
rect 3430 3682 3433 3688
rect 3438 3671 3441 3858
rect 3430 3668 3441 3671
rect 3446 3672 3449 3788
rect 3462 3691 3465 3818
rect 3462 3688 3470 3691
rect 3398 3662 3401 3668
rect 3406 3662 3409 3668
rect 3394 3658 3398 3661
rect 3422 3621 3425 3648
rect 3430 3642 3433 3668
rect 3462 3662 3465 3668
rect 3486 3662 3489 3838
rect 3526 3752 3529 3858
rect 3534 3782 3537 3858
rect 3542 3762 3545 3768
rect 3494 3722 3497 3747
rect 3510 3742 3513 3748
rect 3550 3742 3553 4048
rect 3590 4012 3593 4048
rect 3630 4042 3633 4058
rect 3590 3992 3593 4008
rect 3608 4003 3610 4007
rect 3614 4003 3617 4007
rect 3621 4003 3624 4007
rect 3574 3962 3577 3968
rect 3598 3952 3601 3958
rect 3630 3952 3633 4018
rect 3662 3951 3665 3958
rect 3558 3902 3561 3918
rect 3566 3752 3569 3859
rect 3574 3832 3577 3948
rect 3670 3942 3673 4018
rect 3614 3872 3617 3938
rect 3574 3792 3577 3828
rect 3582 3761 3585 3838
rect 3578 3758 3585 3761
rect 3598 3832 3601 3858
rect 3638 3842 3641 3858
rect 3654 3842 3657 3848
rect 3526 3732 3529 3738
rect 3558 3732 3561 3748
rect 3526 3692 3529 3718
rect 3534 3672 3537 3708
rect 3506 3668 3510 3671
rect 3442 3658 3446 3661
rect 3454 3652 3457 3658
rect 3394 3618 3401 3621
rect 3422 3618 3433 3621
rect 3350 3592 3353 3608
rect 3390 3552 3393 3608
rect 3398 3572 3401 3618
rect 3430 3592 3433 3618
rect 3406 3548 3414 3551
rect 3270 3462 3273 3468
rect 3154 3458 3158 3461
rect 3194 3458 3198 3461
rect 3234 3458 3238 3461
rect 3206 3451 3209 3458
rect 3202 3448 3209 3451
rect 3174 3432 3177 3438
rect 3246 3412 3249 3458
rect 3254 3452 3257 3458
rect 3262 3422 3265 3458
rect 3286 3452 3289 3488
rect 3294 3462 3297 3488
rect 3146 3338 3150 3341
rect 3146 3318 3150 3321
rect 3146 3278 3150 3281
rect 3126 3262 3129 3268
rect 3134 3262 3137 3268
rect 3106 3258 3110 3261
rect 3094 3192 3097 3258
rect 3098 3178 3102 3181
rect 3046 3162 3049 3178
rect 3070 3152 3073 3168
rect 3154 3148 3158 3151
rect 3062 3142 3065 3148
rect 3026 3138 3030 3141
rect 3014 3128 3025 3131
rect 2894 3058 2902 3061
rect 2886 3042 2889 3048
rect 2894 3031 2897 3058
rect 2918 3052 2921 3058
rect 2950 3052 2953 3059
rect 2902 3042 2905 3048
rect 2886 3028 2897 3031
rect 2870 2902 2873 2938
rect 2886 2872 2889 3028
rect 2934 2962 2937 3008
rect 2894 2952 2897 2958
rect 2918 2942 2921 2958
rect 2958 2952 2961 2998
rect 2982 2962 2985 3058
rect 2998 2952 3001 3128
rect 3014 3102 3017 3118
rect 3022 3092 3025 3128
rect 3058 3088 3062 3091
rect 3014 3062 3017 3088
rect 3046 3072 3049 3078
rect 3034 3068 3038 3071
rect 3022 3052 3025 3058
rect 3062 3052 3065 3078
rect 3070 3062 3073 3098
rect 3078 3092 3081 3138
rect 3096 3103 3098 3107
rect 3102 3103 3105 3107
rect 3109 3103 3112 3107
rect 3134 3062 3137 3118
rect 3142 3062 3145 3068
rect 3166 3062 3169 3378
rect 3278 3372 3281 3418
rect 3302 3392 3305 3538
rect 3318 3462 3321 3528
rect 3350 3462 3353 3518
rect 3358 3472 3361 3538
rect 3366 3492 3369 3528
rect 3342 3452 3345 3458
rect 3318 3392 3321 3448
rect 3358 3442 3361 3458
rect 3374 3432 3377 3478
rect 3382 3462 3385 3538
rect 3398 3452 3401 3518
rect 3406 3482 3409 3548
rect 3414 3532 3417 3538
rect 3422 3512 3425 3538
rect 3430 3482 3433 3528
rect 3438 3492 3441 3558
rect 3454 3552 3457 3558
rect 3470 3542 3473 3658
rect 3478 3562 3481 3618
rect 3502 3612 3505 3668
rect 3514 3658 3518 3661
rect 3494 3562 3497 3568
rect 3526 3552 3529 3558
rect 3478 3542 3481 3548
rect 3510 3542 3513 3548
rect 3446 3482 3449 3518
rect 3454 3472 3457 3478
rect 3406 3452 3409 3458
rect 3310 3372 3313 3378
rect 3282 3358 3286 3361
rect 3318 3352 3321 3388
rect 3326 3362 3329 3368
rect 3182 3263 3185 3268
rect 3206 3262 3209 3348
rect 3222 3332 3225 3348
rect 3262 3342 3265 3348
rect 3270 3322 3273 3348
rect 3270 3292 3273 3318
rect 3214 3272 3217 3278
rect 3210 3258 3214 3261
rect 3198 3142 3201 3208
rect 3214 3162 3217 3198
rect 3214 3152 3217 3158
rect 3182 3132 3185 3138
rect 3214 3062 3217 3068
rect 3090 3058 3094 3061
rect 3102 3042 3105 3058
rect 3110 3052 3113 3058
rect 3134 3002 3137 3058
rect 2950 2942 2953 2948
rect 2974 2942 2977 2948
rect 2994 2938 2998 2941
rect 2842 2868 2846 2871
rect 2782 2862 2785 2868
rect 2790 2862 2793 2868
rect 2750 2842 2753 2859
rect 2814 2852 2817 2868
rect 2794 2838 2798 2841
rect 2762 2768 2766 2771
rect 2798 2762 2801 2768
rect 2778 2758 2782 2761
rect 2814 2752 2817 2828
rect 2830 2792 2833 2868
rect 2842 2858 2846 2861
rect 2762 2738 2766 2741
rect 2774 2732 2777 2748
rect 2822 2742 2825 2788
rect 2830 2762 2833 2768
rect 2838 2751 2841 2838
rect 2846 2762 2849 2818
rect 2838 2748 2846 2751
rect 2854 2742 2857 2868
rect 2886 2862 2889 2868
rect 2846 2732 2849 2738
rect 2854 2732 2857 2738
rect 2726 2662 2729 2668
rect 2766 2662 2769 2718
rect 2822 2692 2825 2698
rect 2790 2652 2793 2658
rect 2622 2592 2625 2618
rect 2646 2572 2649 2618
rect 2654 2572 2657 2598
rect 2634 2558 2638 2561
rect 2662 2552 2665 2588
rect 2694 2552 2697 2558
rect 2702 2552 2705 2588
rect 2622 2452 2625 2538
rect 2630 2532 2633 2548
rect 2654 2532 2657 2538
rect 2630 2432 2633 2528
rect 2642 2478 2649 2481
rect 2646 2472 2649 2478
rect 2638 2462 2641 2468
rect 2646 2451 2649 2458
rect 2642 2448 2649 2451
rect 2654 2402 2657 2488
rect 2662 2391 2665 2538
rect 2686 2522 2689 2538
rect 2678 2492 2681 2518
rect 2694 2502 2697 2538
rect 2702 2502 2705 2548
rect 2710 2512 2713 2518
rect 2706 2468 2710 2471
rect 2686 2462 2689 2468
rect 2706 2458 2710 2461
rect 2694 2452 2697 2458
rect 2654 2388 2665 2391
rect 2702 2418 2710 2421
rect 2550 2362 2553 2368
rect 2586 2348 2590 2351
rect 2618 2348 2622 2351
rect 2502 2342 2505 2348
rect 2518 2342 2521 2348
rect 2486 2272 2489 2318
rect 2502 2292 2505 2328
rect 2510 2262 2513 2318
rect 2518 2272 2521 2338
rect 2534 2332 2537 2338
rect 2542 2262 2545 2348
rect 2570 2338 2574 2341
rect 2550 2282 2553 2318
rect 2566 2272 2569 2278
rect 2534 2252 2537 2258
rect 2470 2172 2473 2218
rect 2502 2212 2505 2248
rect 2478 2152 2481 2188
rect 2510 2162 2513 2188
rect 2498 2148 2502 2151
rect 2482 2138 2486 2141
rect 2398 2062 2401 2088
rect 2422 2072 2425 2088
rect 2502 2082 2505 2108
rect 2518 2092 2521 2208
rect 2526 2142 2529 2158
rect 2534 2142 2537 2218
rect 2542 2152 2545 2258
rect 2554 2248 2561 2251
rect 2534 2131 2537 2138
rect 2530 2128 2537 2131
rect 2434 2078 2438 2081
rect 2462 2062 2465 2068
rect 2442 2058 2449 2061
rect 2354 1947 2358 1950
rect 2390 1932 2393 1938
rect 2270 1902 2273 1918
rect 2358 1882 2361 1928
rect 2378 1888 2382 1891
rect 2230 1872 2233 1878
rect 2294 1862 2297 1878
rect 2398 1872 2401 2018
rect 2406 1952 2409 2028
rect 2438 1952 2441 2038
rect 2406 1942 2409 1948
rect 2414 1942 2417 1948
rect 2438 1942 2441 1948
rect 2426 1938 2430 1941
rect 2350 1862 2353 1868
rect 2406 1862 2409 1868
rect 2414 1862 2417 1918
rect 2422 1872 2425 1938
rect 2430 1892 2433 1928
rect 2438 1872 2441 1888
rect 2274 1858 2278 1861
rect 2362 1858 2366 1861
rect 2382 1852 2385 1858
rect 2430 1842 2433 1848
rect 2222 1752 2225 1808
rect 2246 1792 2249 1838
rect 2310 1772 2313 1838
rect 2446 1792 2449 2058
rect 2486 2052 2489 2068
rect 2510 2062 2513 2078
rect 2534 2072 2537 2108
rect 2558 2092 2561 2248
rect 2594 2218 2598 2221
rect 2606 2212 2609 2238
rect 2584 2203 2586 2207
rect 2590 2203 2593 2207
rect 2597 2203 2600 2207
rect 2590 2182 2593 2188
rect 2542 2072 2545 2088
rect 2454 1932 2457 1948
rect 2454 1852 2457 1858
rect 2462 1772 2465 1988
rect 2478 1952 2481 1958
rect 2486 1952 2489 2028
rect 2518 1992 2521 2068
rect 2550 2062 2553 2078
rect 2590 2072 2593 2108
rect 2582 2062 2585 2068
rect 2614 2062 2617 2338
rect 2630 2292 2633 2308
rect 2626 2148 2630 2151
rect 2638 2141 2641 2318
rect 2646 2262 2649 2378
rect 2654 2272 2657 2388
rect 2670 2351 2673 2418
rect 2678 2392 2681 2418
rect 2694 2352 2697 2368
rect 2666 2348 2673 2351
rect 2678 2272 2681 2308
rect 2678 2262 2681 2268
rect 2646 2252 2649 2258
rect 2646 2152 2649 2248
rect 2638 2138 2649 2141
rect 2542 2012 2545 2058
rect 2584 2003 2586 2007
rect 2590 2003 2593 2007
rect 2597 2003 2600 2007
rect 2494 1952 2497 1958
rect 2502 1952 2505 1968
rect 2562 1958 2566 1961
rect 2526 1942 2529 1948
rect 2542 1941 2545 1958
rect 2582 1942 2585 1948
rect 2542 1938 2553 1941
rect 2562 1938 2566 1941
rect 2470 1932 2473 1938
rect 2494 1892 2497 1898
rect 2478 1842 2481 1848
rect 2486 1842 2489 1858
rect 2262 1752 2265 1758
rect 2310 1752 2313 1768
rect 2414 1762 2417 1768
rect 2234 1748 2238 1751
rect 2226 1738 2230 1741
rect 2162 1688 2166 1691
rect 2174 1672 2177 1688
rect 2166 1658 2174 1661
rect 2150 1642 2153 1648
rect 2158 1642 2161 1648
rect 2142 1628 2153 1631
rect 2078 1552 2081 1578
rect 2090 1548 2094 1551
rect 2072 1503 2074 1507
rect 2078 1503 2081 1507
rect 2085 1503 2088 1507
rect 2102 1472 2105 1578
rect 2110 1552 2113 1558
rect 2110 1472 2113 1518
rect 2118 1502 2121 1618
rect 2142 1562 2145 1618
rect 2150 1602 2153 1628
rect 2150 1552 2153 1578
rect 2130 1528 2134 1531
rect 2142 1522 2145 1548
rect 2158 1532 2161 1548
rect 2158 1492 2161 1518
rect 2122 1488 2126 1491
rect 2166 1482 2169 1658
rect 2182 1592 2185 1678
rect 2190 1561 2193 1718
rect 2198 1682 2201 1728
rect 2278 1722 2281 1728
rect 2210 1718 2214 1721
rect 2318 1692 2321 1748
rect 2374 1732 2377 1758
rect 2390 1742 2393 1748
rect 2218 1688 2222 1691
rect 2242 1678 2246 1681
rect 2222 1662 2225 1668
rect 2230 1592 2233 1658
rect 2186 1558 2193 1561
rect 2222 1558 2249 1561
rect 2154 1468 2158 1471
rect 2038 1392 2041 1408
rect 2086 1372 2089 1468
rect 2094 1452 2097 1468
rect 2102 1452 2105 1458
rect 2126 1452 2129 1468
rect 2118 1442 2121 1448
rect 2142 1442 2145 1448
rect 2062 1352 2065 1358
rect 2070 1352 2073 1368
rect 2030 1292 2033 1348
rect 2054 1292 2057 1348
rect 2086 1332 2089 1358
rect 2072 1303 2074 1307
rect 2078 1303 2081 1307
rect 2085 1303 2088 1307
rect 2094 1292 2097 1308
rect 2102 1292 2105 1418
rect 2110 1352 2113 1358
rect 2126 1342 2129 1368
rect 2110 1321 2113 1338
rect 2110 1318 2121 1321
rect 2026 1268 2030 1271
rect 1974 1262 1977 1268
rect 1982 1262 1985 1268
rect 2046 1262 2049 1288
rect 1966 1248 1977 1251
rect 1866 1068 1873 1071
rect 1882 1068 1886 1071
rect 1898 1068 1902 1071
rect 1854 1032 1857 1058
rect 1838 842 1841 888
rect 1854 812 1857 1028
rect 1862 992 1865 1048
rect 1870 902 1873 1068
rect 1910 1062 1913 1068
rect 1918 1062 1921 1068
rect 1930 1048 1934 1051
rect 1870 882 1873 898
rect 1878 871 1881 1048
rect 1902 1042 1905 1048
rect 1870 868 1881 871
rect 1862 752 1865 798
rect 1858 568 1862 571
rect 1870 571 1873 868
rect 1894 852 1897 858
rect 1878 742 1881 818
rect 1894 792 1897 848
rect 1894 662 1897 698
rect 1902 672 1905 968
rect 1914 948 1918 951
rect 1942 942 1945 988
rect 1958 942 1961 1078
rect 1966 992 1969 1148
rect 1974 1112 1977 1248
rect 1982 1062 1985 1138
rect 1990 1132 1993 1148
rect 1998 1142 2001 1248
rect 2006 1222 2009 1248
rect 2002 1088 2006 1091
rect 2022 1072 2025 1078
rect 2030 1062 2033 1188
rect 2038 1132 2041 1138
rect 2046 1121 2049 1238
rect 2054 1212 2057 1268
rect 2054 1152 2057 1158
rect 2038 1118 2049 1121
rect 2018 1058 2022 1061
rect 1974 1012 1977 1058
rect 1982 1032 1985 1058
rect 2030 1042 2033 1048
rect 1982 972 1985 978
rect 2002 958 2006 961
rect 1910 892 1913 908
rect 1918 872 1921 938
rect 1958 892 1961 938
rect 1966 912 1969 948
rect 2014 942 2017 968
rect 2022 952 2025 998
rect 2038 992 2041 1118
rect 2062 1092 2065 1248
rect 2078 1242 2081 1268
rect 2090 1258 2094 1261
rect 2098 1248 2102 1251
rect 2110 1232 2113 1258
rect 2118 1202 2121 1318
rect 2126 1292 2129 1298
rect 2142 1292 2145 1328
rect 2150 1302 2153 1458
rect 2162 1448 2169 1451
rect 2158 1342 2161 1348
rect 2166 1292 2169 1448
rect 2174 1362 2177 1558
rect 2198 1552 2201 1558
rect 2222 1552 2225 1558
rect 2246 1552 2249 1558
rect 2234 1548 2238 1551
rect 2190 1522 2193 1548
rect 2206 1532 2209 1548
rect 2254 1542 2257 1658
rect 2262 1542 2265 1678
rect 2350 1672 2353 1678
rect 2270 1562 2273 1628
rect 2286 1582 2289 1588
rect 2214 1522 2217 1538
rect 2270 1532 2273 1558
rect 2282 1548 2286 1551
rect 2282 1538 2286 1541
rect 2194 1468 2198 1471
rect 2182 1442 2185 1468
rect 2190 1452 2193 1458
rect 2206 1452 2209 1498
rect 2214 1492 2217 1508
rect 2246 1472 2249 1478
rect 2254 1462 2257 1528
rect 2246 1452 2249 1458
rect 2218 1448 2225 1451
rect 2206 1442 2209 1448
rect 2158 1262 2161 1268
rect 2142 1242 2145 1248
rect 2126 1212 2129 1218
rect 2118 1162 2121 1168
rect 2106 1158 2110 1161
rect 2090 1148 2097 1151
rect 2074 1138 2078 1141
rect 2072 1103 2074 1107
rect 2078 1103 2081 1107
rect 2085 1103 2088 1107
rect 2046 1052 2049 1088
rect 2074 1068 2078 1071
rect 2094 1062 2097 1148
rect 2126 1151 2129 1208
rect 2158 1162 2161 1248
rect 2174 1162 2177 1338
rect 2182 1272 2185 1298
rect 2190 1272 2193 1418
rect 2198 1372 2201 1418
rect 2222 1372 2225 1448
rect 2214 1362 2217 1368
rect 2218 1348 2222 1351
rect 2210 1318 2214 1321
rect 2198 1292 2201 1318
rect 2214 1292 2217 1308
rect 2230 1292 2233 1438
rect 2238 1352 2241 1448
rect 2254 1422 2257 1458
rect 2262 1452 2265 1458
rect 2270 1452 2273 1518
rect 2282 1478 2286 1481
rect 2294 1442 2297 1578
rect 2302 1552 2305 1558
rect 2310 1442 2313 1668
rect 2318 1642 2321 1659
rect 2350 1652 2353 1658
rect 2374 1652 2377 1718
rect 2398 1692 2401 1758
rect 2430 1752 2433 1768
rect 2438 1752 2441 1758
rect 2462 1752 2465 1758
rect 2518 1752 2521 1778
rect 2542 1761 2545 1918
rect 2538 1758 2545 1761
rect 2550 1782 2553 1938
rect 2566 1852 2569 1858
rect 2550 1752 2553 1778
rect 2574 1761 2577 1918
rect 2590 1872 2593 1878
rect 2584 1803 2586 1807
rect 2590 1803 2593 1807
rect 2597 1803 2600 1807
rect 2570 1758 2577 1761
rect 2558 1752 2561 1758
rect 2410 1748 2414 1751
rect 2490 1748 2494 1751
rect 2570 1748 2574 1751
rect 2470 1741 2473 1748
rect 2462 1738 2473 1741
rect 2478 1742 2481 1748
rect 2502 1742 2505 1748
rect 2542 1742 2545 1748
rect 2422 1732 2425 1738
rect 2418 1718 2425 1721
rect 2422 1692 2425 1718
rect 2430 1692 2433 1728
rect 2462 1692 2465 1738
rect 2510 1732 2513 1738
rect 2474 1688 2478 1691
rect 2438 1682 2441 1688
rect 2406 1672 2409 1678
rect 2386 1668 2390 1671
rect 2450 1668 2454 1671
rect 2318 1592 2321 1608
rect 2342 1552 2345 1598
rect 2334 1542 2337 1548
rect 2342 1542 2345 1548
rect 2318 1502 2321 1518
rect 2334 1452 2337 1458
rect 2286 1362 2289 1408
rect 2298 1358 2302 1361
rect 2314 1358 2318 1361
rect 2330 1358 2334 1361
rect 2342 1352 2345 1478
rect 2350 1422 2353 1648
rect 2362 1638 2366 1641
rect 2398 1612 2401 1648
rect 2422 1642 2425 1648
rect 2430 1642 2433 1658
rect 2410 1588 2414 1591
rect 2358 1542 2361 1548
rect 2358 1522 2361 1538
rect 2358 1412 2361 1468
rect 2242 1348 2246 1351
rect 2322 1348 2326 1351
rect 2270 1342 2273 1348
rect 2350 1342 2353 1348
rect 2322 1338 2326 1341
rect 2246 1322 2249 1328
rect 2326 1322 2329 1328
rect 2286 1292 2289 1318
rect 2182 1182 2185 1268
rect 2190 1192 2193 1268
rect 2230 1262 2233 1288
rect 2310 1272 2313 1288
rect 2238 1251 2241 1268
rect 2246 1262 2249 1268
rect 2270 1262 2273 1268
rect 2218 1248 2225 1251
rect 2238 1248 2249 1251
rect 2206 1242 2209 1248
rect 2122 1148 2129 1151
rect 2174 1152 2177 1158
rect 2102 1142 2105 1148
rect 2190 1142 2193 1148
rect 2110 1131 2113 1138
rect 2102 1128 2113 1131
rect 2102 1082 2105 1128
rect 2118 1072 2121 1098
rect 2090 1048 2094 1051
rect 2054 982 2057 1048
rect 2110 1042 2113 1048
rect 2118 1002 2121 1058
rect 2150 1052 2153 1059
rect 2050 978 2054 981
rect 2150 962 2153 1028
rect 2110 952 2113 958
rect 2022 941 2025 948
rect 2022 938 2033 941
rect 2022 912 2025 928
rect 1958 862 1961 878
rect 1966 872 1969 908
rect 1974 752 1977 858
rect 2006 792 2009 908
rect 2022 872 2025 898
rect 2014 842 2017 848
rect 2022 792 2025 868
rect 2030 862 2033 938
rect 2072 903 2074 907
rect 2078 903 2081 907
rect 2085 903 2088 907
rect 2038 872 2041 878
rect 2078 872 2081 888
rect 2070 862 2073 868
rect 2030 752 2033 858
rect 2054 842 2057 848
rect 2070 752 2073 788
rect 2078 752 2081 808
rect 2094 792 2097 938
rect 2106 888 2110 891
rect 2126 872 2129 908
rect 2134 892 2137 938
rect 2150 891 2153 958
rect 2146 888 2153 891
rect 2158 881 2161 1068
rect 2170 958 2174 961
rect 2178 958 2182 961
rect 2198 952 2201 1218
rect 2222 1092 2225 1248
rect 2238 1192 2241 1198
rect 2246 1181 2249 1248
rect 2254 1222 2257 1258
rect 2278 1252 2281 1268
rect 2270 1192 2273 1248
rect 2294 1212 2297 1258
rect 2302 1252 2305 1268
rect 2238 1178 2249 1181
rect 2238 1102 2241 1178
rect 2258 1148 2262 1151
rect 2278 1142 2281 1148
rect 2246 1112 2249 1128
rect 2286 1112 2289 1118
rect 2270 1092 2273 1108
rect 2302 1102 2305 1118
rect 2210 1088 2214 1091
rect 2234 1068 2238 1071
rect 2250 1068 2254 1071
rect 2258 1058 2262 1061
rect 2218 1048 2222 1051
rect 2194 948 2198 951
rect 2166 912 2169 948
rect 2206 942 2209 998
rect 2222 992 2225 1028
rect 2246 992 2249 1058
rect 2270 1052 2273 1088
rect 2302 1072 2305 1098
rect 2318 1072 2321 1158
rect 2342 1152 2345 1158
rect 2350 1142 2353 1268
rect 2362 1258 2366 1261
rect 2374 1172 2377 1538
rect 2390 1492 2393 1588
rect 2398 1522 2401 1548
rect 2406 1512 2409 1548
rect 2422 1532 2425 1608
rect 2406 1472 2409 1508
rect 2414 1462 2417 1518
rect 2422 1502 2425 1528
rect 2454 1522 2457 1548
rect 2430 1492 2433 1508
rect 2438 1491 2441 1518
rect 2454 1492 2457 1498
rect 2438 1488 2446 1491
rect 2422 1482 2425 1488
rect 2462 1472 2465 1648
rect 2486 1522 2489 1548
rect 2434 1468 2438 1471
rect 2398 1402 2401 1418
rect 2414 1362 2417 1418
rect 2390 1272 2393 1328
rect 2414 1292 2417 1358
rect 2438 1352 2441 1468
rect 2450 1458 2454 1461
rect 2470 1392 2473 1518
rect 2502 1482 2505 1678
rect 2534 1663 2537 1718
rect 2550 1672 2553 1688
rect 2526 1552 2529 1558
rect 2550 1552 2553 1668
rect 2566 1652 2569 1658
rect 2586 1618 2590 1621
rect 2584 1603 2586 1607
rect 2590 1603 2593 1607
rect 2597 1603 2600 1607
rect 2510 1462 2513 1508
rect 2518 1482 2521 1528
rect 2550 1462 2553 1518
rect 2566 1492 2569 1588
rect 2486 1412 2489 1458
rect 2606 1432 2609 2038
rect 2614 1932 2617 2058
rect 2622 1982 2625 1998
rect 2614 1862 2617 1918
rect 2622 1872 2625 1968
rect 2630 1872 2633 2068
rect 2638 1972 2641 2118
rect 2646 2002 2649 2138
rect 2654 2012 2657 2058
rect 2662 1992 2665 2218
rect 2670 2122 2673 2128
rect 2686 1992 2689 2348
rect 2694 2292 2697 2298
rect 2702 2282 2705 2418
rect 2718 2411 2721 2648
rect 2742 2562 2745 2628
rect 2774 2562 2777 2568
rect 2790 2562 2793 2588
rect 2806 2561 2809 2668
rect 2822 2652 2825 2688
rect 2830 2662 2833 2668
rect 2838 2651 2841 2718
rect 2834 2648 2841 2651
rect 2846 2662 2849 2708
rect 2870 2702 2873 2838
rect 2886 2832 2889 2858
rect 2894 2812 2897 2868
rect 2902 2862 2905 2908
rect 2918 2862 2921 2868
rect 2942 2862 2945 2888
rect 2894 2762 2897 2768
rect 2882 2758 2886 2761
rect 2878 2742 2881 2748
rect 2878 2722 2881 2728
rect 2854 2672 2857 2678
rect 2866 2668 2870 2671
rect 2886 2662 2889 2738
rect 2902 2672 2905 2778
rect 2934 2682 2937 2728
rect 2950 2692 2953 2918
rect 2986 2868 2990 2871
rect 2966 2862 2969 2868
rect 3022 2862 3025 2988
rect 3030 2892 3033 2898
rect 3038 2862 3041 2878
rect 3046 2862 3049 2978
rect 3130 2958 3134 2961
rect 3054 2942 3057 2958
rect 3070 2951 3073 2958
rect 3122 2948 3126 2951
rect 3106 2938 3110 2941
rect 3142 2941 3145 3048
rect 3150 2952 3153 2958
rect 3142 2938 3153 2941
rect 3054 2872 3057 2938
rect 3066 2888 3070 2891
rect 3078 2882 3081 2908
rect 3096 2903 3098 2907
rect 3102 2903 3105 2907
rect 3109 2903 3112 2907
rect 2986 2858 2990 2861
rect 2918 2672 2921 2678
rect 2894 2662 2897 2668
rect 2846 2572 2849 2658
rect 2862 2652 2865 2658
rect 2910 2652 2913 2658
rect 2890 2648 2894 2651
rect 2798 2558 2809 2561
rect 2758 2552 2761 2558
rect 2798 2552 2801 2558
rect 2814 2552 2817 2558
rect 2830 2552 2833 2558
rect 2746 2548 2750 2551
rect 2778 2548 2782 2551
rect 2850 2548 2854 2551
rect 2822 2542 2825 2548
rect 2726 2522 2729 2538
rect 2758 2532 2761 2538
rect 2726 2472 2729 2518
rect 2734 2462 2737 2478
rect 2742 2472 2745 2498
rect 2742 2462 2745 2468
rect 2710 2408 2721 2411
rect 2710 2392 2713 2408
rect 2750 2392 2753 2528
rect 2782 2512 2785 2518
rect 2794 2478 2798 2481
rect 2758 2458 2766 2461
rect 2758 2442 2761 2458
rect 2774 2452 2777 2458
rect 2782 2452 2785 2458
rect 2766 2448 2774 2451
rect 2706 2258 2710 2261
rect 2718 2152 2721 2288
rect 2726 2272 2729 2348
rect 2734 2292 2737 2378
rect 2766 2352 2769 2448
rect 2806 2422 2809 2538
rect 2838 2522 2841 2528
rect 2850 2518 2854 2521
rect 2814 2462 2817 2468
rect 2862 2461 2865 2598
rect 2870 2592 2873 2618
rect 2886 2462 2889 2568
rect 2894 2472 2897 2548
rect 2910 2532 2913 2548
rect 2918 2522 2921 2668
rect 2930 2658 2934 2661
rect 2958 2592 2961 2818
rect 2966 2732 2969 2748
rect 2974 2692 2977 2858
rect 3014 2852 3017 2858
rect 3018 2738 3022 2741
rect 2998 2732 3001 2738
rect 2998 2682 3001 2728
rect 3030 2661 3033 2788
rect 3046 2772 3049 2858
rect 3054 2742 3057 2868
rect 3142 2862 3145 2868
rect 3074 2848 3078 2851
rect 3086 2781 3089 2818
rect 3094 2792 3097 2848
rect 3110 2842 3113 2858
rect 3086 2778 3097 2781
rect 3086 2762 3089 2768
rect 3082 2738 3086 2741
rect 3094 2721 3097 2778
rect 3142 2762 3145 2778
rect 3086 2718 3097 2721
rect 3062 2692 3065 2698
rect 3070 2672 3073 2678
rect 3086 2672 3089 2718
rect 3118 2712 3121 2738
rect 3126 2732 3129 2738
rect 3096 2703 3098 2707
rect 3102 2703 3105 2707
rect 3109 2703 3112 2707
rect 3150 2692 3153 2938
rect 3130 2678 3134 2681
rect 3110 2662 3113 2668
rect 3026 2658 3033 2661
rect 2966 2612 2969 2658
rect 2982 2562 2985 2608
rect 2934 2542 2937 2558
rect 2962 2548 2966 2551
rect 2950 2542 2953 2548
rect 2974 2541 2977 2548
rect 2982 2541 2985 2558
rect 2974 2538 2985 2541
rect 2998 2542 3001 2658
rect 3086 2652 3089 2658
rect 3110 2622 3113 2658
rect 3158 2642 3161 3018
rect 3214 2952 3217 2978
rect 3186 2938 3190 2941
rect 3166 2902 3169 2938
rect 3174 2922 3177 2938
rect 3198 2932 3201 2948
rect 3166 2862 3169 2888
rect 3190 2792 3193 2888
rect 3206 2872 3209 2888
rect 3210 2858 3214 2861
rect 3222 2861 3225 3188
rect 3242 3178 3246 3181
rect 3254 3171 3257 3278
rect 3310 3272 3313 3338
rect 3318 3302 3321 3338
rect 3334 3302 3337 3418
rect 3382 3382 3385 3448
rect 3398 3412 3401 3418
rect 3414 3372 3417 3468
rect 3430 3462 3433 3468
rect 3438 3442 3441 3448
rect 3454 3442 3457 3458
rect 3422 3392 3425 3428
rect 3374 3352 3377 3368
rect 3358 3342 3361 3348
rect 3398 3308 3406 3311
rect 3370 3288 3374 3291
rect 3266 3268 3270 3271
rect 3310 3262 3313 3268
rect 3322 3258 3326 3261
rect 3270 3252 3273 3258
rect 3254 3168 3265 3171
rect 3234 3148 3238 3151
rect 3246 3142 3249 3148
rect 3238 3062 3241 3128
rect 3238 2942 3241 2978
rect 3246 2952 3249 2968
rect 3262 2952 3265 3168
rect 3278 3151 3281 3178
rect 3286 3092 3289 3138
rect 3294 3132 3297 3138
rect 3310 3122 3313 3258
rect 3334 3092 3337 3228
rect 3314 3068 3318 3071
rect 3330 3068 3334 3071
rect 3342 3062 3345 3198
rect 3350 3162 3353 3278
rect 3398 3272 3401 3308
rect 3406 3282 3409 3288
rect 3422 3272 3425 3278
rect 3374 3262 3377 3268
rect 3438 3262 3441 3438
rect 3462 3432 3465 3438
rect 3454 3342 3457 3348
rect 3394 3258 3398 3261
rect 3458 3258 3462 3261
rect 3374 3232 3377 3248
rect 3390 3202 3393 3258
rect 3390 3162 3393 3178
rect 3350 3152 3353 3158
rect 3398 3152 3401 3218
rect 3370 3148 3374 3151
rect 3398 3142 3401 3148
rect 3362 3138 3366 3141
rect 3354 3088 3358 3091
rect 3350 3082 3353 3088
rect 3306 3058 3310 3061
rect 3342 3052 3345 3058
rect 3310 3048 3318 3051
rect 3234 2918 3238 2921
rect 3222 2858 3230 2861
rect 3210 2848 3214 2851
rect 3170 2788 3174 2791
rect 3166 2752 3169 2778
rect 3222 2772 3225 2858
rect 3238 2851 3241 2888
rect 3254 2881 3257 2948
rect 3234 2848 3241 2851
rect 3246 2878 3257 2881
rect 3246 2832 3249 2878
rect 3262 2872 3265 2938
rect 3270 2862 3273 2998
rect 3286 2952 3289 2958
rect 3278 2862 3281 2918
rect 3310 2872 3313 3048
rect 3342 2972 3345 3048
rect 3326 2942 3329 2947
rect 3222 2752 3225 2768
rect 3254 2752 3257 2828
rect 3262 2752 3265 2768
rect 3250 2748 3254 2751
rect 3182 2702 3185 2728
rect 3198 2682 3201 2708
rect 3166 2652 3169 2658
rect 3138 2628 3142 2631
rect 3078 2602 3081 2618
rect 3006 2542 3009 2548
rect 2966 2532 2969 2538
rect 2902 2472 2905 2498
rect 2862 2458 2873 2461
rect 2782 2392 2785 2408
rect 2798 2352 2801 2408
rect 2822 2382 2825 2458
rect 2830 2452 2833 2458
rect 2870 2452 2873 2458
rect 2918 2452 2921 2508
rect 2950 2481 2953 2498
rect 2950 2478 2961 2481
rect 2958 2472 2961 2478
rect 2950 2462 2953 2468
rect 2966 2462 2969 2488
rect 2838 2412 2841 2418
rect 2734 2172 2737 2218
rect 2702 2052 2705 2118
rect 2734 2112 2737 2118
rect 2710 2082 2713 2088
rect 2734 2082 2737 2108
rect 2714 2068 2718 2071
rect 2734 2052 2737 2058
rect 2730 2038 2737 2041
rect 2734 1992 2737 2038
rect 2638 1952 2641 1968
rect 2646 1952 2649 1978
rect 2666 1958 2670 1961
rect 2718 1952 2721 1968
rect 2638 1902 2641 1938
rect 2646 1912 2649 1948
rect 2702 1942 2705 1948
rect 2710 1922 2713 1948
rect 2702 1872 2705 1878
rect 2682 1868 2686 1871
rect 2614 1832 2617 1858
rect 2622 1772 2625 1868
rect 2726 1862 2729 1928
rect 2718 1762 2721 1828
rect 2734 1782 2737 1918
rect 2742 1792 2745 2348
rect 2774 2342 2777 2348
rect 2750 2302 2753 2318
rect 2750 2252 2753 2258
rect 2758 2182 2761 2308
rect 2790 2292 2793 2328
rect 2814 2272 2817 2358
rect 2822 2352 2825 2358
rect 2882 2348 2886 2351
rect 2770 2268 2774 2271
rect 2766 2262 2769 2268
rect 2806 2262 2809 2268
rect 2822 2262 2825 2298
rect 2838 2252 2841 2348
rect 2854 2312 2857 2338
rect 2854 2262 2857 2278
rect 2846 2242 2849 2258
rect 2790 2202 2793 2218
rect 2758 2142 2761 2178
rect 2766 2072 2769 2088
rect 2762 2058 2766 2061
rect 2774 2052 2777 2158
rect 2786 2148 2790 2151
rect 2790 2072 2793 2078
rect 2798 2072 2801 2228
rect 2862 2142 2865 2308
rect 2886 2292 2889 2338
rect 2902 2282 2905 2428
rect 2926 2392 2929 2458
rect 2934 2452 2937 2458
rect 2974 2362 2977 2538
rect 2982 2452 2985 2498
rect 3014 2472 3017 2578
rect 3022 2532 3025 2538
rect 3014 2462 3017 2468
rect 3030 2462 3033 2588
rect 3086 2562 3089 2568
rect 3174 2552 3177 2608
rect 3198 2562 3201 2608
rect 3130 2547 3134 2550
rect 3186 2548 3190 2551
rect 3150 2532 3153 2538
rect 3166 2522 3169 2538
rect 3042 2518 3046 2521
rect 3046 2492 3049 2498
rect 3086 2492 3089 2508
rect 3096 2503 3098 2507
rect 3102 2503 3105 2507
rect 3109 2503 3112 2507
rect 3058 2468 3062 2471
rect 3038 2462 3041 2468
rect 3070 2462 3073 2488
rect 3158 2472 3161 2498
rect 3182 2492 3185 2518
rect 3198 2502 3201 2558
rect 3206 2492 3209 2718
rect 3214 2662 3217 2698
rect 3270 2582 3273 2858
rect 3278 2792 3281 2838
rect 3310 2832 3313 2858
rect 3318 2852 3321 2878
rect 3326 2872 3329 2928
rect 3342 2882 3345 2968
rect 3354 2888 3358 2891
rect 3334 2862 3337 2868
rect 3342 2862 3345 2868
rect 3358 2852 3361 2878
rect 3382 2861 3385 3138
rect 3398 3062 3401 3138
rect 3414 3132 3417 3148
rect 3406 3072 3409 3128
rect 3422 3121 3425 3258
rect 3470 3252 3473 3538
rect 3518 3462 3521 3538
rect 3534 3532 3537 3648
rect 3542 3532 3545 3718
rect 3574 3692 3577 3748
rect 3598 3742 3601 3828
rect 3662 3812 3665 3888
rect 3686 3862 3689 4068
rect 3706 4058 3710 4061
rect 3694 3892 3697 3918
rect 3608 3803 3610 3807
rect 3614 3803 3617 3807
rect 3621 3803 3624 3807
rect 3642 3768 3646 3771
rect 3686 3762 3689 3768
rect 3674 3758 3678 3761
rect 3590 3712 3593 3718
rect 3606 3692 3609 3758
rect 3614 3742 3617 3748
rect 3670 3742 3673 3748
rect 3686 3742 3689 3758
rect 3630 3692 3633 3738
rect 3662 3732 3665 3738
rect 3654 3722 3657 3728
rect 3550 3662 3553 3688
rect 3566 3682 3569 3688
rect 3562 3668 3566 3671
rect 3534 3482 3537 3518
rect 3542 3462 3545 3478
rect 3478 3441 3481 3448
rect 3478 3438 3489 3441
rect 3478 3352 3481 3368
rect 3486 3292 3489 3438
rect 3518 3372 3521 3398
rect 3534 3342 3537 3428
rect 3566 3372 3569 3658
rect 3574 3652 3577 3688
rect 3630 3662 3633 3688
rect 3638 3672 3641 3698
rect 3582 3622 3585 3658
rect 3590 3641 3593 3658
rect 3590 3638 3598 3641
rect 3582 3602 3585 3618
rect 3646 3612 3649 3658
rect 3608 3603 3610 3607
rect 3614 3603 3617 3607
rect 3621 3603 3624 3607
rect 3654 3552 3657 3718
rect 3662 3652 3665 3688
rect 3686 3662 3689 3718
rect 3694 3712 3697 3818
rect 3702 3792 3705 3888
rect 3710 3872 3713 4058
rect 3742 4052 3745 4088
rect 3766 4062 3769 4068
rect 3758 4052 3761 4058
rect 3774 4052 3777 4118
rect 3798 4072 3801 4258
rect 3806 4252 3809 4278
rect 3814 4262 3817 4268
rect 3814 4222 3817 4248
rect 3822 4232 3825 4508
rect 3830 4382 3833 4548
rect 3870 4472 3873 4598
rect 3886 4532 3889 4548
rect 3878 4492 3881 4518
rect 3838 4442 3841 4448
rect 3830 4342 3833 4348
rect 3846 4272 3849 4428
rect 3854 4402 3857 4458
rect 3862 4452 3865 4458
rect 3854 4352 3857 4378
rect 3842 4268 3846 4271
rect 3830 4232 3833 4258
rect 3822 4142 3825 4228
rect 3830 4152 3833 4228
rect 3846 4212 3849 4258
rect 3854 4212 3857 4348
rect 3870 4282 3873 4468
rect 3878 4452 3881 4458
rect 3886 4332 3889 4458
rect 3894 4352 3897 4668
rect 3926 4662 3929 4738
rect 3994 4718 3998 4721
rect 4006 4682 4009 4698
rect 4006 4672 4009 4678
rect 3962 4668 3966 4671
rect 3926 4652 3929 4658
rect 3910 4622 3913 4648
rect 3926 4632 3929 4638
rect 3934 4622 3937 4668
rect 3942 4662 3945 4668
rect 3974 4662 3977 4668
rect 4010 4658 4014 4661
rect 3982 4652 3985 4658
rect 3942 4642 3945 4648
rect 3982 4622 3985 4648
rect 3902 4542 3905 4548
rect 3910 4492 3913 4558
rect 3926 4552 3929 4558
rect 3918 4532 3921 4538
rect 3934 4512 3937 4618
rect 3902 4472 3905 4488
rect 3942 4482 3945 4558
rect 3950 4472 3953 4518
rect 3966 4512 3969 4548
rect 3974 4542 3977 4608
rect 3982 4552 3985 4618
rect 3998 4541 4001 4658
rect 4030 4652 4033 4718
rect 4038 4692 4041 4748
rect 4070 4742 4073 4758
rect 4086 4692 4089 4758
rect 4094 4722 4097 4818
rect 4106 4778 4110 4781
rect 4158 4762 4161 4768
rect 4102 4711 4105 4748
rect 4110 4732 4113 4738
rect 4094 4708 4105 4711
rect 4078 4682 4081 4688
rect 4054 4652 4057 4658
rect 4014 4562 4017 4568
rect 4006 4552 4009 4558
rect 3998 4538 4009 4541
rect 3902 4452 3905 4458
rect 3910 4442 3913 4448
rect 3926 4412 3929 4468
rect 3966 4462 3969 4508
rect 3974 4502 3977 4538
rect 3982 4532 3985 4538
rect 3998 4462 4001 4468
rect 3914 4338 3918 4341
rect 3894 4322 3897 4338
rect 3886 4312 3889 4318
rect 3926 4312 3929 4358
rect 3866 4268 3870 4271
rect 3878 4262 3881 4268
rect 3850 4188 3854 4191
rect 3846 4152 3849 4158
rect 3814 4132 3817 4138
rect 3862 4092 3865 4258
rect 3878 4242 3881 4248
rect 3854 4062 3857 4068
rect 3794 4058 3798 4061
rect 3806 4052 3809 4058
rect 3790 4042 3793 4048
rect 3758 4032 3761 4038
rect 3814 4032 3817 4058
rect 3838 4042 3841 4058
rect 3722 3988 3726 3991
rect 3850 3978 3854 3981
rect 3850 3958 3854 3961
rect 3734 3912 3737 3918
rect 3750 3872 3753 3878
rect 3758 3862 3761 3908
rect 3766 3872 3769 3948
rect 3710 3801 3713 3858
rect 3718 3852 3721 3858
rect 3710 3798 3718 3801
rect 3710 3762 3713 3768
rect 3710 3752 3713 3758
rect 3718 3752 3721 3758
rect 3726 3752 3729 3858
rect 3750 3752 3753 3768
rect 3738 3748 3742 3751
rect 3746 3738 3753 3741
rect 3698 3688 3702 3691
rect 3694 3662 3697 3668
rect 3690 3638 3694 3641
rect 3602 3548 3606 3551
rect 3646 3548 3654 3551
rect 3630 3542 3633 3548
rect 3574 3492 3577 3508
rect 3582 3482 3585 3538
rect 3578 3468 3582 3471
rect 3626 3468 3630 3471
rect 3638 3462 3641 3478
rect 3638 3452 3641 3458
rect 3594 3448 3598 3451
rect 3608 3403 3610 3407
rect 3614 3403 3617 3407
rect 3621 3403 3624 3407
rect 3646 3402 3649 3548
rect 3662 3542 3665 3578
rect 3682 3538 3686 3541
rect 3694 3512 3697 3558
rect 3662 3482 3665 3488
rect 3670 3482 3673 3508
rect 3710 3502 3713 3718
rect 3718 3672 3721 3708
rect 3718 3542 3721 3668
rect 3734 3592 3737 3608
rect 3742 3552 3745 3658
rect 3750 3622 3753 3738
rect 3766 3702 3769 3868
rect 3774 3862 3777 3868
rect 3782 3832 3785 3938
rect 3790 3932 3793 3948
rect 3814 3942 3817 3948
rect 3830 3932 3833 3938
rect 3802 3888 3806 3891
rect 3782 3752 3785 3828
rect 3790 3802 3793 3848
rect 3814 3762 3817 3858
rect 3822 3852 3825 3868
rect 3838 3862 3841 3878
rect 3846 3832 3849 3918
rect 3870 3871 3873 4218
rect 3886 4082 3889 4308
rect 3910 4272 3913 4298
rect 3934 4292 3937 4458
rect 3942 4422 3945 4438
rect 3966 4382 3969 4438
rect 4006 4412 4009 4538
rect 4014 4532 4017 4558
rect 4030 4552 4033 4648
rect 4062 4582 4065 4668
rect 4086 4642 4089 4648
rect 4038 4531 4041 4548
rect 4030 4528 4041 4531
rect 4062 4532 4065 4538
rect 4014 4482 4017 4518
rect 4030 4482 4033 4528
rect 3974 4352 3977 4358
rect 3942 4342 3945 4348
rect 3954 4338 3958 4341
rect 3966 4332 3969 4348
rect 4014 4342 4017 4468
rect 4030 4382 4033 4478
rect 4054 4462 4057 4518
rect 4062 4482 4065 4488
rect 4046 4452 4049 4458
rect 4046 4372 4049 4418
rect 4030 4362 4033 4368
rect 4054 4352 4057 4408
rect 4054 4342 4057 4348
rect 3994 4338 3998 4341
rect 4026 4338 4030 4341
rect 3958 4292 3961 4318
rect 3974 4292 3977 4318
rect 4006 4312 4009 4338
rect 3990 4282 3993 4298
rect 3938 4268 3942 4271
rect 3898 4248 3902 4251
rect 3910 4232 3913 4268
rect 3918 4262 3921 4268
rect 3958 4252 3961 4268
rect 3930 4248 3934 4251
rect 3954 4248 3958 4251
rect 4014 4251 4017 4318
rect 4026 4268 4030 4271
rect 4010 4248 4017 4251
rect 4022 4252 4025 4258
rect 4038 4252 4041 4318
rect 3982 4242 3985 4248
rect 3894 4152 3897 4208
rect 3950 4182 3953 4218
rect 3998 4182 4001 4218
rect 3918 4151 3921 4168
rect 3966 4162 3969 4168
rect 3974 4162 3977 4178
rect 4002 4168 4006 4171
rect 3950 4152 3953 4158
rect 3974 4152 3977 4158
rect 3970 4138 3974 4141
rect 3982 4122 3985 4138
rect 3934 4062 3937 4088
rect 3950 4062 3953 4068
rect 3906 4058 3910 4061
rect 3878 3892 3881 3898
rect 3862 3868 3873 3871
rect 3862 3862 3865 3868
rect 3870 3832 3873 3858
rect 3782 3672 3785 3748
rect 3798 3682 3801 3748
rect 3810 3747 3814 3750
rect 3830 3692 3833 3748
rect 3854 3742 3857 3818
rect 3862 3742 3865 3828
rect 3870 3732 3873 3828
rect 3846 3722 3849 3728
rect 3854 3692 3857 3718
rect 3878 3712 3881 3738
rect 3758 3642 3761 3658
rect 3798 3602 3801 3678
rect 3834 3668 3838 3671
rect 3814 3662 3817 3668
rect 3846 3662 3849 3668
rect 3854 3662 3857 3678
rect 3886 3662 3889 4058
rect 3942 4032 3945 4058
rect 3894 3821 3897 4018
rect 3926 3992 3929 4018
rect 3918 3922 3921 3947
rect 3934 3942 3937 3948
rect 3950 3932 3953 3978
rect 3958 3932 3961 4118
rect 3974 4062 3977 4068
rect 3990 4051 3993 4118
rect 4006 4112 4009 4138
rect 4014 4082 4017 4228
rect 4010 4068 4014 4071
rect 3998 4062 4001 4068
rect 3986 4048 3993 4051
rect 4022 4042 4025 4218
rect 4030 4052 4033 4088
rect 4046 4071 4049 4288
rect 4062 4272 4065 4398
rect 4070 4292 4073 4618
rect 4078 4572 4081 4628
rect 4094 4602 4097 4708
rect 4112 4703 4114 4707
rect 4118 4703 4121 4707
rect 4125 4703 4128 4707
rect 4134 4682 4137 4738
rect 4142 4701 4145 4748
rect 4142 4698 4150 4701
rect 4110 4672 4113 4678
rect 4150 4662 4153 4698
rect 4158 4692 4161 4758
rect 4166 4742 4169 4808
rect 4182 4752 4185 4858
rect 4222 4822 4225 4878
rect 4238 4872 4241 4878
rect 4362 4868 4366 4871
rect 4506 4868 4510 4871
rect 5034 4868 5038 4871
rect 4246 4862 4249 4868
rect 4286 4863 4289 4868
rect 4198 4812 4201 4818
rect 4194 4778 4198 4781
rect 4186 4748 4190 4751
rect 4190 4732 4193 4738
rect 4170 4688 4174 4691
rect 4158 4672 4161 4678
rect 4106 4658 4110 4661
rect 4134 4632 4137 4648
rect 4150 4632 4153 4638
rect 4158 4622 4161 4668
rect 4178 4658 4182 4661
rect 4166 4642 4169 4648
rect 4082 4558 4086 4561
rect 4090 4548 4094 4551
rect 4102 4512 4105 4548
rect 4110 4542 4113 4588
rect 4130 4568 4134 4571
rect 4082 4458 4086 4461
rect 4094 4392 4097 4458
rect 4102 4412 4105 4508
rect 4112 4503 4114 4507
rect 4118 4503 4121 4507
rect 4125 4503 4128 4507
rect 4118 4472 4121 4478
rect 4142 4472 4145 4578
rect 4106 4388 4110 4391
rect 4082 4358 4086 4361
rect 4098 4348 4102 4351
rect 4078 4342 4081 4348
rect 4118 4342 4121 4468
rect 4126 4322 4129 4468
rect 4150 4462 4153 4598
rect 4190 4592 4193 4668
rect 4206 4642 4209 4788
rect 4246 4692 4249 4748
rect 4254 4672 4257 4858
rect 4318 4832 4321 4858
rect 4354 4818 4358 4821
rect 4278 4742 4281 4758
rect 4318 4742 4321 4748
rect 4330 4718 4337 4721
rect 4302 4702 4305 4718
rect 4278 4672 4281 4688
rect 4262 4663 4265 4668
rect 4202 4618 4206 4621
rect 4246 4572 4249 4618
rect 4278 4582 4281 4668
rect 4302 4661 4305 4698
rect 4318 4672 4321 4678
rect 4326 4662 4329 4668
rect 4302 4658 4310 4661
rect 4286 4572 4289 4638
rect 4294 4622 4297 4648
rect 4326 4642 4329 4648
rect 4334 4641 4337 4718
rect 4358 4692 4361 4738
rect 4354 4668 4358 4671
rect 4346 4658 4350 4661
rect 4358 4642 4361 4648
rect 4334 4638 4342 4641
rect 4310 4632 4313 4638
rect 4186 4548 4190 4551
rect 4214 4542 4217 4548
rect 4270 4542 4273 4548
rect 4278 4542 4281 4568
rect 4306 4548 4310 4551
rect 4298 4538 4302 4541
rect 4214 4522 4217 4538
rect 4134 4362 4137 4388
rect 4138 4348 4142 4351
rect 4112 4303 4114 4307
rect 4118 4303 4121 4307
rect 4125 4303 4128 4307
rect 4102 4262 4105 4298
rect 4142 4262 4145 4318
rect 4150 4302 4153 4458
rect 4158 4452 4161 4458
rect 4166 4452 4169 4458
rect 4158 4412 4161 4438
rect 4158 4352 4161 4408
rect 4166 4362 4169 4368
rect 4158 4332 4161 4338
rect 4158 4302 4161 4328
rect 4166 4262 4169 4328
rect 4198 4292 4201 4498
rect 4214 4472 4217 4518
rect 4206 4452 4209 4458
rect 4230 4392 4233 4538
rect 4254 4492 4257 4518
rect 4274 4458 4278 4461
rect 4262 4412 4265 4418
rect 4278 4412 4281 4448
rect 4278 4392 4281 4408
rect 4214 4292 4217 4368
rect 4226 4348 4230 4351
rect 4246 4342 4249 4378
rect 4286 4361 4289 4518
rect 4326 4482 4329 4578
rect 4294 4472 4297 4478
rect 4294 4452 4297 4458
rect 4334 4442 4337 4458
rect 4342 4372 4345 4638
rect 4366 4541 4369 4868
rect 4574 4862 4577 4868
rect 4602 4858 4606 4861
rect 4702 4862 4705 4868
rect 4918 4862 4921 4868
rect 4558 4822 4561 4828
rect 4414 4771 4417 4818
rect 4438 4791 4441 4818
rect 4438 4788 4449 4791
rect 4406 4768 4417 4771
rect 4374 4662 4377 4698
rect 4390 4692 4393 4747
rect 4406 4742 4409 4768
rect 4446 4762 4449 4788
rect 4446 4742 4449 4758
rect 4526 4752 4529 4758
rect 4542 4752 4545 4758
rect 4422 4682 4425 4688
rect 4382 4672 4385 4678
rect 4414 4672 4417 4678
rect 4382 4662 4385 4668
rect 4406 4662 4409 4668
rect 4390 4642 4393 4648
rect 4374 4632 4377 4638
rect 4414 4602 4417 4668
rect 4438 4662 4441 4668
rect 4446 4662 4449 4698
rect 4462 4652 4465 4728
rect 4470 4692 4473 4748
rect 4510 4722 4513 4728
rect 4486 4662 4489 4668
rect 4494 4652 4497 4668
rect 4510 4662 4513 4678
rect 4518 4672 4521 4738
rect 4526 4682 4529 4748
rect 4558 4742 4561 4818
rect 4574 4742 4577 4747
rect 4538 4738 4542 4741
rect 4534 4672 4537 4708
rect 4582 4672 4585 4718
rect 4466 4648 4473 4651
rect 4414 4572 4417 4578
rect 4386 4568 4390 4571
rect 4402 4568 4406 4571
rect 4422 4542 4425 4638
rect 4470 4572 4473 4648
rect 4518 4632 4521 4668
rect 4446 4562 4449 4568
rect 4478 4552 4481 4558
rect 4430 4542 4433 4548
rect 4494 4542 4497 4548
rect 4502 4542 4505 4618
rect 4526 4612 4529 4658
rect 4550 4652 4553 4658
rect 4558 4572 4561 4628
rect 4566 4582 4569 4658
rect 4518 4562 4521 4568
rect 4538 4558 4542 4561
rect 4566 4552 4569 4558
rect 4510 4542 4513 4548
rect 4534 4542 4537 4548
rect 4366 4538 4374 4541
rect 4562 4538 4566 4541
rect 4366 4532 4369 4538
rect 4398 4532 4401 4538
rect 4454 4532 4457 4538
rect 4390 4492 4393 4528
rect 4482 4518 4486 4521
rect 4390 4452 4393 4488
rect 4398 4472 4401 4518
rect 4446 4472 4449 4518
rect 4454 4472 4457 4488
rect 4462 4481 4465 4498
rect 4470 4491 4473 4518
rect 4470 4488 4481 4491
rect 4462 4478 4473 4481
rect 4374 4382 4377 4438
rect 4286 4358 4294 4361
rect 4310 4352 4313 4358
rect 4262 4342 4265 4348
rect 4318 4342 4321 4358
rect 4326 4342 4329 4348
rect 4278 4338 4286 4341
rect 4278 4332 4281 4338
rect 4350 4332 4353 4358
rect 4374 4352 4377 4378
rect 4386 4358 4390 4361
rect 4358 4342 4361 4348
rect 4254 4272 4257 4278
rect 4178 4268 4182 4271
rect 4266 4268 4270 4271
rect 4082 4258 4086 4261
rect 4054 4112 4057 4218
rect 4062 4152 4065 4258
rect 4070 4252 4073 4258
rect 4082 4168 4086 4171
rect 4082 4138 4086 4141
rect 4066 4088 4070 4091
rect 4046 4068 4054 4071
rect 4066 4068 4070 4071
rect 3998 4002 4001 4018
rect 3994 3978 4001 3981
rect 3998 3952 4001 3978
rect 4022 3952 4025 4018
rect 3970 3948 3974 3951
rect 3990 3942 3993 3948
rect 3974 3902 3977 3938
rect 3990 3932 3993 3938
rect 3982 3922 3985 3928
rect 3974 3882 3977 3898
rect 3986 3868 3990 3871
rect 3942 3863 3945 3868
rect 3958 3822 3961 3868
rect 3894 3818 3902 3821
rect 3894 3762 3897 3778
rect 3950 3772 3953 3798
rect 3990 3772 3993 3858
rect 3998 3852 4001 3948
rect 3898 3748 3902 3751
rect 3934 3732 3937 3738
rect 3918 3692 3921 3718
rect 3922 3678 3929 3681
rect 3914 3668 3918 3671
rect 3926 3662 3929 3678
rect 3942 3672 3945 3678
rect 3874 3658 3878 3661
rect 3854 3652 3857 3658
rect 3886 3642 3889 3658
rect 3902 3602 3905 3618
rect 3934 3612 3937 3658
rect 3942 3652 3945 3658
rect 3774 3572 3777 3598
rect 3902 3562 3905 3568
rect 3914 3558 3918 3561
rect 3750 3552 3753 3558
rect 3834 3548 3838 3551
rect 3862 3551 3865 3558
rect 3926 3552 3929 3558
rect 3934 3552 3937 3558
rect 3942 3552 3945 3558
rect 3682 3488 3686 3491
rect 3666 3468 3670 3471
rect 3542 3342 3545 3368
rect 3582 3362 3585 3368
rect 3598 3362 3601 3368
rect 3570 3358 3574 3361
rect 3550 3352 3553 3358
rect 3586 3348 3593 3351
rect 3574 3342 3577 3348
rect 3578 3338 3582 3341
rect 3486 3262 3489 3278
rect 3502 3272 3505 3278
rect 3498 3258 3502 3261
rect 3442 3248 3446 3251
rect 3430 3222 3433 3228
rect 3446 3152 3449 3158
rect 3470 3152 3473 3158
rect 3434 3138 3438 3141
rect 3458 3138 3462 3141
rect 3434 3128 3438 3131
rect 3422 3118 3433 3121
rect 3406 3012 3409 3068
rect 3414 3042 3417 3059
rect 3430 3022 3433 3118
rect 3446 3082 3449 3088
rect 3470 3081 3473 3118
rect 3478 3102 3481 3218
rect 3494 3092 3497 3258
rect 3510 3232 3513 3258
rect 3526 3222 3529 3318
rect 3542 3302 3545 3338
rect 3566 3332 3569 3338
rect 3534 3262 3537 3278
rect 3550 3262 3553 3328
rect 3590 3322 3593 3348
rect 3598 3311 3601 3358
rect 3614 3321 3617 3378
rect 3630 3342 3633 3348
rect 3654 3332 3657 3348
rect 3614 3318 3625 3321
rect 3590 3308 3601 3311
rect 3558 3262 3561 3308
rect 3542 3212 3545 3258
rect 3566 3182 3569 3218
rect 3574 3162 3577 3298
rect 3582 3262 3585 3268
rect 3574 3152 3577 3158
rect 3534 3142 3537 3148
rect 3582 3142 3585 3238
rect 3470 3078 3481 3081
rect 3462 3072 3465 3078
rect 3470 3062 3473 3068
rect 3458 3058 3462 3061
rect 3478 3051 3481 3078
rect 3494 3072 3497 3078
rect 3502 3072 3505 3078
rect 3518 3062 3521 3068
rect 3526 3062 3529 3068
rect 3474 3048 3481 3051
rect 3486 3052 3489 3058
rect 3502 3032 3505 3038
rect 3390 2962 3393 2968
rect 3462 2951 3465 2958
rect 3430 2942 3433 2948
rect 3494 2942 3497 2948
rect 3510 2942 3513 3058
rect 3534 3042 3537 3068
rect 3546 3048 3550 3051
rect 3558 3002 3561 3138
rect 3566 3062 3569 3068
rect 3574 3052 3577 3058
rect 3518 2952 3521 2978
rect 3534 2952 3537 2968
rect 3542 2952 3545 2958
rect 3530 2938 3534 2941
rect 3398 2892 3401 2918
rect 3494 2892 3497 2928
rect 3474 2888 3478 2891
rect 3462 2882 3465 2888
rect 3422 2862 3425 2868
rect 3446 2862 3449 2878
rect 3510 2872 3513 2938
rect 3478 2862 3481 2868
rect 3518 2862 3521 2928
rect 3534 2892 3537 2918
rect 3550 2892 3553 2958
rect 3566 2942 3569 2998
rect 3582 2982 3585 3108
rect 3590 3082 3593 3308
rect 3622 3292 3625 3318
rect 3610 3288 3614 3291
rect 3662 3282 3665 3438
rect 3678 3352 3681 3418
rect 3718 3392 3721 3538
rect 3742 3472 3745 3548
rect 3790 3542 3793 3548
rect 3894 3542 3897 3548
rect 3754 3538 3758 3541
rect 3902 3532 3905 3548
rect 3942 3532 3945 3548
rect 3950 3532 3953 3718
rect 3966 3692 3969 3748
rect 3982 3742 3985 3747
rect 3974 3652 3977 3678
rect 3990 3672 3993 3768
rect 3998 3702 4001 3838
rect 4006 3802 4009 3918
rect 4038 3912 4041 4058
rect 4046 4052 4049 4058
rect 4078 4052 4081 4088
rect 4094 4062 4097 4218
rect 4126 4152 4129 4208
rect 4112 4103 4114 4107
rect 4118 4103 4121 4107
rect 4125 4103 4128 4107
rect 4086 4052 4089 4058
rect 4046 3901 4049 3998
rect 4102 3982 4105 4018
rect 4118 3992 4121 4058
rect 4126 4002 4129 4058
rect 4134 4022 4137 4258
rect 4206 4252 4209 4258
rect 4198 4232 4201 4248
rect 4222 4242 4225 4268
rect 4230 4262 4233 4268
rect 4242 4258 4246 4261
rect 4278 4252 4281 4308
rect 4286 4282 4289 4328
rect 4338 4318 4342 4321
rect 4366 4312 4369 4348
rect 4286 4262 4289 4268
rect 4234 4248 4238 4251
rect 4270 4248 4278 4251
rect 4154 4218 4158 4221
rect 4202 4168 4206 4171
rect 4190 4162 4193 4168
rect 4154 4147 4158 4150
rect 4206 4132 4209 4148
rect 4214 4142 4217 4178
rect 4222 4162 4225 4168
rect 4238 4152 4241 4158
rect 4226 4148 4230 4151
rect 4246 4142 4249 4148
rect 4246 4118 4254 4121
rect 4206 4092 4209 4108
rect 4246 4082 4249 4118
rect 4222 4078 4238 4081
rect 4222 4072 4225 4078
rect 4186 4068 4190 4071
rect 4234 4068 4238 4071
rect 4166 4052 4169 4058
rect 4150 4042 4153 4048
rect 4106 3958 4110 3961
rect 4038 3898 4049 3901
rect 4014 3862 4017 3868
rect 4022 3852 4025 3858
rect 4014 3752 4017 3818
rect 3998 3672 4001 3698
rect 3958 3592 3961 3618
rect 3974 3572 3977 3648
rect 3990 3631 3993 3658
rect 3982 3628 3993 3631
rect 3742 3452 3745 3458
rect 3706 3368 3710 3371
rect 3734 3358 3742 3361
rect 3750 3361 3753 3498
rect 3766 3452 3769 3518
rect 3782 3472 3785 3478
rect 3806 3462 3809 3468
rect 3814 3462 3817 3508
rect 3902 3502 3905 3528
rect 3822 3462 3825 3468
rect 3870 3462 3873 3478
rect 3910 3472 3913 3478
rect 3894 3462 3897 3468
rect 3922 3458 3926 3461
rect 3790 3442 3793 3458
rect 3846 3452 3849 3458
rect 3802 3448 3806 3451
rect 3902 3422 3905 3458
rect 3914 3448 3918 3451
rect 3930 3448 3934 3451
rect 3942 3442 3945 3468
rect 3950 3462 3953 3518
rect 3958 3472 3961 3568
rect 3966 3512 3969 3528
rect 3982 3522 3985 3628
rect 3966 3452 3969 3498
rect 3974 3452 3977 3518
rect 3990 3482 3993 3538
rect 3998 3532 4001 3668
rect 4014 3662 4017 3688
rect 4038 3662 4041 3898
rect 4054 3892 4057 3948
rect 4118 3942 4121 3958
rect 4134 3942 4137 3948
rect 4062 3862 4065 3888
rect 4086 3882 4089 3938
rect 4102 3922 4105 3938
rect 4112 3903 4114 3907
rect 4118 3903 4121 3907
rect 4125 3903 4128 3907
rect 4134 3892 4137 3898
rect 4070 3792 4073 3858
rect 4086 3822 4089 3858
rect 4102 3762 4105 3848
rect 4126 3762 4129 3798
rect 4126 3752 4129 3758
rect 4054 3742 4057 3748
rect 4078 3742 4081 3748
rect 4122 3738 4126 3741
rect 4046 3682 4049 3718
rect 4074 3668 4078 3671
rect 4058 3658 4062 3661
rect 4006 3652 4009 3658
rect 4022 3592 4025 3618
rect 4054 3572 4057 3648
rect 4086 3632 4089 3738
rect 4094 3642 4097 3658
rect 4102 3631 4105 3718
rect 4112 3703 4114 3707
rect 4118 3703 4121 3707
rect 4125 3703 4128 3707
rect 4134 3672 4137 3878
rect 4142 3872 4145 3998
rect 4150 3952 4153 4028
rect 4182 3992 4185 4038
rect 4190 4022 4193 4058
rect 4214 4022 4217 4048
rect 4254 4002 4257 4068
rect 4262 4062 4265 4128
rect 4262 4002 4265 4058
rect 4270 4022 4273 4248
rect 4278 4052 4281 4058
rect 4286 4012 4289 4258
rect 4302 4222 4305 4278
rect 4322 4268 4326 4271
rect 4334 4262 4337 4288
rect 4374 4272 4377 4348
rect 4398 4262 4401 4468
rect 4462 4462 4465 4468
rect 4470 4462 4473 4478
rect 4410 4458 4414 4461
rect 4426 4448 4430 4451
rect 4410 4438 4414 4441
rect 4446 4412 4449 4458
rect 4430 4352 4433 4358
rect 4318 4252 4321 4258
rect 4366 4252 4369 4259
rect 4438 4232 4441 4238
rect 4434 4218 4438 4221
rect 4446 4202 4449 4408
rect 4454 4342 4457 4348
rect 4350 4152 4353 4158
rect 4274 3988 4278 3991
rect 4166 3962 4169 3968
rect 4150 3872 4153 3948
rect 4142 3842 4145 3868
rect 4154 3858 4158 3861
rect 4166 3852 4169 3918
rect 4174 3912 4177 3958
rect 4174 3902 4177 3908
rect 4182 3892 4185 3968
rect 4194 3958 4198 3961
rect 4242 3958 4246 3961
rect 4214 3951 4217 3958
rect 4214 3948 4225 3951
rect 4198 3942 4201 3948
rect 4190 3922 4193 3938
rect 4198 3922 4201 3938
rect 4214 3882 4217 3938
rect 4222 3892 4225 3948
rect 4250 3948 4254 3951
rect 4150 3762 4153 3818
rect 4166 3791 4169 3838
rect 4162 3788 4169 3791
rect 4174 3772 4177 3818
rect 4190 3812 4193 3868
rect 4198 3842 4201 3868
rect 4210 3858 4214 3861
rect 4222 3852 4225 3888
rect 4230 3882 4233 3948
rect 4262 3942 4265 3948
rect 4250 3938 4254 3941
rect 4238 3861 4241 3918
rect 4258 3888 4262 3891
rect 4250 3868 4254 3871
rect 4294 3862 4297 4138
rect 4302 4112 4305 4148
rect 4334 4112 4337 4138
rect 4318 4082 4321 4088
rect 4314 4068 4318 4071
rect 4302 4062 4305 4068
rect 4334 4062 4337 4088
rect 4306 4048 4310 4051
rect 4302 3952 4305 3958
rect 4318 3942 4321 3948
rect 4326 3942 4329 4018
rect 4350 3962 4353 4148
rect 4358 4142 4361 4198
rect 4382 4152 4385 4198
rect 4454 4182 4457 4268
rect 4462 4252 4465 4458
rect 4478 4362 4481 4488
rect 4490 4468 4494 4471
rect 4510 4462 4513 4488
rect 4494 4422 4497 4448
rect 4518 4432 4521 4468
rect 4522 4418 4526 4421
rect 4498 4358 4502 4361
rect 4510 4352 4513 4358
rect 4506 4348 4510 4351
rect 4518 4342 4521 4388
rect 4478 4292 4481 4338
rect 4534 4332 4537 4418
rect 4542 4412 4545 4538
rect 4574 4482 4577 4668
rect 4590 4642 4593 4658
rect 4598 4622 4601 4728
rect 4606 4692 4609 4848
rect 4622 4792 4625 4818
rect 4632 4803 4634 4807
rect 4638 4803 4641 4807
rect 4645 4803 4648 4807
rect 4678 4792 4681 4838
rect 4686 4832 4689 4859
rect 4866 4858 4870 4861
rect 4750 4842 4753 4858
rect 4774 4852 4777 4858
rect 4846 4852 4849 4858
rect 4934 4852 4937 4859
rect 5026 4858 5030 4861
rect 5070 4852 5073 4858
rect 5102 4852 5105 4859
rect 5006 4842 5009 4848
rect 4810 4818 4814 4821
rect 4622 4772 4625 4778
rect 4694 4772 4697 4818
rect 4902 4812 4905 4818
rect 5022 4802 5025 4818
rect 5038 4812 5041 4818
rect 4614 4652 4617 4708
rect 4622 4672 4625 4748
rect 4638 4712 4641 4718
rect 4662 4692 4665 4758
rect 4750 4752 4753 4778
rect 4830 4752 4833 4768
rect 4682 4748 4686 4751
rect 4842 4748 4846 4751
rect 4686 4702 4689 4738
rect 4634 4668 4638 4671
rect 4638 4652 4641 4658
rect 4654 4652 4657 4688
rect 4682 4668 4686 4671
rect 4678 4652 4681 4658
rect 4694 4652 4697 4718
rect 4710 4711 4713 4738
rect 4722 4718 4729 4721
rect 4710 4708 4721 4711
rect 4606 4642 4609 4648
rect 4582 4572 4585 4618
rect 4614 4572 4617 4648
rect 4678 4642 4681 4648
rect 4632 4603 4634 4607
rect 4638 4603 4641 4607
rect 4645 4603 4648 4607
rect 4614 4532 4617 4558
rect 4590 4512 4593 4518
rect 4582 4462 4585 4468
rect 4542 4392 4545 4398
rect 4550 4332 4553 4408
rect 4558 4332 4561 4338
rect 4494 4322 4497 4328
rect 4526 4282 4529 4318
rect 4566 4292 4569 4458
rect 4606 4452 4609 4518
rect 4630 4482 4633 4568
rect 4654 4492 4657 4638
rect 4678 4582 4681 4638
rect 4606 4412 4609 4448
rect 4654 4442 4657 4448
rect 4574 4312 4577 4358
rect 4598 4352 4601 4358
rect 4622 4342 4625 4418
rect 4632 4403 4634 4407
rect 4638 4403 4641 4407
rect 4645 4403 4648 4407
rect 4662 4352 4665 4548
rect 4678 4492 4681 4578
rect 4686 4522 4689 4547
rect 4674 4468 4678 4471
rect 4694 4462 4697 4488
rect 4702 4472 4705 4668
rect 4710 4652 4713 4658
rect 4710 4612 4713 4618
rect 4718 4542 4721 4708
rect 4726 4682 4729 4718
rect 4766 4692 4769 4748
rect 4854 4742 4857 4768
rect 4862 4752 4865 4758
rect 4902 4752 4905 4778
rect 4994 4758 4998 4761
rect 4922 4748 4926 4751
rect 4986 4748 4990 4751
rect 4814 4722 4817 4728
rect 4950 4722 4953 4738
rect 4866 4718 4870 4721
rect 4858 4678 4862 4681
rect 4818 4668 4822 4671
rect 4746 4658 4750 4661
rect 4774 4652 4777 4668
rect 4790 4652 4793 4658
rect 4730 4568 4734 4571
rect 4742 4562 4745 4568
rect 4722 4538 4726 4541
rect 4738 4528 4745 4531
rect 4710 4492 4713 4518
rect 4734 4472 4737 4518
rect 4674 4448 4678 4451
rect 4694 4442 4697 4448
rect 4702 4402 4705 4468
rect 4722 4458 4726 4461
rect 4710 4442 4713 4448
rect 4734 4412 4737 4468
rect 4742 4452 4745 4528
rect 4750 4462 4753 4648
rect 4782 4482 4785 4618
rect 4798 4562 4801 4648
rect 4814 4642 4817 4658
rect 4814 4602 4817 4618
rect 4830 4592 4833 4668
rect 4886 4662 4889 4668
rect 4942 4662 4945 4678
rect 4950 4672 4953 4718
rect 4966 4702 4969 4738
rect 4842 4658 4846 4661
rect 4838 4562 4841 4598
rect 4802 4547 4806 4550
rect 4842 4548 4846 4551
rect 4822 4532 4825 4538
rect 4854 4502 4857 4658
rect 4862 4642 4865 4648
rect 4862 4552 4865 4588
rect 4870 4542 4873 4658
rect 4878 4652 4881 4658
rect 4878 4552 4881 4648
rect 4890 4638 4894 4641
rect 4930 4568 4934 4571
rect 4894 4562 4897 4568
rect 4906 4548 4910 4551
rect 4862 4532 4865 4538
rect 4854 4492 4857 4498
rect 4862 4492 4865 4498
rect 4798 4482 4801 4488
rect 4818 4468 4822 4471
rect 4754 4458 4758 4461
rect 4810 4458 4814 4461
rect 4838 4452 4841 4458
rect 4846 4452 4849 4458
rect 4826 4438 4830 4441
rect 4738 4358 4742 4361
rect 4694 4351 4697 4358
rect 4634 4318 4638 4321
rect 4566 4272 4569 4288
rect 4478 4242 4481 4258
rect 4486 4252 4489 4268
rect 4494 4262 4497 4268
rect 4506 4258 4510 4261
rect 4510 4232 4513 4248
rect 4462 4172 4465 4218
rect 4374 4142 4377 4148
rect 4402 4138 4406 4141
rect 4422 4132 4425 4158
rect 4402 4128 4406 4131
rect 4430 4122 4433 4128
rect 4446 4122 4449 4148
rect 4454 4142 4457 4168
rect 4478 4152 4481 4198
rect 4494 4192 4497 4228
rect 4510 4218 4518 4221
rect 4486 4142 4489 4188
rect 4510 4162 4513 4218
rect 4478 4132 4481 4138
rect 4510 4132 4513 4158
rect 4518 4142 4521 4208
rect 4526 4182 4529 4268
rect 4562 4258 4566 4261
rect 4526 4152 4529 4178
rect 4566 4162 4569 4178
rect 4574 4162 4577 4168
rect 4542 4152 4545 4158
rect 4566 4152 4569 4158
rect 4538 4138 4542 4141
rect 4554 4138 4558 4141
rect 4414 4072 4417 4108
rect 4442 4088 4446 4091
rect 4430 4072 4433 4078
rect 4446 4062 4449 4068
rect 4390 4052 4393 4058
rect 4462 4051 4465 4118
rect 4486 4082 4489 4128
rect 4482 4068 4486 4071
rect 4558 4062 4561 4098
rect 4474 4058 4478 4061
rect 4458 4048 4465 4051
rect 4398 3992 4401 4048
rect 4446 4042 4449 4048
rect 4382 3952 4385 3958
rect 4354 3948 4358 3951
rect 4350 3932 4353 3948
rect 4374 3942 4377 3948
rect 4390 3942 4393 3948
rect 4334 3912 4337 3928
rect 4238 3858 4246 3861
rect 4238 3802 4241 3858
rect 4250 3848 4254 3851
rect 4150 3742 4153 3748
rect 4182 3672 4185 3678
rect 4198 3672 4201 3748
rect 4206 3742 4209 3748
rect 4222 3742 4225 3758
rect 4222 3682 4225 3688
rect 4214 3678 4222 3681
rect 4154 3658 4158 3661
rect 4214 3652 4217 3678
rect 4238 3672 4241 3768
rect 4254 3752 4257 3828
rect 4294 3762 4297 3858
rect 4318 3852 4321 3858
rect 4306 3758 4310 3761
rect 4314 3748 4318 3751
rect 4262 3742 4265 3748
rect 4286 3732 4289 3748
rect 4326 3742 4329 3768
rect 4342 3762 4345 3908
rect 4366 3902 4369 3918
rect 4398 3872 4401 3958
rect 4406 3932 4409 3998
rect 4414 3942 4417 3968
rect 4430 3962 4433 4038
rect 4506 4028 4510 4031
rect 4478 3952 4481 3958
rect 4486 3952 4489 3988
rect 4442 3948 4446 3951
rect 4466 3948 4470 3951
rect 4410 3928 4414 3931
rect 4430 3872 4433 3918
rect 4454 3891 4457 3918
rect 4494 3892 4497 4018
rect 4526 3972 4529 4018
rect 4566 4002 4569 4118
rect 4582 4082 4585 4318
rect 4662 4292 4665 4348
rect 4726 4322 4729 4358
rect 4670 4282 4673 4318
rect 4702 4292 4705 4308
rect 4742 4272 4745 4348
rect 4750 4342 4753 4398
rect 4758 4382 4761 4418
rect 4762 4358 4766 4361
rect 4770 4348 4774 4351
rect 4758 4342 4761 4348
rect 4750 4332 4753 4338
rect 4774 4322 4777 4348
rect 4782 4342 4785 4408
rect 4790 4312 4793 4358
rect 4798 4352 4801 4358
rect 4806 4352 4809 4358
rect 4678 4262 4681 4268
rect 4766 4263 4769 4298
rect 4798 4272 4801 4278
rect 4626 4258 4630 4261
rect 4694 4252 4697 4258
rect 4618 4248 4622 4251
rect 4674 4248 4678 4251
rect 4630 4222 4633 4228
rect 4718 4221 4721 4238
rect 4782 4232 4785 4268
rect 4806 4262 4809 4348
rect 4814 4342 4817 4428
rect 4838 4412 4841 4448
rect 4822 4352 4825 4358
rect 4814 4292 4817 4338
rect 4822 4302 4825 4318
rect 4814 4272 4817 4288
rect 4830 4272 4833 4278
rect 4802 4258 4806 4261
rect 4838 4261 4841 4348
rect 4846 4342 4849 4378
rect 4854 4352 4857 4488
rect 4870 4481 4873 4538
rect 4878 4502 4881 4548
rect 4918 4492 4921 4548
rect 4926 4532 4929 4538
rect 4966 4532 4969 4538
rect 4974 4532 4977 4748
rect 4990 4672 4993 4678
rect 4990 4652 4993 4658
rect 4998 4622 5001 4718
rect 5014 4692 5017 4758
rect 5042 4748 5046 4751
rect 5030 4722 5033 4748
rect 5126 4722 5129 4748
rect 5050 4668 5054 4671
rect 5022 4662 5025 4668
rect 5074 4658 5078 4661
rect 5014 4622 5017 4648
rect 5022 4571 5025 4658
rect 5030 4652 5033 4658
rect 5054 4652 5057 4658
rect 5034 4648 5041 4651
rect 5022 4568 5033 4571
rect 4986 4548 4990 4551
rect 5030 4542 5033 4568
rect 5038 4552 5041 4648
rect 5046 4632 5049 4648
rect 5050 4558 5054 4561
rect 4862 4478 4873 4481
rect 4862 4432 4865 4478
rect 4998 4472 5001 4528
rect 5062 4492 5065 4658
rect 5074 4648 5078 4651
rect 5082 4628 5086 4631
rect 5078 4592 5081 4618
rect 5094 4562 5097 4718
rect 5134 4672 5137 4858
rect 5150 4842 5153 4848
rect 5154 4818 5158 4821
rect 5130 4658 5134 4661
rect 5142 4622 5145 4748
rect 5150 4682 5153 4738
rect 5162 4558 5166 4561
rect 5078 4492 5081 4548
rect 5178 4538 5182 4541
rect 5086 4512 5089 4538
rect 5022 4472 5025 4478
rect 5062 4472 5065 4478
rect 5078 4472 5081 4478
rect 5094 4472 5097 4538
rect 4930 4468 4934 4471
rect 4862 4402 4865 4418
rect 4862 4352 4865 4358
rect 4854 4332 4857 4338
rect 4870 4332 4873 4468
rect 4890 4458 4897 4461
rect 4878 4352 4881 4358
rect 4894 4352 4897 4458
rect 4922 4448 4926 4451
rect 4902 4422 4905 4448
rect 4934 4372 4937 4458
rect 4990 4452 4993 4458
rect 4946 4418 4950 4421
rect 4906 4358 4910 4361
rect 4858 4268 4862 4271
rect 4838 4258 4846 4261
rect 4822 4222 4825 4248
rect 4718 4218 4729 4221
rect 4858 4218 4862 4221
rect 4632 4203 4634 4207
rect 4638 4203 4641 4207
rect 4645 4203 4648 4207
rect 4626 4148 4630 4151
rect 4654 4112 4657 4138
rect 4646 4092 4649 4098
rect 4582 4062 4585 4068
rect 4598 4032 4601 4078
rect 4526 3962 4529 3968
rect 4502 3922 4505 3928
rect 4454 3888 4462 3891
rect 4478 3872 4481 3888
rect 4398 3862 4401 3868
rect 4486 3862 4489 3868
rect 4370 3858 4374 3861
rect 4434 3858 4438 3861
rect 4458 3858 4462 3861
rect 4474 3858 4478 3861
rect 4502 3861 4505 3918
rect 4498 3858 4505 3861
rect 4390 3852 4393 3858
rect 4414 3841 4417 3858
rect 4414 3838 4422 3841
rect 4378 3828 4382 3831
rect 4270 3702 4273 3718
rect 4274 3688 4278 3691
rect 4258 3668 4262 3671
rect 4238 3662 4241 3668
rect 4266 3658 4270 3661
rect 4254 3652 4257 3658
rect 4102 3628 4110 3631
rect 4050 3548 4054 3551
rect 4078 3542 4081 3568
rect 4094 3552 4097 3588
rect 3998 3512 4001 3518
rect 4038 3482 4041 3538
rect 4034 3459 4038 3462
rect 4086 3462 4089 3518
rect 4094 3472 4097 3528
rect 4102 3502 4105 3618
rect 4118 3572 4121 3638
rect 4110 3522 4113 3528
rect 4112 3503 4114 3507
rect 4118 3503 4121 3507
rect 4125 3503 4128 3507
rect 4134 3472 4137 3598
rect 4182 3562 4185 3568
rect 4158 3552 4161 3558
rect 4190 3552 4193 3628
rect 4206 3572 4209 3618
rect 4222 3562 4225 3568
rect 4178 3548 4182 3551
rect 4142 3532 4145 3538
rect 4142 3462 4145 3518
rect 4150 3462 4153 3468
rect 4098 3458 4102 3461
rect 4118 3452 4121 3458
rect 4098 3448 4102 3451
rect 3830 3412 3833 3418
rect 3750 3358 3761 3361
rect 3722 3348 3726 3351
rect 3710 3341 3713 3348
rect 3710 3338 3718 3341
rect 3734 3332 3737 3358
rect 3746 3348 3750 3351
rect 3718 3282 3721 3308
rect 3598 3272 3601 3278
rect 3654 3262 3657 3268
rect 3726 3262 3729 3268
rect 3670 3258 3678 3261
rect 3670 3252 3673 3258
rect 3682 3248 3686 3251
rect 3608 3203 3610 3207
rect 3614 3203 3617 3207
rect 3621 3203 3624 3207
rect 3610 3148 3614 3151
rect 3622 3142 3625 3148
rect 3622 3082 3625 3138
rect 3630 3132 3633 3238
rect 3638 3192 3641 3238
rect 3694 3232 3697 3258
rect 3670 3191 3673 3218
rect 3670 3188 3681 3191
rect 3618 3068 3622 3071
rect 3590 3062 3593 3068
rect 3646 3052 3649 3118
rect 3586 2947 3590 2950
rect 3598 2901 3601 3018
rect 3630 3012 3633 3038
rect 3608 3003 3610 3007
rect 3614 3003 3617 3007
rect 3621 3003 3624 3007
rect 3614 2932 3617 2938
rect 3590 2898 3601 2901
rect 3378 2858 3385 2861
rect 3506 2858 3510 2861
rect 3366 2842 3369 2858
rect 3398 2832 3401 2858
rect 3386 2828 3390 2831
rect 3286 2792 3289 2818
rect 3350 2792 3353 2808
rect 3290 2738 3294 2741
rect 3302 2672 3305 2698
rect 3334 2672 3337 2678
rect 3294 2652 3297 2658
rect 3222 2542 3225 2548
rect 3214 2532 3217 2538
rect 3278 2492 3281 2618
rect 3318 2592 3321 2648
rect 3334 2632 3337 2648
rect 3342 2552 3345 2788
rect 3366 2732 3369 2738
rect 3362 2668 3366 2671
rect 3374 2662 3377 2768
rect 3430 2752 3433 2818
rect 3446 2792 3449 2848
rect 3430 2712 3433 2738
rect 3430 2682 3433 2708
rect 3394 2668 3398 2671
rect 3386 2658 3390 2661
rect 3430 2652 3433 2659
rect 3370 2648 3374 2651
rect 3390 2642 3393 2648
rect 3358 2602 3361 2618
rect 3322 2548 3326 2551
rect 3286 2532 3289 2538
rect 3294 2532 3297 2548
rect 3374 2542 3377 2547
rect 3310 2512 3313 2528
rect 3326 2522 3329 2538
rect 3334 2532 3337 2538
rect 3266 2488 3270 2491
rect 3294 2472 3297 2488
rect 3334 2472 3337 2498
rect 3130 2468 3134 2471
rect 3146 2468 3150 2471
rect 3170 2468 3174 2471
rect 3242 2468 3246 2471
rect 3078 2462 3081 2468
rect 2990 2392 2993 2458
rect 2998 2372 3001 2418
rect 3014 2412 3017 2458
rect 3022 2452 3025 2458
rect 3062 2452 3065 2458
rect 3014 2372 3017 2378
rect 2942 2358 2950 2361
rect 2942 2352 2945 2358
rect 2974 2352 2977 2358
rect 2954 2348 2958 2351
rect 2926 2318 2934 2321
rect 2926 2282 2929 2318
rect 2886 2232 2889 2238
rect 2894 2162 2897 2268
rect 2918 2262 2921 2278
rect 2942 2272 2945 2338
rect 2974 2282 2977 2348
rect 2986 2338 2990 2341
rect 2962 2278 2966 2281
rect 2998 2281 3001 2348
rect 2998 2278 3006 2281
rect 2974 2262 2977 2268
rect 2990 2262 2993 2278
rect 2998 2262 3001 2278
rect 3014 2272 3017 2278
rect 2902 2222 2905 2258
rect 2942 2242 2945 2258
rect 3010 2228 3014 2231
rect 2926 2152 2929 2168
rect 2958 2152 2961 2228
rect 2966 2182 2969 2218
rect 2982 2152 2985 2158
rect 2998 2152 3001 2168
rect 3006 2162 3009 2168
rect 2886 2142 2889 2148
rect 2894 2142 2897 2148
rect 2838 2132 2841 2138
rect 2866 2128 2870 2131
rect 2822 2072 2825 2088
rect 2830 2062 2833 2068
rect 2814 2052 2817 2058
rect 2822 2051 2825 2058
rect 2846 2052 2849 2118
rect 2878 2072 2881 2118
rect 2910 2082 2913 2148
rect 2866 2058 2870 2061
rect 2910 2052 2913 2059
rect 2822 2048 2838 2051
rect 2858 2048 2862 2051
rect 2874 2048 2878 2051
rect 2750 1942 2753 2038
rect 2758 2012 2761 2018
rect 2782 2012 2785 2018
rect 2814 1972 2817 2048
rect 2830 2012 2833 2018
rect 2774 1962 2777 1968
rect 2758 1952 2761 1958
rect 2750 1892 2753 1938
rect 2806 1902 2809 1948
rect 2838 1942 2841 1947
rect 2870 1932 2873 1958
rect 2878 1921 2881 1978
rect 2918 1952 2921 2148
rect 2942 2142 2945 2148
rect 2950 2142 2953 2148
rect 2926 2062 2929 2138
rect 2934 2112 2937 2138
rect 2974 2132 2977 2138
rect 2934 2082 2937 2108
rect 2982 2072 2985 2118
rect 2990 2112 2993 2138
rect 3006 2112 3009 2118
rect 2998 1992 3001 2058
rect 3014 2042 3017 2168
rect 3022 2152 3025 2388
rect 3030 2332 3033 2348
rect 3046 2312 3049 2318
rect 3030 2262 3033 2308
rect 3046 2262 3049 2278
rect 3030 2172 3033 2218
rect 3046 2192 3049 2258
rect 3054 2192 3057 2318
rect 3062 2282 3065 2448
rect 3086 2352 3089 2398
rect 3094 2372 3097 2468
rect 3182 2461 3185 2468
rect 3198 2462 3201 2468
rect 3170 2458 3185 2461
rect 3102 2452 3105 2458
rect 3118 2392 3121 2458
rect 3142 2422 3145 2438
rect 3142 2352 3145 2418
rect 3150 2392 3153 2458
rect 3182 2442 3185 2448
rect 3190 2412 3193 2458
rect 3206 2442 3209 2458
rect 3190 2392 3193 2398
rect 3206 2362 3209 2408
rect 3166 2352 3169 2358
rect 3174 2342 3177 2348
rect 3070 2332 3073 2338
rect 3118 2312 3121 2318
rect 3096 2303 3098 2307
rect 3102 2303 3105 2307
rect 3109 2303 3112 2307
rect 3070 2292 3073 2298
rect 3062 2232 3065 2258
rect 3058 2158 3062 2161
rect 3042 2138 3054 2141
rect 3022 2082 3025 2138
rect 3054 2122 3057 2128
rect 3070 2081 3073 2268
rect 3094 2262 3097 2268
rect 3086 2242 3089 2258
rect 3102 2252 3105 2258
rect 3078 2152 3081 2168
rect 3118 2152 3121 2308
rect 3186 2268 3190 2271
rect 3138 2248 3142 2251
rect 3106 2148 3110 2151
rect 3078 2132 3081 2138
rect 3070 2078 3081 2081
rect 3078 2072 3081 2078
rect 3030 2052 3033 2068
rect 3070 2062 3073 2068
rect 2986 1958 2990 1961
rect 2946 1948 2950 1951
rect 2978 1948 2982 1951
rect 2886 1942 2889 1948
rect 2894 1942 2897 1948
rect 2910 1942 2913 1948
rect 2870 1918 2881 1921
rect 2786 1888 2790 1891
rect 2806 1882 2809 1898
rect 2870 1892 2873 1918
rect 2802 1868 2806 1871
rect 2866 1868 2870 1871
rect 2662 1752 2665 1758
rect 2722 1748 2726 1751
rect 2738 1748 2742 1751
rect 2706 1738 2710 1741
rect 2614 1672 2617 1708
rect 2670 1692 2673 1728
rect 2630 1652 2633 1678
rect 2622 1562 2625 1618
rect 2630 1552 2633 1558
rect 2638 1542 2641 1558
rect 2646 1552 2649 1678
rect 2670 1672 2673 1688
rect 2682 1658 2686 1661
rect 2694 1612 2697 1658
rect 2718 1652 2721 1718
rect 2730 1688 2734 1691
rect 2750 1682 2753 1828
rect 2798 1762 2801 1818
rect 2774 1758 2782 1761
rect 2774 1752 2777 1758
rect 2774 1692 2777 1738
rect 2782 1712 2785 1748
rect 2814 1742 2817 1868
rect 2886 1862 2889 1868
rect 2854 1852 2857 1858
rect 2838 1802 2841 1818
rect 2766 1682 2769 1688
rect 2734 1662 2737 1668
rect 2750 1662 2753 1678
rect 2786 1668 2790 1671
rect 2730 1648 2734 1651
rect 2750 1552 2753 1588
rect 2722 1548 2726 1551
rect 2618 1538 2622 1541
rect 2642 1538 2646 1541
rect 2638 1492 2641 1498
rect 2634 1468 2638 1471
rect 2654 1462 2657 1548
rect 2670 1532 2673 1538
rect 2670 1492 2673 1498
rect 2618 1458 2622 1461
rect 2650 1458 2654 1461
rect 2650 1448 2654 1451
rect 2482 1368 2486 1371
rect 2426 1348 2430 1351
rect 2470 1342 2473 1358
rect 2558 1352 2561 1368
rect 2510 1342 2513 1348
rect 2454 1332 2457 1338
rect 2478 1292 2481 1338
rect 2410 1258 2414 1261
rect 2390 1152 2393 1218
rect 2422 1211 2425 1278
rect 2462 1262 2465 1288
rect 2434 1258 2438 1261
rect 2450 1238 2454 1241
rect 2418 1208 2425 1211
rect 2406 1162 2409 1168
rect 2414 1151 2417 1208
rect 2422 1162 2425 1168
rect 2446 1162 2449 1168
rect 2414 1148 2422 1151
rect 2410 1138 2414 1141
rect 2282 1058 2286 1061
rect 2254 1042 2257 1048
rect 2278 1042 2281 1048
rect 2226 948 2230 951
rect 2178 938 2182 941
rect 2174 932 2177 938
rect 2150 878 2161 881
rect 2138 868 2142 871
rect 2126 812 2129 868
rect 2134 792 2137 848
rect 1926 692 1929 748
rect 1942 742 1945 747
rect 1974 742 1977 748
rect 1906 658 1910 661
rect 1922 648 1926 651
rect 1866 568 1873 571
rect 1878 561 1881 618
rect 1870 558 1881 561
rect 1838 531 1841 548
rect 1862 542 1865 558
rect 1830 528 1841 531
rect 1798 492 1801 508
rect 1822 472 1825 488
rect 1830 462 1833 528
rect 1570 368 1574 371
rect 1666 368 1670 371
rect 1750 362 1753 368
rect 1674 358 1678 361
rect 1566 292 1569 358
rect 1694 352 1697 358
rect 1734 352 1737 358
rect 1606 332 1609 347
rect 1750 342 1753 348
rect 1758 342 1761 368
rect 1766 362 1769 368
rect 1706 338 1710 341
rect 1606 292 1609 308
rect 1582 262 1585 278
rect 1606 272 1609 288
rect 1598 262 1601 268
rect 1550 192 1553 248
rect 1582 232 1585 258
rect 1598 242 1601 248
rect 1606 222 1609 258
rect 1614 242 1617 248
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1573 203 1576 207
rect 1554 188 1558 191
rect 1582 112 1585 148
rect 1606 142 1609 218
rect 1622 142 1625 338
rect 1710 282 1713 328
rect 1726 282 1729 338
rect 1734 292 1737 338
rect 1662 263 1665 268
rect 1630 242 1633 248
rect 1686 232 1689 258
rect 1742 252 1745 278
rect 1758 271 1761 338
rect 1766 322 1769 348
rect 1822 311 1825 458
rect 1830 322 1833 458
rect 1846 452 1849 478
rect 1858 468 1862 471
rect 1870 352 1873 558
rect 1878 532 1881 548
rect 1886 542 1889 578
rect 1926 552 1929 558
rect 1902 542 1905 548
rect 1886 501 1889 538
rect 1934 522 1937 668
rect 1942 662 1945 668
rect 1958 652 1961 708
rect 1966 672 1969 728
rect 1990 682 1993 688
rect 1974 662 1977 678
rect 1998 672 2001 718
rect 2006 712 2009 718
rect 2006 662 2009 668
rect 2014 661 2017 708
rect 2010 658 2017 661
rect 1946 648 1950 651
rect 1994 648 2006 651
rect 1966 572 1969 638
rect 1982 592 1985 628
rect 2006 562 2009 568
rect 2014 562 2017 658
rect 2022 582 2025 718
rect 2030 652 2033 688
rect 2038 682 2041 748
rect 2094 742 2097 788
rect 2122 758 2126 761
rect 2122 748 2126 751
rect 2150 742 2153 878
rect 2182 862 2185 918
rect 2206 902 2209 938
rect 2214 932 2217 938
rect 2238 892 2241 958
rect 2250 918 2254 921
rect 2222 872 2225 888
rect 2262 882 2265 918
rect 2278 892 2281 938
rect 2254 872 2257 878
rect 2166 742 2169 747
rect 2094 732 2097 738
rect 2150 732 2153 738
rect 2054 712 2057 718
rect 2072 703 2074 707
rect 2078 703 2081 707
rect 2085 703 2088 707
rect 2126 692 2129 728
rect 2130 688 2134 691
rect 2022 562 2025 568
rect 2014 552 2017 558
rect 2038 552 2041 658
rect 2054 642 2057 668
rect 2070 652 2073 659
rect 2086 642 2089 678
rect 2026 548 2030 551
rect 1878 498 1889 501
rect 1878 472 1881 498
rect 1886 482 1889 488
rect 1950 482 1953 538
rect 1934 462 1937 468
rect 1878 432 1881 458
rect 1910 392 1913 418
rect 1966 392 1969 528
rect 1990 492 1993 538
rect 2014 522 2017 538
rect 2006 462 2009 478
rect 2014 472 2017 518
rect 2038 502 2041 548
rect 2046 542 2049 578
rect 2090 568 2094 571
rect 2118 562 2121 638
rect 2054 552 2057 558
rect 2110 542 2113 548
rect 2118 542 2121 548
rect 2126 542 2129 678
rect 2174 672 2177 698
rect 2190 692 2193 748
rect 2222 682 2225 868
rect 2274 858 2278 861
rect 2238 772 2241 848
rect 2238 752 2241 758
rect 2254 752 2257 808
rect 2262 742 2265 828
rect 2286 792 2289 1008
rect 2294 1002 2297 1058
rect 2334 1052 2337 1059
rect 2342 992 2345 1128
rect 2382 1082 2385 1138
rect 2406 1122 2409 1128
rect 2394 1088 2398 1091
rect 2382 1052 2385 1078
rect 2406 1072 2409 1098
rect 2422 1061 2425 1148
rect 2430 1092 2433 1148
rect 2454 1141 2457 1178
rect 2462 1162 2465 1168
rect 2470 1162 2473 1258
rect 2450 1138 2457 1141
rect 2422 1058 2430 1061
rect 2406 1052 2409 1058
rect 2406 1002 2409 1048
rect 2430 1042 2433 1048
rect 2382 951 2385 958
rect 2294 892 2297 948
rect 2326 942 2329 948
rect 2342 921 2345 948
rect 2350 942 2353 948
rect 2334 918 2345 921
rect 2350 922 2353 928
rect 2302 862 2305 868
rect 2310 862 2313 898
rect 2334 892 2337 918
rect 2318 862 2321 888
rect 2366 882 2369 918
rect 2382 892 2385 928
rect 2346 858 2350 861
rect 2270 752 2273 758
rect 2318 752 2321 798
rect 2326 752 2329 808
rect 2342 772 2345 808
rect 2390 792 2393 928
rect 2406 892 2409 998
rect 2414 792 2417 1028
rect 2438 932 2441 1068
rect 2462 1052 2465 1118
rect 2470 1082 2473 1108
rect 2470 1052 2473 1078
rect 2446 1042 2449 1048
rect 2486 992 2489 1338
rect 2494 1332 2497 1338
rect 2534 1332 2537 1338
rect 2510 1262 2513 1328
rect 2526 1262 2529 1318
rect 2510 1152 2513 1258
rect 2526 1132 2529 1148
rect 2498 1058 2502 1061
rect 2506 1048 2510 1051
rect 2518 992 2521 1028
rect 2454 952 2457 968
rect 2486 952 2489 958
rect 2462 942 2465 948
rect 2442 918 2446 921
rect 2438 872 2441 878
rect 2454 872 2457 938
rect 2470 863 2473 918
rect 2502 892 2505 928
rect 2510 922 2513 958
rect 2534 942 2537 1278
rect 2542 1211 2545 1348
rect 2550 1342 2553 1348
rect 2566 1332 2569 1418
rect 2574 1272 2577 1428
rect 2584 1403 2586 1407
rect 2590 1403 2593 1407
rect 2597 1403 2600 1407
rect 2606 1382 2609 1418
rect 2654 1392 2657 1428
rect 2610 1358 2614 1361
rect 2590 1292 2593 1348
rect 2630 1342 2633 1368
rect 2638 1352 2641 1358
rect 2646 1342 2649 1348
rect 2610 1338 2614 1341
rect 2590 1282 2593 1288
rect 2574 1262 2577 1268
rect 2610 1248 2614 1251
rect 2542 1208 2550 1211
rect 2550 1082 2553 1138
rect 2542 1072 2545 1078
rect 2566 1062 2569 1218
rect 2574 1192 2577 1248
rect 2584 1203 2586 1207
rect 2590 1203 2593 1207
rect 2597 1203 2600 1207
rect 2606 1142 2609 1228
rect 2622 1162 2625 1318
rect 2630 1272 2633 1278
rect 2646 1262 2649 1298
rect 2638 1202 2641 1258
rect 2654 1242 2657 1258
rect 2662 1222 2665 1468
rect 2686 1462 2689 1548
rect 2702 1492 2705 1518
rect 2734 1512 2737 1518
rect 2682 1458 2686 1461
rect 2670 1362 2673 1418
rect 2670 1192 2673 1348
rect 2678 1272 2681 1408
rect 2686 1372 2689 1438
rect 2702 1422 2705 1428
rect 2738 1368 2742 1371
rect 2686 1332 2689 1368
rect 2718 1352 2721 1358
rect 2698 1348 2702 1351
rect 2726 1342 2729 1348
rect 2734 1342 2737 1348
rect 2702 1292 2705 1308
rect 2750 1302 2753 1548
rect 2782 1542 2785 1558
rect 2790 1552 2793 1578
rect 2806 1562 2809 1718
rect 2794 1548 2801 1551
rect 2758 1462 2761 1538
rect 2778 1528 2782 1531
rect 2766 1462 2769 1518
rect 2774 1462 2777 1468
rect 2774 1352 2777 1458
rect 2782 1352 2785 1358
rect 2690 1288 2694 1291
rect 2790 1272 2793 1508
rect 2798 1452 2801 1548
rect 2822 1542 2825 1698
rect 2838 1692 2841 1738
rect 2854 1702 2857 1748
rect 2862 1692 2865 1748
rect 2886 1732 2889 1858
rect 2902 1842 2905 1878
rect 2910 1872 2913 1888
rect 2918 1852 2921 1948
rect 2966 1942 2969 1948
rect 2998 1942 3001 1968
rect 2958 1932 2961 1938
rect 2926 1892 2929 1928
rect 2934 1782 2937 1788
rect 2906 1758 2910 1761
rect 2918 1752 2921 1758
rect 2934 1752 2937 1768
rect 2942 1742 2945 1758
rect 2950 1741 2953 1858
rect 2958 1752 2961 1758
rect 2966 1752 2969 1938
rect 2974 1852 2977 1859
rect 2990 1762 2993 1918
rect 3006 1872 3009 1878
rect 3014 1832 3017 2038
rect 3038 2012 3041 2058
rect 3030 1951 3033 1978
rect 3030 1902 3033 1928
rect 3038 1892 3041 1948
rect 3022 1872 3025 1878
rect 3030 1861 3033 1868
rect 3026 1858 3033 1861
rect 3022 1832 3025 1848
rect 3038 1842 3041 1848
rect 3046 1782 3049 1988
rect 3054 1932 3057 2018
rect 3062 2012 3065 2058
rect 3086 1982 3089 2138
rect 3114 2128 3118 2131
rect 3096 2103 3098 2107
rect 3102 2103 3105 2107
rect 3109 2103 3112 2107
rect 3126 2081 3129 2218
rect 3134 2152 3137 2218
rect 3150 2192 3153 2248
rect 3158 2242 3161 2258
rect 3134 2132 3137 2138
rect 3142 2112 3145 2138
rect 3166 2132 3169 2168
rect 3174 2102 3177 2258
rect 3126 2078 3137 2081
rect 3122 2068 3126 2071
rect 3094 2052 3097 2058
rect 3102 1952 3105 2008
rect 3110 1952 3113 1958
rect 3086 1918 3094 1921
rect 3054 1842 3057 1878
rect 3062 1862 3065 1908
rect 3078 1872 3081 1898
rect 3086 1852 3089 1918
rect 3096 1903 3098 1907
rect 3102 1903 3105 1907
rect 3109 1903 3112 1907
rect 3098 1848 3102 1851
rect 3078 1832 3081 1848
rect 3110 1842 3113 1868
rect 3062 1782 3065 1818
rect 2978 1758 2982 1761
rect 3014 1752 3017 1778
rect 3058 1768 3081 1771
rect 2986 1748 2990 1751
rect 2950 1738 2961 1741
rect 2870 1672 2873 1678
rect 2942 1663 2945 1708
rect 2958 1682 2961 1738
rect 2966 1702 2969 1738
rect 2982 1732 2985 1738
rect 3014 1732 3017 1748
rect 2958 1672 2961 1678
rect 2974 1672 2977 1688
rect 2878 1642 2881 1648
rect 2838 1612 2841 1618
rect 2806 1498 2814 1501
rect 2806 1492 2809 1498
rect 2814 1482 2817 1498
rect 2822 1492 2825 1528
rect 2838 1491 2841 1608
rect 2846 1552 2849 1558
rect 2854 1502 2857 1638
rect 2910 1562 2913 1658
rect 2982 1622 2985 1728
rect 2998 1712 3001 1718
rect 3022 1672 3025 1728
rect 3030 1712 3033 1728
rect 3038 1692 3041 1758
rect 3070 1752 3073 1758
rect 3078 1752 3081 1768
rect 3102 1752 3105 1788
rect 3058 1748 3062 1751
rect 3062 1732 3065 1738
rect 3096 1703 3098 1707
rect 3102 1703 3105 1707
rect 3109 1703 3112 1707
rect 3046 1672 3049 1678
rect 3058 1668 3062 1671
rect 3010 1658 3014 1661
rect 2990 1652 2993 1658
rect 2942 1592 2945 1618
rect 2990 1592 2993 1648
rect 2922 1578 2926 1581
rect 2866 1558 2870 1561
rect 2866 1548 2870 1551
rect 2910 1542 2913 1558
rect 2962 1548 2966 1551
rect 2874 1538 2878 1541
rect 2926 1532 2929 1538
rect 2890 1518 2894 1521
rect 2870 1502 2873 1518
rect 2902 1512 2905 1528
rect 2838 1488 2849 1491
rect 2846 1472 2849 1488
rect 2870 1462 2873 1488
rect 2826 1458 2830 1461
rect 2910 1422 2913 1518
rect 2934 1502 2937 1548
rect 2982 1541 2985 1548
rect 3014 1542 3017 1618
rect 3022 1612 3025 1668
rect 3062 1652 3065 1668
rect 3034 1648 3038 1651
rect 3030 1542 3033 1558
rect 3070 1552 3073 1678
rect 3110 1592 3113 1688
rect 3118 1672 3121 2048
rect 3134 1952 3137 2078
rect 3142 2072 3145 2078
rect 3182 2062 3185 2068
rect 3142 1962 3145 2058
rect 3158 1972 3161 1978
rect 3134 1892 3137 1948
rect 3142 1902 3145 1958
rect 3154 1938 3158 1941
rect 3166 1872 3169 1978
rect 3174 1952 3177 2048
rect 3138 1868 3142 1871
rect 3178 1868 3182 1871
rect 3154 1858 3158 1861
rect 3134 1852 3137 1858
rect 3134 1781 3137 1848
rect 3150 1792 3153 1848
rect 3190 1792 3193 2108
rect 3198 2032 3201 2338
rect 3206 2302 3209 2318
rect 3214 2221 3217 2468
rect 3254 2462 3257 2468
rect 3266 2458 3270 2461
rect 3222 2452 3225 2458
rect 3238 2442 3241 2448
rect 3254 2402 3257 2458
rect 3270 2442 3273 2448
rect 3286 2442 3289 2468
rect 3306 2458 3310 2461
rect 3306 2448 3310 2451
rect 3318 2442 3321 2448
rect 3278 2392 3281 2408
rect 3230 2352 3233 2358
rect 3254 2342 3257 2358
rect 3262 2352 3265 2358
rect 3270 2352 3273 2378
rect 3226 2338 3230 2341
rect 3238 2332 3241 2338
rect 3246 2332 3249 2338
rect 3238 2302 3241 2328
rect 3262 2312 3265 2348
rect 3294 2342 3297 2398
rect 3326 2362 3329 2458
rect 3334 2402 3337 2418
rect 3310 2352 3313 2358
rect 3302 2342 3305 2348
rect 3334 2342 3337 2358
rect 3342 2352 3345 2458
rect 3350 2352 3353 2508
rect 3358 2501 3361 2538
rect 3358 2498 3369 2501
rect 3358 2472 3361 2488
rect 3366 2472 3369 2498
rect 3358 2381 3361 2458
rect 3366 2402 3369 2458
rect 3366 2392 3369 2398
rect 3358 2378 3369 2381
rect 3314 2338 3318 2341
rect 3278 2332 3281 2338
rect 3326 2312 3329 2318
rect 3230 2262 3233 2278
rect 3298 2268 3302 2271
rect 3214 2218 3225 2221
rect 3222 2192 3225 2218
rect 3222 2122 3225 2148
rect 3230 2142 3233 2258
rect 3262 2252 3265 2259
rect 3294 2232 3297 2258
rect 3302 2242 3305 2248
rect 3262 2152 3265 2158
rect 3310 2152 3313 2278
rect 3318 2152 3321 2308
rect 3334 2302 3337 2338
rect 3350 2302 3353 2348
rect 3358 2342 3361 2348
rect 3366 2342 3369 2378
rect 3374 2372 3377 2528
rect 3382 2492 3385 2558
rect 3390 2512 3393 2568
rect 3454 2552 3457 2858
rect 3462 2632 3465 2798
rect 3478 2792 3481 2838
rect 3494 2792 3497 2818
rect 3510 2792 3513 2838
rect 3518 2752 3521 2858
rect 3550 2852 3553 2858
rect 3526 2752 3529 2808
rect 3550 2762 3553 2768
rect 3490 2748 3494 2751
rect 3470 2742 3473 2748
rect 3494 2742 3497 2748
rect 3526 2722 3529 2748
rect 3534 2742 3537 2748
rect 3478 2652 3481 2718
rect 3518 2662 3521 2668
rect 3542 2662 3545 2728
rect 3558 2712 3561 2868
rect 3558 2662 3561 2698
rect 3462 2542 3465 2628
rect 3486 2562 3489 2658
rect 3526 2572 3529 2618
rect 3542 2592 3545 2658
rect 3566 2652 3569 2868
rect 3574 2852 3577 2868
rect 3574 2822 3577 2848
rect 3578 2768 3582 2771
rect 3590 2761 3593 2898
rect 3602 2888 3606 2891
rect 3630 2862 3633 2988
rect 3678 2972 3681 3188
rect 3694 3182 3697 3228
rect 3734 3201 3737 3248
rect 3742 3212 3745 3318
rect 3758 3272 3761 3358
rect 3782 3342 3785 3388
rect 3766 3322 3769 3328
rect 3806 3312 3809 3358
rect 3830 3352 3833 3398
rect 3878 3382 3881 3418
rect 3838 3342 3841 3348
rect 3890 3338 3894 3341
rect 3822 3332 3825 3338
rect 3846 3312 3849 3318
rect 3750 3262 3753 3268
rect 3766 3262 3769 3288
rect 3790 3272 3793 3298
rect 3862 3272 3865 3338
rect 3902 3332 3905 3348
rect 3798 3262 3801 3268
rect 3750 3222 3753 3258
rect 3786 3248 3790 3251
rect 3802 3248 3806 3251
rect 3814 3242 3817 3248
rect 3766 3232 3769 3238
rect 3846 3232 3849 3259
rect 3734 3198 3745 3201
rect 3742 3172 3745 3198
rect 3698 3148 3702 3151
rect 3750 3151 3753 3218
rect 3762 3168 3766 3171
rect 3790 3162 3793 3168
rect 3814 3152 3817 3198
rect 3826 3168 3830 3171
rect 3862 3152 3865 3268
rect 3898 3248 3902 3251
rect 3750 3148 3758 3151
rect 3806 3142 3809 3148
rect 3702 3082 3705 3138
rect 3742 3132 3745 3138
rect 3734 3092 3737 3118
rect 3718 3072 3721 3078
rect 3690 3058 3694 3061
rect 3686 2972 3689 3048
rect 3750 2992 3753 3078
rect 3766 3002 3769 3138
rect 3814 3122 3817 3148
rect 3826 3138 3830 3141
rect 3830 3082 3833 3088
rect 3814 3072 3817 3078
rect 3774 3062 3777 3068
rect 3798 3063 3801 3068
rect 3846 3062 3849 3098
rect 3862 3072 3865 3148
rect 3870 3072 3873 3098
rect 3854 3062 3857 3068
rect 3878 3062 3881 3158
rect 3886 3152 3889 3158
rect 3894 3142 3897 3148
rect 3902 3092 3905 3098
rect 3886 3032 3889 3058
rect 3910 3042 3913 3438
rect 3966 3412 3969 3448
rect 3974 3412 3977 3418
rect 3990 3392 3993 3438
rect 4070 3412 4073 3448
rect 4086 3442 4089 3448
rect 4174 3442 4177 3448
rect 3942 3362 3945 3378
rect 4006 3372 4009 3408
rect 4102 3392 4105 3398
rect 4142 3392 4145 3438
rect 4066 3368 4070 3371
rect 3974 3352 3977 3368
rect 4174 3362 4177 3368
rect 4190 3362 4193 3548
rect 4202 3538 4206 3541
rect 4234 3538 4238 3541
rect 4202 3468 4206 3471
rect 4202 3458 4206 3461
rect 4198 3432 4201 3438
rect 4214 3412 4217 3418
rect 4086 3352 4089 3358
rect 3962 3348 3966 3351
rect 4162 3348 4166 3351
rect 4186 3348 4190 3351
rect 4030 3342 4033 3348
rect 3962 3338 3966 3341
rect 4074 3338 4078 3341
rect 3926 3292 3929 3338
rect 3942 3262 3945 3318
rect 3990 3302 3993 3318
rect 3986 3268 3990 3271
rect 3966 3262 3969 3268
rect 3994 3258 3998 3261
rect 3974 3252 3977 3258
rect 4006 3252 4009 3318
rect 4022 3282 4025 3338
rect 4062 3332 4065 3338
rect 4150 3332 4153 3338
rect 4118 3322 4121 3328
rect 4046 3292 4049 3318
rect 4102 3292 4105 3318
rect 4112 3303 4114 3307
rect 4118 3303 4121 3307
rect 4125 3303 4128 3307
rect 4050 3258 4054 3261
rect 4114 3258 4118 3261
rect 3934 3152 3937 3218
rect 3950 3212 3953 3218
rect 3990 3201 3993 3218
rect 3990 3198 4001 3201
rect 3986 3188 3990 3191
rect 3950 3162 3953 3188
rect 3962 3148 3966 3151
rect 3926 3142 3929 3148
rect 3922 3078 3926 3081
rect 3934 3072 3937 3148
rect 3974 3122 3977 3148
rect 3982 3112 3985 3138
rect 3990 3062 3993 3068
rect 3946 3058 3950 3061
rect 3718 2982 3721 2988
rect 3730 2958 3734 2961
rect 3722 2948 3726 2951
rect 3686 2942 3689 2948
rect 3710 2942 3713 2948
rect 3702 2921 3705 2938
rect 3702 2918 3713 2921
rect 3650 2878 3654 2881
rect 3608 2803 3610 2807
rect 3614 2803 3617 2807
rect 3621 2803 3624 2807
rect 3638 2772 3641 2858
rect 3622 2762 3625 2768
rect 3590 2758 3601 2761
rect 3590 2722 3593 2748
rect 3598 2742 3601 2758
rect 3626 2748 3633 2751
rect 3582 2662 3585 2678
rect 3602 2668 3606 2671
rect 3602 2658 3606 2661
rect 3590 2632 3593 2658
rect 3566 2612 3569 2618
rect 3608 2603 3610 2607
rect 3614 2603 3617 2607
rect 3621 2603 3624 2607
rect 3514 2558 3518 2561
rect 3486 2552 3489 2558
rect 3462 2532 3465 2538
rect 3434 2518 3438 2521
rect 3390 2442 3393 2468
rect 3398 2462 3401 2498
rect 3446 2472 3449 2478
rect 3414 2462 3417 2468
rect 3382 2352 3385 2428
rect 3398 2352 3401 2388
rect 3406 2382 3409 2458
rect 3422 2452 3425 2458
rect 3398 2332 3401 2348
rect 3370 2328 3374 2331
rect 3326 2262 3329 2298
rect 3382 2282 3385 2298
rect 3398 2292 3401 2298
rect 3338 2268 3342 2271
rect 3406 2262 3409 2318
rect 3326 2232 3329 2248
rect 3270 2142 3273 2148
rect 3326 2142 3329 2198
rect 3342 2142 3345 2258
rect 3350 2252 3353 2258
rect 3358 2252 3361 2258
rect 3366 2252 3369 2258
rect 3394 2248 3398 2251
rect 3414 2202 3417 2438
rect 3430 2412 3433 2468
rect 3442 2458 3446 2461
rect 3442 2448 3446 2451
rect 3454 2451 3457 2518
rect 3470 2512 3473 2538
rect 3486 2492 3489 2538
rect 3466 2488 3470 2491
rect 3462 2472 3465 2478
rect 3454 2448 3462 2451
rect 3426 2388 3430 2391
rect 3462 2352 3465 2368
rect 3422 2332 3425 2338
rect 3462 2282 3465 2348
rect 3462 2242 3465 2259
rect 3382 2162 3385 2178
rect 3398 2172 3401 2178
rect 3410 2168 3417 2171
rect 3354 2148 3358 2151
rect 3402 2148 3406 2151
rect 3354 2138 3358 2141
rect 3298 2128 3302 2131
rect 3274 2118 3278 2121
rect 3326 2112 3329 2118
rect 3254 2082 3257 2088
rect 3206 2062 3209 2068
rect 3226 1958 3230 1961
rect 3230 1942 3233 1948
rect 3198 1862 3201 1918
rect 3214 1882 3217 1938
rect 3230 1902 3233 1918
rect 3262 1892 3265 2078
rect 3278 2062 3281 2108
rect 3366 2092 3369 2148
rect 3414 2142 3417 2168
rect 3438 2162 3441 2168
rect 3422 2152 3425 2158
rect 3446 2152 3449 2208
rect 3470 2192 3473 2208
rect 3478 2202 3481 2488
rect 3494 2462 3497 2558
rect 3506 2548 3510 2551
rect 3518 2542 3521 2548
rect 3510 2462 3513 2478
rect 3534 2462 3537 2588
rect 3550 2551 3553 2558
rect 3542 2492 3545 2498
rect 3550 2481 3553 2528
rect 3542 2478 3553 2481
rect 3530 2458 3534 2461
rect 3490 2348 3494 2351
rect 3494 2252 3497 2268
rect 3502 2262 3505 2298
rect 3502 2242 3505 2248
rect 3510 2191 3513 2388
rect 3542 2372 3545 2478
rect 3566 2472 3569 2558
rect 3590 2472 3593 2488
rect 3598 2462 3601 2598
rect 3630 2572 3633 2748
rect 3646 2732 3649 2738
rect 3646 2672 3649 2678
rect 3638 2632 3641 2648
rect 3654 2622 3657 2818
rect 3662 2762 3665 2768
rect 3662 2722 3665 2748
rect 3670 2691 3673 2888
rect 3686 2851 3689 2918
rect 3698 2868 3702 2871
rect 3682 2848 3689 2851
rect 3694 2852 3697 2858
rect 3710 2851 3713 2918
rect 3750 2912 3753 2918
rect 3758 2892 3761 2978
rect 3766 2862 3769 2948
rect 3774 2942 3777 3008
rect 3786 2958 3790 2961
rect 3818 2958 3822 2961
rect 3790 2952 3793 2958
rect 3818 2948 3822 2951
rect 3746 2858 3750 2861
rect 3702 2848 3713 2851
rect 3694 2742 3697 2748
rect 3662 2688 3673 2691
rect 3678 2692 3681 2728
rect 3686 2722 3689 2728
rect 3650 2548 3654 2551
rect 3662 2542 3665 2688
rect 3670 2662 3673 2678
rect 3694 2672 3697 2728
rect 3678 2662 3681 2668
rect 3690 2658 3694 2661
rect 3694 2632 3697 2638
rect 3650 2538 3654 2541
rect 3670 2532 3673 2608
rect 3678 2582 3681 2588
rect 3678 2542 3681 2578
rect 3702 2552 3705 2848
rect 3718 2842 3721 2848
rect 3730 2768 3734 2771
rect 3710 2652 3713 2698
rect 3718 2672 3721 2678
rect 3726 2672 3729 2738
rect 3718 2622 3721 2668
rect 3742 2651 3745 2678
rect 3758 2662 3761 2708
rect 3774 2672 3777 2938
rect 3838 2932 3841 2958
rect 3874 2947 3878 2950
rect 3854 2932 3857 2938
rect 3830 2872 3833 2918
rect 3886 2872 3889 2888
rect 3886 2862 3889 2868
rect 3802 2858 3806 2861
rect 3842 2858 3846 2861
rect 3870 2852 3873 2858
rect 3782 2842 3785 2848
rect 3894 2842 3897 3028
rect 3918 2892 3921 3058
rect 3926 2872 3929 3018
rect 3934 3012 3937 3058
rect 3934 2962 3937 2968
rect 3942 2962 3945 3048
rect 3950 2992 3953 3038
rect 3958 2962 3961 3018
rect 3982 2992 3985 3058
rect 3906 2868 3910 2871
rect 3918 2852 3921 2858
rect 3818 2838 3822 2841
rect 3782 2752 3785 2838
rect 3854 2772 3857 2818
rect 3830 2762 3833 2768
rect 3794 2747 3798 2750
rect 3794 2738 3798 2741
rect 3834 2738 3838 2741
rect 3846 2722 3849 2748
rect 3854 2742 3857 2748
rect 3862 2742 3865 2758
rect 3878 2752 3881 2758
rect 3886 2752 3889 2768
rect 3894 2751 3897 2838
rect 3902 2792 3905 2808
rect 3910 2772 3913 2798
rect 3894 2748 3902 2751
rect 3866 2728 3870 2731
rect 3886 2712 3889 2738
rect 3782 2672 3785 2708
rect 3798 2682 3801 2688
rect 3778 2658 3782 2661
rect 3738 2648 3745 2651
rect 3790 2642 3793 2658
rect 3806 2642 3809 2688
rect 3850 2658 3854 2661
rect 3790 2622 3793 2638
rect 3726 2562 3729 2618
rect 3742 2592 3745 2598
rect 3710 2552 3713 2558
rect 3718 2552 3721 2558
rect 3750 2552 3753 2608
rect 3774 2562 3777 2578
rect 3790 2552 3793 2598
rect 3690 2548 3694 2551
rect 3690 2538 3694 2541
rect 3662 2511 3665 2518
rect 3654 2508 3665 2511
rect 3626 2458 3630 2461
rect 3550 2452 3553 2458
rect 3578 2448 3582 2451
rect 3526 2332 3529 2348
rect 3526 2252 3529 2308
rect 3534 2212 3537 2348
rect 3542 2332 3545 2338
rect 3550 2331 3553 2448
rect 3558 2352 3561 2438
rect 3582 2412 3585 2418
rect 3550 2328 3561 2331
rect 3542 2272 3545 2298
rect 3558 2292 3561 2328
rect 3574 2302 3577 2348
rect 3550 2262 3553 2278
rect 3566 2262 3569 2298
rect 3574 2282 3577 2298
rect 3562 2228 3566 2231
rect 3574 2212 3577 2258
rect 3510 2188 3521 2191
rect 3478 2152 3481 2158
rect 3510 2152 3513 2158
rect 3422 2122 3425 2138
rect 3446 2092 3449 2138
rect 3290 2088 3294 2091
rect 3382 2082 3385 2088
rect 3418 2068 3422 2071
rect 3442 2068 3446 2071
rect 3334 2062 3337 2068
rect 3282 2058 3289 2061
rect 3274 2048 3278 2051
rect 3198 1792 3201 1838
rect 3134 1778 3145 1781
rect 3126 1732 3129 1778
rect 3134 1742 3137 1748
rect 3126 1682 3129 1728
rect 3142 1712 3145 1778
rect 3170 1748 3174 1751
rect 3218 1748 3222 1751
rect 3206 1732 3209 1748
rect 3230 1732 3233 1868
rect 3242 1858 3246 1861
rect 3274 1788 3278 1791
rect 3270 1752 3273 1758
rect 3238 1742 3241 1748
rect 3266 1738 3270 1741
rect 3170 1728 3177 1731
rect 3118 1582 3121 1658
rect 3046 1542 3049 1548
rect 3070 1542 3073 1548
rect 2982 1538 2993 1541
rect 2950 1522 2953 1528
rect 2958 1512 2961 1528
rect 2970 1488 2974 1491
rect 2926 1471 2929 1488
rect 2934 1472 2937 1478
rect 2926 1468 2934 1471
rect 2974 1462 2977 1468
rect 2954 1458 2958 1461
rect 2982 1452 2985 1458
rect 2822 1272 2825 1368
rect 2866 1358 2870 1361
rect 2886 1352 2889 1358
rect 2842 1348 2846 1351
rect 2858 1348 2862 1351
rect 2870 1342 2873 1348
rect 2842 1338 2846 1341
rect 2878 1322 2881 1338
rect 2894 1332 2897 1418
rect 2838 1292 2841 1308
rect 2638 1152 2641 1168
rect 2654 1142 2657 1168
rect 2542 992 2545 998
rect 2550 982 2553 1058
rect 2566 1052 2569 1058
rect 2558 952 2561 1018
rect 2566 962 2569 1038
rect 2574 962 2577 1118
rect 2606 1092 2609 1118
rect 2622 1112 2625 1118
rect 2614 1078 2633 1081
rect 2590 1062 2593 1068
rect 2614 1062 2617 1078
rect 2630 1072 2633 1078
rect 2622 1062 2625 1068
rect 2630 1052 2633 1058
rect 2584 1003 2586 1007
rect 2590 1003 2593 1007
rect 2597 1003 2600 1007
rect 2566 952 2569 958
rect 2614 952 2617 1048
rect 2638 992 2641 1138
rect 2654 1092 2657 1138
rect 2662 1112 2665 1148
rect 2678 1142 2681 1258
rect 2750 1252 2753 1258
rect 2710 1192 2713 1238
rect 2730 1168 2734 1171
rect 2718 1158 2726 1161
rect 2694 1152 2697 1158
rect 2706 1148 2710 1151
rect 2686 1122 2689 1148
rect 2702 1132 2705 1138
rect 2718 1092 2721 1158
rect 2766 1152 2769 1208
rect 2774 1152 2777 1268
rect 2790 1262 2793 1268
rect 2806 1262 2809 1268
rect 2846 1262 2849 1268
rect 2838 1242 2841 1248
rect 2782 1152 2785 1158
rect 2798 1152 2801 1198
rect 2846 1152 2849 1158
rect 2862 1152 2865 1218
rect 2766 1142 2769 1148
rect 2742 1091 2745 1128
rect 2750 1122 2753 1128
rect 2738 1088 2745 1091
rect 2702 1072 2705 1088
rect 2774 1082 2777 1148
rect 2786 1138 2790 1141
rect 2774 1072 2777 1078
rect 2722 1068 2726 1071
rect 2662 1062 2665 1068
rect 2670 1062 2673 1068
rect 2682 1058 2686 1061
rect 2786 1058 2790 1061
rect 2694 1052 2697 1058
rect 2678 1032 2681 1048
rect 2658 948 2662 951
rect 2534 922 2537 938
rect 2530 888 2534 891
rect 2454 792 2457 848
rect 2558 842 2561 948
rect 2574 872 2577 938
rect 2582 902 2585 918
rect 2566 852 2569 858
rect 2598 852 2601 868
rect 2366 762 2369 768
rect 2290 748 2294 751
rect 2318 742 2321 748
rect 2366 742 2369 748
rect 2374 742 2377 788
rect 2414 752 2417 758
rect 2138 668 2142 671
rect 2142 542 2145 668
rect 2150 652 2153 658
rect 2166 652 2169 658
rect 2182 651 2185 668
rect 2222 652 2225 659
rect 2178 648 2185 651
rect 2190 572 2193 648
rect 2238 592 2241 738
rect 2262 712 2265 738
rect 2306 728 2310 731
rect 2286 682 2289 688
rect 2318 672 2321 718
rect 2334 692 2337 698
rect 2358 692 2361 718
rect 2374 692 2377 708
rect 2354 678 2358 681
rect 2346 668 2350 671
rect 2294 662 2297 668
rect 2218 568 2222 571
rect 2158 542 2161 558
rect 2170 548 2174 551
rect 2054 532 2057 538
rect 2072 503 2074 507
rect 2078 503 2081 507
rect 2085 503 2088 507
rect 2022 462 2025 468
rect 2038 452 2041 488
rect 2054 462 2057 468
rect 2062 462 2065 498
rect 2070 472 2073 478
rect 1918 358 1926 361
rect 1910 352 1913 358
rect 1838 342 1841 348
rect 1822 308 1833 311
rect 1806 272 1809 288
rect 1754 268 1761 271
rect 1802 268 1806 271
rect 1722 238 1726 241
rect 1686 172 1689 228
rect 1750 192 1753 268
rect 1794 258 1798 261
rect 1758 222 1761 258
rect 1802 248 1806 251
rect 1774 242 1777 248
rect 1810 238 1814 241
rect 1706 168 1710 171
rect 1766 162 1769 168
rect 1722 158 1726 161
rect 1738 158 1742 161
rect 1754 158 1758 161
rect 1778 158 1785 161
rect 1646 152 1649 158
rect 1714 148 1718 151
rect 1754 148 1758 151
rect 1706 138 1710 141
rect 1742 132 1745 138
rect 1598 82 1601 88
rect 1614 72 1617 78
rect 1638 72 1641 128
rect 1690 88 1694 91
rect 1706 88 1710 91
rect 1582 62 1585 68
rect 1766 63 1769 118
rect 1774 102 1777 118
rect 1782 102 1785 158
rect 1790 152 1793 198
rect 1822 152 1825 268
rect 1830 192 1833 308
rect 1846 262 1849 338
rect 1870 282 1873 348
rect 1890 328 1897 331
rect 1846 232 1849 258
rect 1846 162 1849 198
rect 1854 142 1857 278
rect 1870 252 1873 258
rect 1894 182 1897 328
rect 1918 292 1921 358
rect 1942 332 1945 338
rect 1926 272 1929 278
rect 1958 272 1961 288
rect 1938 268 1942 271
rect 1966 262 1969 388
rect 1974 352 1977 368
rect 1990 342 1993 418
rect 1982 262 1985 268
rect 1954 248 1958 251
rect 1910 242 1913 248
rect 1990 242 1993 248
rect 1942 202 1945 218
rect 1914 178 1918 181
rect 1886 172 1889 178
rect 1862 152 1865 158
rect 1878 142 1881 158
rect 1950 152 1953 228
rect 1906 148 1910 151
rect 1802 138 1806 141
rect 1906 138 1910 141
rect 1802 128 1806 131
rect 1798 92 1801 98
rect 1538 58 1542 61
rect 1570 58 1574 61
rect 1634 59 1638 62
rect 1782 62 1785 68
rect 1814 62 1817 78
rect 1822 72 1825 118
rect 1910 72 1913 78
rect 1958 72 1961 208
rect 2006 171 2009 398
rect 2054 382 2057 408
rect 2026 378 2030 381
rect 2054 372 2057 378
rect 2038 342 2041 348
rect 2026 338 2030 341
rect 2014 312 2017 328
rect 2014 272 2017 308
rect 2014 222 2017 258
rect 2022 242 2025 248
rect 2030 192 2033 338
rect 1998 168 2009 171
rect 1974 152 1977 158
rect 1998 112 2001 168
rect 1990 92 1993 98
rect 1830 62 1833 68
rect 1894 62 1897 68
rect 1934 62 1937 68
rect 1998 62 2001 108
rect 2014 82 2017 88
rect 2022 62 2025 68
rect 1798 52 1801 58
rect 2030 52 2033 108
rect 2038 92 2041 338
rect 2054 212 2057 258
rect 2050 148 2054 151
rect 2046 62 2049 78
rect 2062 71 2065 358
rect 2086 351 2089 428
rect 2094 372 2097 378
rect 2086 348 2094 351
rect 2072 303 2074 307
rect 2078 303 2081 307
rect 2085 303 2088 307
rect 2094 302 2097 348
rect 2102 342 2105 498
rect 2126 482 2129 538
rect 2118 463 2121 468
rect 2110 392 2113 418
rect 2126 382 2129 478
rect 2134 342 2137 348
rect 2142 342 2145 538
rect 2206 492 2209 558
rect 2246 552 2249 588
rect 2310 562 2313 658
rect 2318 592 2321 668
rect 2366 652 2369 668
rect 2374 662 2377 688
rect 2382 662 2385 728
rect 2390 692 2393 728
rect 2398 722 2401 738
rect 2406 722 2409 748
rect 2430 742 2433 758
rect 2478 752 2481 798
rect 2486 792 2489 808
rect 2518 752 2521 838
rect 2550 792 2553 818
rect 2584 803 2586 807
rect 2590 803 2593 807
rect 2597 803 2600 807
rect 2542 752 2545 768
rect 2414 692 2417 738
rect 2330 648 2334 651
rect 2334 562 2337 598
rect 2350 592 2353 648
rect 2382 562 2385 658
rect 2302 552 2305 558
rect 2310 552 2313 558
rect 2266 548 2270 551
rect 2330 548 2334 551
rect 2278 542 2281 548
rect 2306 538 2310 541
rect 2178 488 2182 491
rect 2150 462 2153 468
rect 2190 402 2193 458
rect 2230 441 2233 528
rect 2254 462 2257 478
rect 2262 462 2265 468
rect 2222 438 2233 441
rect 2154 368 2158 371
rect 2174 352 2177 388
rect 2178 338 2182 341
rect 2126 332 2129 338
rect 2074 258 2078 261
rect 2118 192 2121 328
rect 2134 312 2137 338
rect 2162 318 2166 321
rect 2198 321 2201 338
rect 2190 318 2201 321
rect 2214 322 2217 347
rect 2190 282 2193 318
rect 2190 272 2193 278
rect 2170 258 2174 261
rect 2150 168 2169 171
rect 2102 162 2105 168
rect 2150 162 2153 168
rect 2126 158 2134 161
rect 2126 152 2129 158
rect 2158 152 2161 158
rect 2166 152 2169 168
rect 2174 152 2177 218
rect 2138 148 2142 151
rect 2182 142 2185 268
rect 2206 182 2209 298
rect 2194 158 2201 161
rect 2198 142 2201 158
rect 2206 152 2209 178
rect 2214 152 2217 288
rect 2222 242 2225 438
rect 2262 372 2265 458
rect 2270 442 2273 538
rect 2306 528 2310 531
rect 2310 492 2313 508
rect 2310 452 2313 488
rect 2318 472 2321 518
rect 2230 272 2233 288
rect 2238 262 2241 318
rect 2270 292 2273 438
rect 2318 402 2321 468
rect 2326 462 2329 518
rect 2342 512 2345 528
rect 2334 472 2337 478
rect 2342 468 2350 471
rect 2330 458 2337 461
rect 2278 372 2281 378
rect 2286 362 2289 368
rect 2302 352 2305 388
rect 2318 362 2321 398
rect 2326 362 2329 368
rect 2318 352 2321 358
rect 2318 332 2321 338
rect 2230 258 2238 261
rect 2250 258 2254 261
rect 2230 252 2233 258
rect 2262 242 2265 248
rect 2226 238 2230 241
rect 2222 162 2225 168
rect 2238 152 2241 218
rect 2122 138 2126 141
rect 2190 132 2193 138
rect 2072 103 2074 107
rect 2078 103 2081 107
rect 2085 103 2088 107
rect 2058 68 2065 71
rect 2070 61 2073 88
rect 2066 58 2073 61
rect 2102 72 2105 108
rect 2174 72 2177 108
rect 2206 82 2209 148
rect 2214 142 2217 148
rect 2222 142 2225 148
rect 2246 142 2249 188
rect 2254 172 2257 228
rect 2278 162 2281 308
rect 2286 302 2289 318
rect 2326 312 2329 348
rect 2334 322 2337 458
rect 2342 452 2345 468
rect 2366 462 2369 558
rect 2382 532 2385 538
rect 2382 472 2385 528
rect 2390 492 2393 648
rect 2398 582 2401 668
rect 2414 602 2417 638
rect 2422 632 2425 668
rect 2398 532 2401 548
rect 2430 522 2433 658
rect 2438 581 2441 748
rect 2446 681 2449 748
rect 2470 732 2473 748
rect 2446 678 2457 681
rect 2454 672 2457 678
rect 2446 662 2449 668
rect 2462 662 2465 678
rect 2458 658 2462 661
rect 2478 652 2481 688
rect 2518 672 2521 748
rect 2590 732 2593 738
rect 2598 702 2601 758
rect 2570 688 2574 691
rect 2606 672 2609 948
rect 2622 942 2625 948
rect 2646 942 2649 948
rect 2618 888 2622 891
rect 2630 862 2633 908
rect 2646 882 2649 888
rect 2646 872 2649 878
rect 2614 792 2617 848
rect 2614 752 2617 758
rect 2622 752 2625 858
rect 2638 802 2641 868
rect 2662 852 2665 858
rect 2670 832 2673 838
rect 2678 792 2681 998
rect 2686 882 2689 938
rect 2698 888 2702 891
rect 2686 852 2689 868
rect 2694 862 2697 868
rect 2694 792 2697 828
rect 2654 762 2657 768
rect 2618 738 2622 741
rect 2646 722 2649 728
rect 2510 663 2513 668
rect 2614 662 2617 668
rect 2622 652 2625 668
rect 2450 648 2454 651
rect 2466 648 2470 651
rect 2598 632 2601 648
rect 2446 592 2449 598
rect 2438 578 2449 581
rect 2446 472 2449 578
rect 2462 552 2465 628
rect 2478 562 2481 568
rect 2474 548 2478 551
rect 2454 491 2457 538
rect 2462 502 2465 548
rect 2514 547 2518 550
rect 2494 532 2497 538
rect 2566 512 2569 628
rect 2574 592 2577 618
rect 2584 603 2586 607
rect 2590 603 2593 607
rect 2597 603 2600 607
rect 2606 591 2609 648
rect 2630 642 2633 698
rect 2646 662 2649 678
rect 2654 672 2657 678
rect 2662 672 2665 788
rect 2678 752 2681 788
rect 2710 782 2713 1048
rect 2766 1032 2769 1058
rect 2750 992 2753 1028
rect 2798 1002 2801 1148
rect 2838 1142 2841 1148
rect 2806 1122 2809 1128
rect 2862 1092 2865 1148
rect 2830 1072 2833 1078
rect 2854 1062 2857 1068
rect 2862 1062 2865 1068
rect 2830 1002 2833 1058
rect 2838 972 2841 1048
rect 2870 972 2873 1298
rect 2902 1282 2905 1348
rect 2910 1342 2913 1398
rect 2966 1392 2969 1438
rect 2990 1432 2993 1538
rect 3018 1528 3022 1531
rect 3042 1528 3054 1531
rect 2998 1522 3001 1528
rect 3006 1512 3009 1528
rect 3070 1522 3073 1538
rect 3006 1492 3009 1508
rect 3030 1492 3033 1508
rect 3046 1482 3049 1488
rect 3042 1468 3046 1471
rect 3014 1451 3017 1468
rect 3026 1458 3033 1461
rect 3014 1448 3022 1451
rect 3030 1442 3033 1458
rect 2926 1382 2929 1388
rect 2934 1352 2937 1388
rect 2958 1372 2961 1378
rect 2942 1352 2945 1358
rect 2926 1332 2929 1338
rect 2878 1262 2881 1268
rect 2898 1258 2902 1261
rect 2894 1172 2897 1218
rect 2910 1212 2913 1328
rect 2950 1312 2953 1348
rect 2998 1302 3001 1418
rect 3006 1352 3009 1358
rect 2926 1282 2929 1288
rect 3006 1272 3009 1338
rect 2946 1268 2950 1271
rect 2986 1268 2990 1271
rect 2978 1258 2982 1261
rect 2910 1192 2913 1208
rect 2902 1142 2905 1158
rect 2926 1152 2929 1258
rect 2990 1252 2993 1258
rect 2946 1148 2950 1151
rect 2878 1082 2881 1108
rect 2870 961 2873 968
rect 2862 958 2873 961
rect 2798 932 2801 948
rect 2806 872 2809 938
rect 2758 842 2761 858
rect 2726 751 2729 758
rect 2670 742 2673 748
rect 2710 732 2713 738
rect 2686 692 2689 728
rect 2726 672 2729 728
rect 2782 692 2785 828
rect 2822 792 2825 958
rect 2862 952 2865 958
rect 2918 952 2921 1138
rect 2926 1072 2929 1148
rect 2934 1102 2937 1148
rect 2958 1142 2961 1248
rect 3006 1241 3009 1268
rect 3022 1252 3025 1259
rect 2998 1238 3009 1241
rect 2998 1162 3001 1238
rect 3054 1232 3057 1448
rect 3062 1382 3065 1518
rect 3074 1468 3078 1471
rect 3070 1392 3073 1408
rect 3062 1362 3065 1368
rect 3078 1332 3081 1358
rect 2966 1142 2969 1148
rect 2998 1142 3001 1158
rect 3018 1147 3022 1150
rect 2942 1132 2945 1138
rect 2982 1132 2985 1138
rect 3046 1132 3049 1138
rect 2934 1082 2937 1098
rect 2938 1058 2942 1061
rect 2926 1052 2929 1058
rect 2942 992 2945 1048
rect 2982 992 2985 1118
rect 2994 1088 2998 1091
rect 3006 1062 3009 1068
rect 3038 1062 3041 1068
rect 3070 1062 3073 1078
rect 3078 1052 3081 1058
rect 3022 1012 3025 1018
rect 2926 952 2929 958
rect 2958 952 2961 958
rect 2966 952 2969 978
rect 3022 962 3025 1008
rect 3054 992 3057 1018
rect 2870 942 2873 948
rect 2854 922 2857 938
rect 2894 932 2897 938
rect 2878 922 2881 928
rect 2830 862 2833 878
rect 2846 832 2849 858
rect 2854 792 2857 898
rect 2890 888 2894 891
rect 2910 872 2913 878
rect 2890 868 2894 871
rect 2898 858 2902 861
rect 2798 752 2801 758
rect 2862 752 2865 808
rect 2894 792 2897 798
rect 2902 752 2905 858
rect 2918 852 2921 948
rect 2950 902 2953 948
rect 2974 932 2977 948
rect 2962 878 2966 881
rect 2926 852 2929 878
rect 2954 868 2958 871
rect 2982 862 2985 928
rect 2998 892 3001 948
rect 3014 942 3017 958
rect 3074 948 3078 951
rect 3030 942 3033 948
rect 3018 918 3022 921
rect 3062 872 3065 928
rect 2806 742 2809 748
rect 2790 722 2793 728
rect 2602 588 2609 591
rect 2614 592 2617 628
rect 2630 622 2633 638
rect 2638 562 2641 658
rect 2502 492 2505 508
rect 2454 488 2465 491
rect 2462 472 2465 488
rect 2510 472 2513 478
rect 2402 468 2406 471
rect 2426 468 2430 471
rect 2350 452 2353 458
rect 2374 442 2377 468
rect 2434 458 2438 461
rect 2382 442 2385 448
rect 2342 372 2345 418
rect 2342 322 2345 348
rect 2350 342 2353 408
rect 2362 388 2366 391
rect 2374 381 2377 438
rect 2406 422 2409 448
rect 2414 442 2417 448
rect 2374 378 2385 381
rect 2374 362 2377 368
rect 2354 338 2358 341
rect 2374 322 2377 348
rect 2382 342 2385 378
rect 2390 362 2393 368
rect 2374 312 2377 318
rect 2382 312 2385 338
rect 2286 272 2289 288
rect 2302 272 2305 278
rect 2318 263 2321 298
rect 2386 288 2390 291
rect 2386 268 2390 271
rect 2398 262 2401 318
rect 2406 292 2409 418
rect 2422 392 2425 458
rect 2438 432 2441 458
rect 2450 448 2454 451
rect 2414 362 2417 368
rect 2414 292 2417 328
rect 2286 222 2289 258
rect 2414 252 2417 288
rect 2438 262 2441 398
rect 2454 351 2457 388
rect 2450 288 2454 291
rect 2462 282 2465 468
rect 2494 462 2497 468
rect 2542 463 2545 468
rect 2470 412 2473 458
rect 2486 452 2489 458
rect 2550 452 2553 468
rect 2494 442 2497 448
rect 2514 368 2518 371
rect 2446 272 2449 278
rect 2486 272 2489 348
rect 2550 332 2553 448
rect 2584 403 2586 407
rect 2590 403 2593 407
rect 2597 403 2600 407
rect 2606 372 2609 528
rect 2622 492 2625 528
rect 2630 462 2633 518
rect 2646 462 2649 658
rect 2662 492 2665 658
rect 2682 648 2686 651
rect 2718 632 2721 659
rect 2790 652 2793 668
rect 2802 658 2806 661
rect 2670 622 2673 628
rect 2694 551 2697 558
rect 2786 548 2793 551
rect 2802 548 2806 551
rect 2742 542 2745 548
rect 2750 542 2753 548
rect 2770 538 2774 541
rect 2654 472 2657 478
rect 2666 468 2670 471
rect 2678 462 2681 528
rect 2694 472 2697 528
rect 2726 522 2729 528
rect 2618 458 2622 461
rect 2678 452 2681 458
rect 2694 452 2697 468
rect 2722 458 2726 461
rect 2618 388 2622 391
rect 2558 352 2561 358
rect 2654 352 2657 398
rect 2662 392 2665 438
rect 2670 361 2673 418
rect 2694 362 2697 368
rect 2670 358 2678 361
rect 2714 358 2718 361
rect 2734 352 2737 388
rect 2690 348 2694 351
rect 2686 332 2689 338
rect 2550 272 2553 328
rect 2638 292 2641 328
rect 2650 288 2654 291
rect 2686 272 2689 308
rect 2438 242 2441 248
rect 2366 191 2369 238
rect 2446 212 2449 268
rect 2710 262 2713 348
rect 2742 342 2745 408
rect 2758 392 2761 528
rect 2782 482 2785 528
rect 2790 471 2793 548
rect 2814 482 2817 668
rect 2822 662 2825 678
rect 2822 492 2825 558
rect 2830 552 2833 748
rect 2846 702 2849 728
rect 2854 662 2857 678
rect 2838 592 2841 618
rect 2870 592 2873 618
rect 2838 562 2841 588
rect 2830 522 2833 538
rect 2878 502 2881 718
rect 2906 668 2910 671
rect 2886 652 2889 658
rect 2886 592 2889 608
rect 2902 532 2905 648
rect 2918 552 2921 848
rect 2942 782 2945 858
rect 2982 842 2985 858
rect 2990 848 2998 851
rect 2926 762 2929 768
rect 2958 742 2961 828
rect 2934 672 2937 678
rect 2942 662 2945 698
rect 2930 658 2934 661
rect 2950 652 2953 658
rect 2930 648 2934 651
rect 2958 612 2961 738
rect 2966 692 2969 788
rect 2974 751 2977 758
rect 2990 692 2993 848
rect 3014 832 3017 868
rect 3038 852 3041 858
rect 3086 792 3089 1548
rect 3096 1503 3098 1507
rect 3102 1503 3105 1507
rect 3109 1503 3112 1507
rect 3118 1502 3121 1578
rect 3126 1552 3129 1578
rect 3134 1552 3137 1618
rect 3142 1512 3145 1708
rect 3174 1702 3177 1728
rect 3222 1722 3225 1728
rect 3158 1682 3161 1688
rect 3166 1672 3169 1688
rect 3174 1661 3177 1698
rect 3182 1692 3185 1718
rect 3190 1692 3193 1718
rect 3170 1658 3177 1661
rect 3222 1652 3225 1658
rect 3230 1651 3233 1728
rect 3246 1662 3249 1738
rect 3226 1648 3233 1651
rect 3162 1578 3166 1581
rect 3174 1552 3177 1578
rect 3182 1552 3185 1608
rect 3206 1592 3209 1598
rect 3154 1548 3158 1551
rect 3190 1542 3193 1558
rect 3206 1552 3209 1558
rect 3214 1542 3217 1608
rect 3230 1542 3233 1648
rect 3270 1642 3273 1718
rect 3286 1702 3289 2058
rect 3398 2062 3401 2068
rect 3314 1947 3318 1950
rect 3334 1942 3337 2058
rect 3350 2042 3353 2059
rect 3442 2058 3446 2061
rect 3410 2038 3414 2041
rect 3430 2032 3433 2058
rect 3446 1992 3449 2038
rect 3454 1962 3457 2148
rect 3462 2072 3465 2108
rect 3486 2092 3489 2148
rect 3494 2142 3497 2148
rect 3502 2092 3505 2108
rect 3482 2068 3486 2071
rect 3462 2052 3465 2068
rect 3518 2062 3521 2188
rect 3550 2132 3553 2148
rect 3574 2132 3577 2158
rect 3526 2112 3529 2128
rect 3550 2092 3553 2128
rect 3474 2058 3478 2061
rect 3498 2048 3502 2051
rect 3354 1958 3358 1961
rect 3406 1952 3409 1958
rect 3478 1952 3481 2008
rect 3486 1952 3489 1978
rect 3378 1948 3382 1951
rect 3434 1948 3438 1951
rect 3334 1912 3337 1938
rect 3358 1932 3361 1948
rect 3366 1942 3369 1948
rect 3422 1942 3425 1948
rect 3462 1942 3465 1948
rect 3378 1938 3382 1941
rect 3390 1932 3393 1938
rect 3350 1891 3353 1918
rect 3342 1888 3353 1891
rect 3310 1732 3313 1748
rect 3318 1681 3321 1858
rect 3326 1852 3329 1858
rect 3334 1852 3337 1858
rect 3342 1852 3345 1888
rect 3358 1872 3361 1908
rect 3438 1892 3441 1898
rect 3342 1751 3345 1758
rect 3358 1742 3361 1868
rect 3386 1858 3390 1861
rect 3470 1852 3473 1948
rect 3478 1862 3481 1908
rect 3486 1792 3489 1928
rect 3494 1872 3497 2028
rect 3510 1952 3513 1958
rect 3518 1952 3521 2058
rect 3502 1942 3505 1948
rect 3502 1852 3505 1858
rect 3374 1742 3377 1748
rect 3382 1731 3385 1778
rect 3398 1752 3401 1758
rect 3378 1728 3385 1731
rect 3390 1722 3393 1738
rect 3406 1732 3409 1788
rect 3518 1782 3521 1948
rect 3534 1932 3537 1938
rect 3542 1932 3545 2048
rect 3558 2022 3561 2118
rect 3566 2063 3569 2118
rect 3582 2052 3585 2348
rect 3598 2332 3601 2448
rect 3654 2442 3657 2508
rect 3666 2498 3673 2501
rect 3670 2463 3673 2498
rect 3634 2438 3638 2441
rect 3608 2403 3610 2407
rect 3614 2403 3617 2407
rect 3621 2403 3624 2407
rect 3638 2362 3641 2418
rect 3634 2348 3638 2351
rect 3602 2328 3606 2331
rect 3622 2312 3625 2318
rect 3630 2302 3633 2338
rect 3646 2322 3649 2328
rect 3630 2282 3633 2298
rect 3662 2292 3665 2418
rect 3678 2372 3681 2468
rect 3702 2462 3705 2548
rect 3774 2542 3777 2548
rect 3746 2538 3750 2541
rect 3758 2531 3761 2538
rect 3750 2528 3761 2531
rect 3742 2492 3745 2498
rect 3702 2312 3705 2348
rect 3678 2272 3681 2298
rect 3590 2262 3593 2268
rect 3608 2203 3610 2207
rect 3614 2203 3617 2207
rect 3621 2203 3624 2207
rect 3630 2172 3633 2178
rect 3590 2142 3593 2158
rect 3610 2148 3614 2151
rect 3622 2142 3625 2148
rect 3638 2142 3641 2258
rect 3646 2252 3649 2258
rect 3702 2222 3705 2238
rect 3646 2152 3649 2158
rect 3654 2152 3657 2188
rect 3670 2152 3673 2188
rect 3678 2152 3681 2168
rect 3690 2148 3694 2151
rect 3646 2062 3649 2128
rect 3702 2112 3705 2218
rect 3710 2171 3713 2328
rect 3726 2272 3729 2448
rect 3734 2442 3737 2448
rect 3742 2392 3745 2448
rect 3742 2362 3745 2378
rect 3750 2362 3753 2528
rect 3766 2492 3769 2518
rect 3806 2492 3809 2588
rect 3814 2562 3817 2598
rect 3862 2582 3865 2668
rect 3894 2662 3897 2678
rect 3902 2652 3905 2748
rect 3910 2722 3913 2748
rect 3926 2742 3929 2858
rect 3942 2852 3945 2958
rect 3974 2952 3977 2988
rect 3998 2952 4001 3198
rect 4006 3142 4009 3168
rect 4014 3062 4017 3068
rect 4022 3062 4025 3248
rect 4030 3072 4033 3078
rect 4038 3062 4041 3178
rect 4046 3152 4049 3158
rect 4070 3142 4073 3258
rect 4054 3091 4057 3128
rect 4054 3088 4065 3091
rect 4062 3072 4065 3088
rect 4050 3068 4054 3071
rect 4086 3062 4089 3068
rect 4026 3058 4030 3061
rect 3962 2948 3966 2951
rect 3950 2852 3953 2918
rect 3958 2882 3961 2938
rect 4006 2912 4009 3018
rect 4054 2992 4057 3008
rect 4022 2982 4025 2988
rect 4086 2982 4089 3038
rect 4066 2948 4070 2951
rect 3934 2832 3937 2838
rect 3946 2758 3953 2761
rect 3950 2752 3953 2758
rect 3938 2748 3942 2751
rect 3958 2742 3961 2868
rect 3966 2862 3969 2908
rect 4022 2892 4025 2908
rect 4038 2892 4041 2948
rect 4094 2942 4097 3128
rect 4110 3121 4113 3248
rect 4134 3152 4137 3298
rect 4142 3281 4145 3318
rect 4142 3278 4153 3281
rect 4150 3272 4153 3278
rect 4158 3272 4161 3328
rect 4198 3322 4201 3348
rect 4206 3342 4209 3378
rect 4222 3361 4225 3518
rect 4254 3442 4257 3458
rect 4262 3382 4265 3658
rect 4278 3482 4281 3538
rect 4218 3358 4225 3361
rect 4258 3348 4262 3351
rect 4226 3338 4230 3341
rect 4246 3332 4249 3348
rect 4258 3338 4262 3341
rect 4230 3328 4238 3331
rect 4214 3292 4217 3318
rect 4230 3282 4233 3328
rect 4246 3302 4249 3318
rect 4206 3272 4209 3278
rect 4214 3272 4217 3278
rect 4142 3262 4145 3268
rect 4158 3262 4161 3268
rect 4174 3242 4177 3268
rect 4238 3262 4241 3268
rect 4202 3248 4206 3251
rect 4214 3242 4217 3258
rect 4174 3202 4177 3238
rect 4230 3222 4233 3258
rect 4246 3252 4249 3258
rect 4254 3222 4257 3338
rect 4286 3282 4289 3308
rect 4294 3261 4297 3738
rect 4334 3722 4337 3738
rect 4342 3702 4345 3748
rect 4358 3742 4361 3818
rect 4366 3762 4369 3768
rect 4382 3742 4385 3808
rect 4422 3761 4425 3818
rect 4446 3812 4449 3858
rect 4506 3848 4510 3851
rect 4414 3758 4425 3761
rect 4402 3748 4406 3751
rect 4382 3702 4385 3738
rect 4390 3732 4393 3738
rect 4358 3672 4361 3678
rect 4302 3552 4305 3558
rect 4310 3542 4313 3658
rect 4318 3652 4321 3658
rect 4374 3652 4377 3658
rect 4358 3571 4361 3628
rect 4350 3568 4361 3571
rect 4342 3542 4345 3548
rect 4350 3462 4353 3568
rect 4358 3552 4361 3558
rect 4358 3462 4361 3468
rect 4310 3422 4313 3458
rect 4318 3432 4321 3458
rect 4302 3332 4305 3348
rect 4290 3258 4297 3261
rect 4190 3192 4193 3198
rect 4158 3152 4161 3178
rect 4198 3152 4201 3168
rect 4102 3118 4113 3121
rect 4102 3092 4105 3118
rect 4112 3103 4114 3107
rect 4118 3103 4121 3107
rect 4125 3103 4128 3107
rect 4106 3048 4110 3051
rect 4134 2972 4137 3128
rect 4158 3072 4161 3148
rect 4206 3142 4209 3158
rect 4246 3152 4249 3158
rect 4262 3152 4265 3218
rect 4294 3161 4297 3218
rect 4302 3212 4305 3218
rect 4310 3192 4313 3338
rect 4326 3301 4329 3418
rect 4358 3392 4361 3458
rect 4354 3368 4358 3371
rect 4366 3352 4369 3608
rect 4390 3592 4393 3618
rect 4398 3592 4401 3718
rect 4414 3662 4417 3758
rect 4454 3752 4457 3848
rect 4462 3792 4465 3848
rect 4422 3722 4425 3748
rect 4406 3642 4409 3658
rect 4422 3582 4425 3618
rect 4430 3571 4433 3748
rect 4438 3712 4441 3738
rect 4442 3658 4446 3661
rect 4454 3652 4457 3668
rect 4470 3662 4473 3788
rect 4490 3658 4494 3661
rect 4470 3652 4473 3658
rect 4494 3642 4497 3648
rect 4510 3572 4513 3618
rect 4426 3568 4433 3571
rect 4382 3562 4385 3568
rect 4386 3548 4390 3551
rect 4390 3472 4393 3528
rect 4374 3341 4377 3418
rect 4390 3402 4393 3468
rect 4398 3462 4401 3518
rect 4422 3452 4425 3488
rect 4438 3462 4441 3478
rect 4446 3472 4449 3568
rect 4470 3552 4473 3558
rect 4518 3552 4521 3948
rect 4534 3942 4537 3988
rect 4578 3968 4582 3971
rect 4590 3962 4593 3998
rect 4598 3972 4601 4028
rect 4546 3948 4550 3951
rect 4558 3942 4561 3948
rect 4530 3928 4534 3931
rect 4590 3922 4593 3938
rect 4534 3862 4537 3898
rect 4542 3872 4545 3898
rect 4550 3882 4553 3888
rect 4598 3882 4601 3918
rect 4606 3872 4609 4058
rect 4614 4052 4617 4058
rect 4654 4052 4657 4068
rect 4632 4003 4634 4007
rect 4638 4003 4641 4007
rect 4645 4003 4648 4007
rect 4614 3932 4617 3948
rect 4622 3942 4625 3948
rect 4642 3938 4646 3941
rect 4526 3751 4529 3858
rect 4542 3852 4545 3868
rect 4582 3822 4585 3868
rect 4570 3748 4574 3751
rect 4558 3742 4561 3748
rect 4542 3642 4545 3738
rect 4582 3671 4585 3818
rect 4590 3752 4593 3758
rect 4598 3742 4601 3748
rect 4606 3732 4609 3738
rect 4614 3721 4617 3868
rect 4622 3772 4625 3918
rect 4654 3912 4657 3918
rect 4662 3902 4665 4058
rect 4670 3972 4673 4218
rect 4714 4178 4718 4181
rect 4682 4158 4686 4161
rect 4690 4148 4694 4151
rect 4702 4092 4705 4148
rect 4714 4138 4718 4141
rect 4678 3982 4681 4018
rect 4706 3958 4710 3961
rect 4686 3952 4689 3958
rect 4674 3938 4678 3941
rect 4686 3931 4689 3948
rect 4698 3938 4702 3941
rect 4686 3928 4697 3931
rect 4666 3868 4670 3871
rect 4630 3863 4633 3868
rect 4678 3852 4681 3918
rect 4694 3862 4697 3928
rect 4702 3872 4705 3888
rect 4718 3882 4721 4038
rect 4726 3862 4729 4218
rect 4870 4192 4873 4328
rect 4878 4232 4881 4238
rect 4770 4148 4774 4151
rect 4818 4148 4822 4151
rect 4798 4142 4801 4148
rect 4742 4092 4745 4098
rect 4750 4082 4753 4128
rect 4814 4112 4817 4148
rect 4886 4142 4889 4188
rect 4894 4162 4897 4348
rect 4902 4272 4905 4348
rect 4914 4338 4918 4341
rect 4918 4312 4921 4318
rect 4918 4262 4921 4278
rect 4894 4152 4897 4158
rect 4874 4138 4878 4141
rect 4734 4072 4737 4078
rect 4762 4068 4766 4071
rect 4794 4068 4798 4071
rect 4778 4058 4782 4061
rect 4750 3982 4753 3988
rect 4734 3972 4737 3978
rect 4734 3952 4737 3958
rect 4758 3932 4761 3968
rect 4766 3952 4769 4058
rect 4774 4048 4782 4051
rect 4774 3992 4777 4048
rect 4782 3952 4785 3958
rect 4814 3942 4817 4108
rect 4878 4102 4881 4138
rect 4886 4092 4889 4138
rect 4910 4132 4913 4158
rect 4926 4151 4929 4368
rect 4950 4291 4953 4338
rect 4942 4288 4953 4291
rect 4942 4272 4945 4288
rect 4958 4272 4961 4288
rect 4966 4262 4969 4398
rect 4974 4352 4977 4358
rect 4998 4342 5001 4468
rect 5050 4458 5054 4461
rect 5038 4442 5041 4448
rect 5054 4442 5057 4448
rect 5014 4382 5017 4388
rect 5094 4371 5097 4468
rect 5110 4452 5113 4459
rect 5158 4411 5161 4538
rect 5174 4502 5177 4518
rect 5174 4482 5177 4488
rect 5150 4408 5161 4411
rect 5094 4368 5105 4371
rect 5050 4358 5054 4361
rect 5022 4332 5025 4358
rect 5078 4352 5081 4368
rect 5034 4348 5038 4351
rect 5070 4342 5073 4348
rect 5102 4342 5105 4368
rect 5118 4342 5121 4347
rect 5030 4332 5033 4338
rect 5086 4322 5089 4338
rect 5014 4272 5017 4318
rect 5102 4272 5105 4338
rect 5150 4272 5153 4408
rect 5182 4362 5185 4368
rect 5122 4268 5126 4271
rect 5002 4258 5006 4261
rect 4978 4248 4982 4251
rect 5006 4232 5009 4238
rect 4938 4158 4942 4161
rect 5006 4152 5009 4158
rect 4926 4148 4934 4151
rect 4942 4148 4950 4151
rect 4942 4142 4945 4148
rect 4934 4138 4942 4141
rect 4858 4058 4862 4061
rect 4870 3982 4873 4088
rect 4886 4072 4889 4078
rect 4822 3952 4825 3958
rect 4766 3932 4769 3938
rect 4814 3872 4817 3878
rect 4830 3872 4833 3948
rect 4858 3868 4862 3871
rect 4758 3862 4761 3868
rect 4766 3862 4769 3868
rect 4822 3862 4825 3868
rect 4830 3862 4833 3868
rect 4870 3862 4873 3978
rect 4878 3962 4881 3968
rect 4890 3948 4894 3951
rect 4878 3872 4881 3888
rect 4886 3862 4889 3938
rect 4894 3862 4897 3948
rect 4902 3922 4905 4018
rect 4926 3992 4929 4018
rect 4910 3922 4913 3958
rect 4918 3952 4921 3958
rect 4926 3952 4929 3978
rect 4918 3932 4921 3938
rect 4934 3892 4937 4138
rect 4950 4122 4953 4128
rect 4982 4062 4985 4068
rect 4998 4062 5001 4068
rect 4958 4022 4961 4058
rect 4942 3952 4945 3958
rect 4950 3892 4953 3918
rect 4966 3872 4969 3968
rect 4990 3882 4993 3888
rect 4934 3862 4937 3868
rect 4632 3803 4634 3807
rect 4638 3803 4641 3807
rect 4645 3803 4648 3807
rect 4694 3792 4697 3858
rect 4726 3832 4729 3858
rect 4806 3852 4809 3858
rect 4870 3852 4873 3858
rect 4710 3782 4713 3818
rect 4750 3772 4753 3838
rect 4706 3758 4710 3761
rect 4734 3752 4737 3758
rect 4706 3748 4710 3751
rect 4646 3742 4649 3748
rect 4686 3732 4689 3738
rect 4606 3718 4617 3721
rect 4606 3682 4609 3718
rect 4606 3672 4609 3678
rect 4582 3668 4593 3671
rect 4582 3652 4585 3658
rect 4542 3572 4545 3638
rect 4514 3548 4518 3551
rect 4530 3548 4534 3551
rect 4494 3542 4497 3548
rect 4466 3488 4470 3491
rect 4510 3472 4513 3538
rect 4458 3468 4462 3471
rect 4434 3458 4438 3461
rect 4470 3452 4473 3458
rect 4410 3448 4414 3451
rect 4398 3362 4401 3418
rect 4438 3412 4441 3418
rect 4446 3392 4449 3448
rect 4430 3362 4433 3368
rect 4410 3358 4414 3361
rect 4502 3352 4505 3358
rect 4386 3348 4390 3351
rect 4434 3348 4438 3351
rect 4510 3342 4513 3468
rect 4518 3462 4521 3538
rect 4534 3532 4537 3538
rect 4526 3522 4529 3528
rect 4542 3522 4545 3548
rect 4558 3521 4561 3558
rect 4570 3538 4574 3541
rect 4546 3518 4553 3521
rect 4558 3518 4566 3521
rect 4374 3338 4385 3341
rect 4366 3332 4369 3338
rect 4382 3332 4385 3338
rect 4402 3328 4406 3331
rect 4318 3298 4329 3301
rect 4310 3182 4313 3188
rect 4294 3158 4305 3161
rect 4214 3112 4217 3118
rect 4166 3062 4169 3108
rect 4230 3102 4233 3128
rect 4214 3092 4217 3098
rect 4206 3018 4214 3021
rect 4206 2972 4209 3018
rect 4222 2972 4225 3078
rect 4262 3062 4265 3138
rect 4286 3132 4289 3148
rect 4294 3142 4297 3148
rect 4270 3092 4273 3118
rect 4234 3058 4238 3061
rect 4250 3058 4254 3061
rect 4238 3042 4241 3048
rect 4238 2992 4241 3018
rect 4102 2952 4105 2958
rect 4146 2948 4150 2951
rect 4114 2938 4118 2941
rect 4082 2928 4086 2931
rect 4118 2922 4121 2928
rect 3998 2878 4025 2881
rect 3998 2871 4001 2878
rect 4022 2872 4025 2878
rect 4078 2872 4081 2898
rect 3990 2868 4001 2871
rect 3990 2862 3993 2868
rect 4006 2862 4009 2868
rect 4086 2862 4089 2918
rect 4112 2903 4114 2907
rect 4118 2903 4121 2907
rect 4125 2903 4128 2907
rect 4058 2858 4062 2861
rect 4106 2858 4110 2861
rect 4134 2861 4137 2908
rect 4142 2871 4145 2898
rect 4150 2892 4153 2948
rect 4178 2938 4182 2941
rect 4166 2922 4169 2928
rect 4166 2882 4169 2918
rect 4182 2892 4185 2898
rect 4190 2882 4193 2968
rect 4206 2932 4209 2938
rect 4158 2872 4161 2878
rect 4142 2868 4150 2871
rect 4126 2858 4137 2861
rect 4146 2858 4150 2861
rect 3998 2822 4001 2858
rect 3974 2802 3977 2818
rect 3974 2752 3977 2758
rect 3998 2752 4001 2758
rect 4014 2752 4017 2768
rect 3986 2738 3990 2741
rect 3926 2722 3929 2738
rect 3950 2732 3953 2738
rect 3910 2692 3913 2698
rect 3926 2692 3929 2698
rect 3946 2688 3950 2691
rect 3910 2682 3913 2688
rect 3934 2672 3937 2678
rect 3998 2662 4001 2698
rect 4006 2692 4009 2738
rect 4022 2732 4025 2848
rect 4038 2842 4041 2858
rect 4070 2752 4073 2858
rect 4126 2852 4129 2858
rect 4198 2852 4201 2918
rect 4214 2912 4217 2918
rect 4222 2872 4225 2898
rect 4246 2892 4249 2908
rect 4254 2892 4257 2948
rect 4262 2932 4265 3058
rect 4270 3032 4273 3068
rect 4286 3052 4289 3088
rect 4302 3071 4305 3158
rect 4298 3068 4305 3071
rect 4318 3072 4321 3298
rect 4366 3263 4369 3318
rect 4398 3302 4401 3318
rect 4438 3302 4441 3338
rect 4446 3312 4449 3318
rect 4542 3302 4545 3358
rect 4550 3351 4553 3518
rect 4566 3492 4569 3518
rect 4582 3472 4585 3568
rect 4590 3552 4593 3668
rect 4622 3662 4625 3668
rect 4630 3641 4633 3718
rect 4662 3692 4665 3728
rect 4694 3722 4697 3748
rect 4718 3731 4721 3748
rect 4726 3742 4729 3748
rect 4750 3742 4753 3748
rect 4734 3732 4737 3738
rect 4766 3732 4769 3778
rect 4782 3742 4785 3848
rect 4846 3842 4849 3848
rect 4882 3838 4886 3841
rect 4806 3751 4809 3818
rect 4806 3748 4814 3751
rect 4718 3728 4729 3731
rect 4622 3638 4633 3641
rect 4598 3582 4601 3588
rect 4590 3502 4593 3548
rect 4598 3542 4601 3578
rect 4598 3522 4601 3528
rect 4606 3522 4609 3598
rect 4622 3562 4625 3638
rect 4634 3628 4638 3631
rect 4654 3612 4657 3668
rect 4662 3662 4665 3688
rect 4678 3682 4681 3718
rect 4686 3692 4689 3698
rect 4714 3688 4718 3691
rect 4710 3662 4713 3668
rect 4670 3622 4673 3658
rect 4694 3652 4697 3658
rect 4686 3642 4689 3648
rect 4726 3642 4729 3728
rect 4706 3638 4710 3641
rect 4632 3603 4634 3607
rect 4638 3603 4641 3607
rect 4645 3603 4648 3607
rect 4634 3558 4638 3561
rect 4666 3558 4670 3561
rect 4614 3552 4617 3558
rect 4678 3542 4681 3558
rect 4702 3552 4705 3598
rect 4726 3592 4729 3628
rect 4710 3562 4713 3568
rect 4606 3462 4609 3488
rect 4558 3362 4561 3368
rect 4570 3358 4574 3361
rect 4550 3348 4558 3351
rect 4602 3348 4606 3351
rect 4566 3332 4569 3338
rect 4454 3282 4457 3288
rect 4398 3272 4401 3278
rect 4434 3268 4441 3271
rect 4382 3142 4385 3268
rect 4438 3262 4441 3268
rect 4410 3258 4414 3261
rect 4430 3252 4433 3258
rect 4446 3222 4449 3268
rect 4334 3062 4337 3068
rect 4314 3058 4318 3061
rect 4354 3058 4358 3061
rect 4302 3052 4305 3058
rect 4278 3042 4281 3048
rect 4318 3042 4321 3048
rect 4278 2992 4281 3018
rect 4326 3002 4329 3058
rect 4342 3042 4345 3058
rect 4346 2978 4350 2981
rect 4294 2932 4297 2978
rect 4310 2952 4313 2958
rect 4330 2948 4334 2951
rect 4342 2942 4345 2948
rect 4330 2938 4334 2941
rect 4298 2888 4302 2891
rect 4286 2882 4289 2888
rect 4230 2872 4233 2878
rect 4290 2868 4294 2871
rect 4262 2862 4265 2868
rect 4210 2858 4214 2861
rect 4254 2852 4257 2858
rect 4098 2848 4102 2851
rect 4162 2848 4166 2851
rect 4086 2802 4089 2818
rect 4122 2748 4126 2751
rect 4138 2748 4142 2751
rect 4062 2742 4065 2748
rect 4074 2728 4078 2731
rect 4006 2662 4009 2688
rect 4030 2672 4033 2728
rect 3938 2658 3942 2661
rect 3814 2542 3817 2548
rect 3842 2538 3846 2541
rect 3830 2532 3833 2538
rect 3854 2531 3857 2568
rect 3906 2548 3910 2551
rect 3918 2542 3921 2578
rect 3950 2572 3953 2628
rect 3974 2592 3977 2608
rect 4014 2582 4017 2668
rect 4046 2612 4049 2678
rect 4062 2662 4065 2678
rect 3950 2542 3953 2568
rect 4014 2552 4017 2578
rect 3842 2528 3857 2531
rect 3798 2482 3801 2488
rect 3758 2462 3761 2468
rect 3782 2462 3785 2468
rect 3766 2452 3769 2458
rect 3782 2412 3785 2458
rect 3798 2392 3801 2478
rect 3918 2472 3921 2508
rect 3858 2468 3862 2471
rect 3914 2468 3918 2471
rect 3846 2462 3849 2468
rect 3814 2452 3817 2458
rect 3822 2442 3825 2458
rect 3886 2422 3889 2458
rect 3758 2342 3761 2388
rect 3782 2362 3785 2368
rect 3790 2352 3793 2388
rect 3846 2362 3849 2398
rect 3878 2382 3881 2418
rect 3894 2372 3897 2468
rect 3902 2452 3905 2468
rect 3934 2462 3937 2468
rect 3910 2452 3913 2458
rect 3930 2448 3934 2451
rect 3938 2438 3942 2441
rect 3950 2441 3953 2538
rect 4022 2532 4025 2578
rect 4038 2551 4041 2598
rect 3958 2502 3961 2518
rect 4054 2512 4057 2648
rect 4062 2618 4070 2621
rect 4062 2602 4065 2618
rect 3958 2478 3974 2481
rect 3958 2472 3961 2478
rect 3978 2468 3982 2471
rect 3958 2452 3961 2458
rect 3950 2438 3961 2441
rect 3870 2362 3873 2368
rect 3814 2342 3817 2358
rect 3846 2352 3849 2358
rect 3834 2348 3841 2351
rect 3866 2348 3870 2351
rect 3910 2351 3913 2358
rect 3826 2338 3830 2341
rect 3766 2332 3769 2338
rect 3838 2332 3841 2348
rect 3742 2262 3745 2318
rect 3798 2292 3801 2318
rect 3878 2302 3881 2338
rect 3782 2272 3785 2288
rect 3750 2268 3777 2271
rect 3806 2271 3809 2288
rect 3798 2268 3809 2271
rect 3814 2272 3817 2298
rect 3902 2292 3905 2298
rect 3826 2288 3830 2291
rect 3750 2262 3753 2268
rect 3774 2261 3777 2268
rect 3774 2258 3782 2261
rect 3798 2261 3801 2268
rect 3838 2262 3841 2268
rect 3790 2258 3801 2261
rect 3726 2242 3729 2258
rect 3758 2252 3761 2258
rect 3790 2252 3793 2258
rect 3806 2252 3809 2258
rect 3846 2252 3849 2278
rect 3862 2262 3865 2288
rect 3886 2272 3889 2288
rect 3910 2282 3913 2308
rect 3766 2242 3769 2248
rect 3822 2242 3825 2248
rect 3862 2242 3865 2258
rect 3894 2242 3897 2258
rect 3918 2242 3921 2248
rect 3870 2232 3873 2238
rect 3742 2182 3745 2188
rect 3722 2178 3726 2181
rect 3710 2168 3721 2171
rect 3710 2091 3713 2128
rect 3706 2088 3713 2091
rect 3670 2062 3673 2068
rect 3608 2003 3610 2007
rect 3614 2003 3617 2007
rect 3621 2003 3624 2007
rect 3550 1948 3558 1951
rect 3550 1932 3553 1948
rect 3574 1942 3577 1948
rect 3582 1942 3585 1998
rect 3646 1992 3649 2048
rect 3654 2012 3657 2058
rect 3686 1992 3689 2078
rect 3718 2072 3721 2168
rect 3726 2092 3729 2158
rect 3734 2142 3737 2178
rect 3766 2162 3769 2218
rect 3774 2202 3777 2218
rect 3786 2158 3790 2161
rect 3766 2152 3769 2158
rect 3790 2152 3793 2158
rect 3746 2148 3750 2151
rect 3806 2142 3809 2168
rect 3754 2138 3758 2141
rect 3774 2132 3777 2138
rect 3814 2112 3817 2158
rect 3830 2141 3833 2158
rect 3838 2152 3841 2188
rect 3862 2152 3865 2158
rect 3830 2138 3838 2141
rect 3850 2138 3862 2141
rect 3822 2122 3825 2138
rect 3722 2068 3726 2071
rect 3710 1982 3713 2068
rect 3782 2062 3785 2078
rect 3846 2062 3849 2068
rect 3726 2052 3729 2058
rect 3790 1982 3793 2058
rect 3814 2018 3822 2021
rect 3798 1992 3801 2018
rect 3590 1952 3593 1978
rect 3750 1968 3766 1971
rect 3750 1961 3753 1968
rect 3742 1958 3753 1961
rect 3786 1958 3790 1961
rect 3590 1942 3593 1948
rect 3558 1932 3561 1938
rect 3542 1902 3545 1918
rect 3574 1892 3577 1908
rect 3606 1892 3609 1958
rect 3622 1952 3625 1958
rect 3718 1952 3721 1958
rect 3742 1952 3745 1958
rect 3766 1952 3769 1958
rect 3806 1952 3809 2018
rect 3814 1972 3817 2018
rect 3846 1992 3849 2058
rect 3826 1958 3830 1961
rect 3854 1961 3857 2128
rect 3866 2078 3870 2081
rect 3866 2068 3870 2071
rect 3878 2062 3881 2228
rect 3890 2168 3921 2171
rect 3918 2162 3921 2168
rect 3906 2158 3910 2161
rect 3890 2148 3894 2151
rect 3886 2092 3889 2108
rect 3910 2082 3913 2098
rect 3902 2072 3905 2078
rect 3910 2062 3913 2078
rect 3926 2072 3929 2278
rect 3934 2242 3937 2348
rect 3958 2122 3961 2438
rect 3966 2412 3969 2468
rect 3990 2462 3993 2468
rect 3998 2442 4001 2458
rect 3982 2352 3985 2418
rect 3998 2352 4001 2358
rect 4006 2342 4009 2508
rect 4054 2472 4057 2508
rect 4034 2468 4038 2471
rect 4014 2462 4017 2468
rect 4070 2462 4073 2608
rect 4078 2592 4081 2708
rect 4112 2703 4114 2707
rect 4118 2703 4121 2707
rect 4125 2703 4128 2707
rect 4086 2672 4089 2678
rect 4134 2662 4137 2698
rect 4142 2672 4145 2718
rect 4094 2622 4097 2658
rect 4142 2652 4145 2658
rect 4158 2642 4161 2708
rect 4166 2662 4169 2798
rect 4174 2762 4177 2848
rect 4214 2832 4217 2838
rect 4182 2752 4185 2808
rect 4198 2692 4201 2818
rect 4246 2802 4249 2848
rect 4206 2752 4209 2798
rect 4230 2792 4233 2798
rect 4234 2748 4241 2751
rect 4186 2658 4190 2661
rect 4178 2648 4185 2651
rect 4094 2552 4097 2588
rect 4110 2572 4113 2618
rect 4158 2562 4161 2618
rect 4158 2552 4161 2558
rect 4166 2552 4169 2558
rect 4130 2548 4134 2551
rect 4106 2538 4110 2541
rect 4082 2528 4086 2531
rect 4112 2503 4114 2507
rect 4118 2503 4121 2507
rect 4125 2503 4128 2507
rect 4078 2492 4081 2498
rect 4102 2472 4105 2488
rect 4090 2468 4094 2471
rect 4110 2462 4113 2468
rect 4030 2422 4033 2458
rect 4038 2442 4041 2448
rect 4014 2352 4017 2378
rect 4022 2352 4025 2358
rect 3986 2338 3990 2341
rect 4022 2332 4025 2338
rect 3974 2312 3977 2318
rect 3998 2272 4001 2298
rect 3974 2252 3977 2258
rect 3974 2152 3977 2158
rect 3998 2142 4001 2268
rect 4030 2262 4033 2358
rect 4046 2352 4049 2458
rect 4086 2452 4089 2458
rect 4066 2448 4070 2451
rect 4054 2352 4057 2358
rect 4038 2342 4041 2348
rect 4070 2342 4073 2408
rect 4094 2392 4097 2448
rect 4118 2412 4121 2468
rect 4126 2352 4129 2458
rect 4134 2352 4137 2498
rect 4142 2472 4145 2538
rect 4150 2471 4153 2548
rect 4174 2512 4177 2538
rect 4162 2478 4166 2481
rect 4150 2468 4161 2471
rect 4150 2442 4153 2458
rect 4158 2452 4161 2468
rect 4046 2332 4049 2338
rect 4054 2292 4057 2338
rect 4078 2302 4081 2328
rect 4078 2272 4081 2298
rect 4046 2252 4049 2258
rect 4070 2252 4073 2258
rect 4022 2192 4025 2218
rect 4054 2172 4057 2218
rect 4062 2172 4065 2238
rect 4086 2192 4089 2348
rect 4112 2303 4114 2307
rect 4118 2303 4121 2307
rect 4125 2303 4128 2307
rect 4078 2152 4081 2188
rect 4110 2152 4113 2158
rect 4026 2148 4030 2151
rect 4038 2142 4041 2148
rect 3966 2092 3969 2098
rect 3946 2068 3950 2071
rect 3926 2062 3929 2068
rect 3998 2062 4001 2138
rect 4014 2132 4017 2138
rect 4046 2132 4049 2138
rect 3938 2058 3942 2061
rect 3878 1992 3881 2058
rect 3846 1958 3857 1961
rect 3658 1948 3662 1951
rect 3754 1948 3758 1951
rect 3630 1912 3633 1948
rect 3670 1942 3673 1948
rect 3758 1932 3761 1938
rect 3794 1928 3798 1931
rect 3534 1882 3537 1888
rect 3546 1878 3550 1881
rect 3578 1868 3582 1871
rect 3550 1792 3553 1868
rect 3558 1862 3561 1868
rect 3590 1862 3593 1868
rect 3558 1802 3561 1858
rect 3598 1852 3601 1878
rect 3638 1872 3641 1878
rect 3582 1792 3585 1828
rect 3418 1778 3422 1781
rect 3450 1758 3473 1761
rect 3398 1692 3401 1728
rect 3422 1722 3425 1748
rect 3430 1732 3433 1758
rect 3470 1752 3473 1758
rect 3518 1758 3526 1761
rect 3562 1758 3566 1761
rect 3458 1748 3462 1751
rect 3498 1748 3502 1751
rect 3310 1678 3321 1681
rect 3414 1682 3417 1688
rect 3310 1672 3313 1678
rect 3322 1668 3326 1671
rect 3386 1668 3390 1671
rect 3302 1652 3305 1658
rect 3382 1648 3390 1651
rect 3286 1611 3289 1648
rect 3306 1638 3310 1641
rect 3278 1608 3289 1611
rect 3254 1552 3257 1558
rect 3158 1492 3161 1538
rect 3190 1492 3193 1508
rect 3246 1492 3249 1538
rect 3278 1522 3281 1608
rect 3382 1602 3385 1648
rect 3310 1592 3313 1598
rect 3330 1578 3334 1581
rect 3318 1552 3321 1558
rect 3342 1552 3345 1578
rect 3382 1572 3385 1598
rect 3406 1592 3409 1668
rect 3446 1662 3449 1748
rect 3510 1742 3513 1748
rect 3458 1738 3465 1741
rect 3454 1692 3457 1728
rect 3462 1692 3465 1738
rect 3518 1712 3521 1758
rect 3526 1712 3529 1718
rect 3482 1688 3486 1691
rect 3438 1652 3441 1658
rect 3446 1648 3454 1651
rect 3414 1592 3417 1608
rect 3362 1558 3366 1561
rect 3342 1532 3345 1538
rect 3350 1532 3353 1538
rect 3094 1472 3097 1488
rect 3102 1482 3105 1488
rect 3158 1482 3161 1488
rect 3110 1472 3113 1478
rect 3182 1472 3185 1478
rect 3130 1468 3134 1471
rect 3154 1468 3158 1471
rect 3094 1402 3097 1448
rect 3110 1412 3113 1468
rect 3122 1418 3126 1421
rect 3094 1362 3097 1398
rect 3118 1348 3126 1351
rect 3110 1322 3113 1328
rect 3096 1303 3098 1307
rect 3102 1303 3105 1307
rect 3109 1303 3112 1307
rect 3098 1268 3102 1271
rect 3102 1142 3105 1198
rect 3096 1103 3098 1107
rect 3102 1103 3105 1107
rect 3109 1103 3112 1107
rect 3110 1032 3113 1068
rect 3118 1062 3121 1348
rect 3134 1342 3137 1468
rect 3198 1462 3201 1488
rect 3222 1482 3225 1488
rect 3206 1462 3209 1468
rect 3230 1462 3233 1468
rect 3154 1458 3158 1461
rect 3166 1458 3174 1461
rect 3150 1422 3153 1448
rect 3166 1332 3169 1458
rect 3254 1442 3257 1458
rect 3182 1332 3185 1408
rect 3198 1392 3201 1428
rect 3190 1372 3193 1388
rect 3214 1372 3217 1418
rect 3190 1362 3193 1368
rect 3262 1342 3265 1408
rect 3202 1338 3206 1341
rect 3218 1338 3222 1341
rect 3138 1328 3142 1331
rect 3186 1328 3190 1331
rect 3150 1292 3153 1298
rect 3126 1272 3129 1288
rect 3154 1268 3158 1271
rect 3166 1262 3169 1328
rect 3222 1322 3225 1328
rect 3250 1318 3254 1321
rect 3154 1248 3158 1251
rect 3158 1238 3166 1241
rect 3158 1192 3161 1238
rect 3150 1152 3153 1188
rect 3174 1162 3177 1318
rect 3190 1272 3193 1318
rect 3182 1252 3185 1258
rect 3190 1241 3193 1258
rect 3186 1238 3193 1241
rect 3198 1192 3201 1308
rect 3214 1282 3217 1298
rect 3226 1288 3230 1291
rect 3238 1252 3241 1308
rect 3246 1292 3249 1298
rect 3262 1282 3265 1338
rect 3270 1282 3273 1488
rect 3282 1358 3286 1361
rect 3290 1318 3294 1321
rect 3258 1268 3262 1271
rect 3226 1248 3230 1251
rect 3206 1242 3209 1248
rect 3154 1138 3161 1141
rect 3126 1112 3129 1118
rect 3146 1058 3150 1061
rect 3158 1051 3161 1138
rect 3150 1048 3161 1051
rect 3094 1002 3097 1018
rect 3094 932 3097 938
rect 3110 932 3113 1028
rect 3150 992 3153 1048
rect 3166 982 3169 1128
rect 3174 1122 3177 1148
rect 3206 1132 3209 1148
rect 3214 1142 3217 1148
rect 3222 1122 3225 1148
rect 3230 1132 3233 1138
rect 3186 1068 3190 1071
rect 3194 1038 3198 1041
rect 3096 903 3098 907
rect 3102 903 3105 907
rect 3109 903 3112 907
rect 3118 902 3121 948
rect 3098 888 3102 891
rect 3118 842 3121 868
rect 3126 862 3129 968
rect 3174 962 3177 1018
rect 3202 948 3206 951
rect 3174 942 3177 948
rect 3158 932 3161 938
rect 3134 922 3137 928
rect 3150 852 3153 888
rect 3174 872 3177 878
rect 3130 848 3134 851
rect 3154 848 3158 851
rect 3038 762 3041 768
rect 3018 758 3022 761
rect 3010 748 3014 751
rect 3006 732 3009 738
rect 3046 672 3049 758
rect 3054 752 3057 778
rect 3102 752 3105 758
rect 3110 752 3113 818
rect 3118 752 3121 838
rect 3166 822 3169 858
rect 2918 542 2921 548
rect 2866 488 2870 491
rect 2862 472 2865 478
rect 2786 468 2793 471
rect 2826 468 2830 471
rect 2774 442 2777 448
rect 2774 382 2777 408
rect 2774 352 2777 378
rect 2782 352 2785 468
rect 2798 462 2801 468
rect 2834 458 2838 461
rect 2850 458 2854 461
rect 2790 402 2793 458
rect 2806 452 2809 458
rect 2814 452 2817 458
rect 2834 448 2838 451
rect 2842 388 2846 391
rect 2806 362 2809 368
rect 2794 358 2798 361
rect 2814 352 2817 388
rect 2810 348 2814 351
rect 2770 338 2774 341
rect 2718 272 2721 338
rect 2602 258 2606 261
rect 2698 258 2702 261
rect 2510 252 2513 258
rect 2358 188 2369 191
rect 2278 152 2281 158
rect 2294 152 2297 178
rect 2326 172 2329 178
rect 2310 162 2313 168
rect 2342 162 2345 168
rect 2326 152 2329 158
rect 2314 148 2318 151
rect 2286 142 2289 148
rect 2358 142 2361 188
rect 2434 168 2438 171
rect 2374 142 2377 147
rect 2274 138 2278 141
rect 2278 132 2281 138
rect 2318 132 2321 138
rect 2254 122 2257 128
rect 2334 92 2337 118
rect 2430 92 2433 128
rect 2446 92 2449 118
rect 2478 82 2481 148
rect 2238 72 2241 78
rect 2350 72 2353 78
rect 2494 72 2497 228
rect 2510 151 2513 158
rect 2526 92 2529 218
rect 2584 203 2586 207
rect 2590 203 2593 207
rect 2597 203 2600 207
rect 2614 152 2617 258
rect 2678 242 2681 248
rect 2686 202 2689 258
rect 2694 242 2697 248
rect 2726 192 2729 268
rect 2734 262 2737 298
rect 2702 182 2705 188
rect 2718 181 2721 188
rect 2710 178 2721 181
rect 2642 168 2646 171
rect 2654 162 2657 178
rect 2686 162 2689 168
rect 2678 152 2681 158
rect 2710 152 2713 178
rect 2602 148 2606 151
rect 2658 148 2662 151
rect 2706 138 2710 141
rect 2678 132 2681 138
rect 2718 132 2721 168
rect 2726 121 2729 178
rect 2734 142 2737 168
rect 2742 152 2745 258
rect 2750 202 2753 328
rect 2798 322 2801 338
rect 2830 332 2833 358
rect 2854 352 2857 458
rect 2862 422 2865 468
rect 2878 382 2881 498
rect 2902 492 2905 528
rect 2918 472 2921 498
rect 2874 348 2878 351
rect 2758 272 2761 308
rect 2790 282 2793 318
rect 2830 292 2833 328
rect 2774 272 2777 278
rect 2758 172 2761 238
rect 2790 232 2793 268
rect 2806 263 2809 278
rect 2854 242 2857 338
rect 2866 288 2870 291
rect 2878 262 2881 308
rect 2854 232 2857 238
rect 2766 162 2769 198
rect 2782 152 2785 188
rect 2818 168 2822 171
rect 2846 168 2854 171
rect 2798 162 2801 168
rect 2830 162 2833 168
rect 2846 152 2849 168
rect 2866 158 2870 161
rect 2810 148 2814 151
rect 2734 132 2737 138
rect 2718 118 2729 121
rect 2538 88 2542 91
rect 2614 72 2617 98
rect 2678 72 2681 78
rect 2102 62 2105 68
rect 2166 62 2169 68
rect 2254 62 2257 68
rect 2446 62 2449 68
rect 2282 58 2286 61
rect 2378 58 2382 61
rect 2474 58 2478 61
rect 2630 62 2633 68
rect 2670 62 2673 68
rect 2686 62 2689 118
rect 2718 92 2721 118
rect 938 48 942 51
rect 962 48 966 51
rect 950 42 953 48
rect 2598 42 2601 59
rect 2702 52 2705 68
rect 2742 62 2745 148
rect 2822 142 2825 148
rect 2786 138 2790 141
rect 2750 82 2753 138
rect 2846 122 2849 148
rect 2858 138 2862 141
rect 2790 82 2793 88
rect 2734 52 2737 58
rect 2650 48 2654 51
rect 2686 42 2689 48
rect 2750 32 2753 68
rect 2766 62 2769 68
rect 2822 63 2825 68
rect 2830 62 2833 118
rect 2862 112 2865 118
rect 2838 72 2841 98
rect 2842 68 2846 71
rect 2774 32 2777 58
rect 2878 52 2881 258
rect 2886 152 2889 418
rect 2918 372 2921 468
rect 2902 272 2905 318
rect 2894 258 2902 261
rect 2894 222 2897 258
rect 2894 192 2897 218
rect 2926 201 2929 568
rect 2966 552 2969 578
rect 2974 552 2977 658
rect 2990 572 2993 638
rect 3006 632 3009 668
rect 3014 662 3017 668
rect 3054 662 3057 748
rect 3070 742 3073 748
rect 3078 722 3081 748
rect 3118 732 3121 748
rect 3096 703 3098 707
rect 3102 703 3105 707
rect 3109 703 3112 707
rect 3062 672 3065 688
rect 3114 668 3118 671
rect 3078 662 3081 668
rect 3126 662 3129 818
rect 3174 782 3177 868
rect 3182 842 3185 868
rect 3190 862 3193 868
rect 3134 762 3137 768
rect 3154 758 3158 761
rect 3178 758 3182 761
rect 3198 751 3201 938
rect 3206 892 3209 898
rect 3214 852 3217 928
rect 3190 748 3201 751
rect 3210 748 3214 751
rect 3150 732 3153 738
rect 3174 732 3177 738
rect 3182 722 3185 738
rect 3122 658 3126 661
rect 3022 652 3025 658
rect 2998 592 3001 608
rect 3046 592 3049 638
rect 3010 588 3014 591
rect 2994 558 3001 561
rect 2954 548 2958 551
rect 2946 538 2950 541
rect 2958 532 2961 538
rect 2934 463 2937 518
rect 2934 392 2937 438
rect 2950 392 2953 518
rect 2966 472 2969 478
rect 2978 458 2982 461
rect 2974 412 2977 418
rect 2958 362 2961 408
rect 2982 362 2985 458
rect 2990 452 2993 528
rect 2998 492 3001 558
rect 2990 442 2993 448
rect 2974 352 2977 358
rect 2962 348 2966 351
rect 2982 342 2985 348
rect 2990 342 2993 418
rect 2998 372 3001 438
rect 3014 432 3017 468
rect 3022 462 3025 578
rect 3038 502 3041 548
rect 3038 482 3041 498
rect 3038 462 3041 468
rect 3054 462 3057 638
rect 3094 582 3097 658
rect 3142 652 3145 688
rect 3166 682 3169 718
rect 3182 691 3185 718
rect 3174 688 3185 691
rect 3174 672 3177 688
rect 3190 682 3193 748
rect 3222 741 3225 1068
rect 3238 1062 3241 1098
rect 3246 902 3249 1268
rect 3278 1261 3281 1318
rect 3310 1292 3313 1528
rect 3350 1472 3353 1488
rect 3318 1463 3321 1468
rect 3334 1432 3337 1468
rect 3358 1452 3361 1548
rect 3366 1492 3369 1548
rect 3398 1492 3401 1548
rect 3406 1542 3409 1578
rect 3430 1562 3433 1568
rect 3418 1528 3422 1531
rect 3446 1492 3449 1648
rect 3470 1562 3473 1678
rect 3510 1662 3513 1668
rect 3494 1551 3497 1578
rect 3510 1542 3513 1658
rect 3526 1552 3529 1558
rect 3534 1552 3537 1748
rect 3574 1672 3577 1778
rect 3590 1752 3593 1828
rect 3614 1822 3617 1868
rect 3638 1842 3641 1858
rect 3608 1803 3610 1807
rect 3614 1803 3617 1807
rect 3621 1803 3624 1807
rect 3646 1792 3649 1918
rect 3678 1882 3681 1928
rect 3806 1882 3809 1948
rect 3838 1942 3841 1958
rect 3830 1932 3833 1938
rect 3838 1911 3841 1918
rect 3830 1908 3841 1911
rect 3674 1878 3678 1881
rect 3814 1862 3817 1878
rect 3658 1858 3662 1861
rect 3738 1858 3742 1861
rect 3666 1848 3670 1851
rect 3718 1842 3721 1858
rect 3658 1778 3662 1781
rect 3606 1732 3609 1778
rect 3630 1742 3633 1758
rect 3646 1752 3649 1758
rect 3654 1748 3662 1751
rect 3706 1748 3710 1751
rect 3646 1692 3649 1718
rect 3542 1652 3545 1659
rect 3574 1631 3577 1658
rect 3606 1652 3609 1688
rect 3646 1672 3649 1678
rect 3654 1662 3657 1748
rect 3686 1732 3689 1748
rect 3718 1742 3721 1838
rect 3790 1802 3793 1818
rect 3750 1742 3753 1788
rect 3806 1782 3809 1858
rect 3830 1852 3833 1908
rect 3782 1772 3785 1778
rect 3830 1772 3833 1818
rect 3838 1752 3841 1898
rect 3846 1872 3849 1958
rect 3866 1948 3870 1951
rect 3854 1942 3857 1948
rect 3862 1892 3865 1928
rect 3870 1892 3873 1898
rect 3858 1848 3862 1851
rect 3870 1792 3873 1878
rect 3878 1872 3881 1918
rect 3886 1902 3889 2048
rect 3906 1958 3910 1961
rect 3894 1932 3897 1958
rect 3918 1952 3921 1968
rect 3950 1951 3953 1958
rect 3910 1941 3913 1948
rect 3910 1938 3918 1941
rect 3958 1932 3961 2058
rect 3982 1982 3985 2038
rect 3982 1952 3985 1978
rect 3998 1962 4001 2028
rect 3770 1748 3774 1751
rect 3646 1658 3654 1661
rect 3638 1652 3641 1658
rect 3582 1642 3585 1648
rect 3574 1628 3585 1631
rect 3582 1582 3585 1628
rect 3608 1603 3610 1607
rect 3614 1603 3617 1607
rect 3621 1603 3624 1607
rect 3570 1578 3574 1581
rect 3546 1558 3558 1561
rect 3582 1552 3585 1578
rect 3614 1552 3617 1558
rect 3542 1542 3545 1548
rect 3590 1542 3593 1548
rect 3390 1462 3393 1488
rect 3442 1468 3446 1471
rect 3458 1468 3462 1471
rect 3398 1462 3401 1468
rect 3406 1462 3409 1468
rect 3374 1452 3377 1458
rect 3422 1452 3425 1458
rect 3394 1448 3406 1451
rect 3318 1342 3321 1348
rect 3278 1258 3286 1261
rect 3294 1252 3297 1258
rect 3302 1242 3305 1268
rect 3286 1202 3289 1218
rect 3290 1188 3294 1191
rect 3266 1148 3270 1151
rect 3254 1141 3257 1148
rect 3254 1138 3265 1141
rect 3254 1092 3257 1118
rect 3262 1102 3265 1138
rect 3262 1072 3265 1078
rect 3254 962 3257 968
rect 3262 952 3265 1058
rect 3278 1052 3281 1148
rect 3274 948 3278 951
rect 3266 938 3270 941
rect 3286 932 3289 1178
rect 3310 1152 3313 1168
rect 3302 1142 3305 1148
rect 3310 1142 3313 1148
rect 3298 1078 3302 1081
rect 3298 958 3302 961
rect 3318 952 3321 1278
rect 3334 1272 3337 1378
rect 3350 1311 3353 1347
rect 3342 1308 3353 1311
rect 3342 1292 3345 1308
rect 3358 1262 3361 1268
rect 3326 1212 3329 1258
rect 3358 1232 3361 1258
rect 3366 1222 3369 1438
rect 3374 1282 3377 1358
rect 3382 1352 3385 1428
rect 3430 1372 3433 1468
rect 3470 1452 3473 1458
rect 3454 1402 3457 1448
rect 3478 1432 3481 1528
rect 3534 1492 3537 1518
rect 3542 1492 3545 1538
rect 3510 1462 3513 1488
rect 3542 1482 3545 1488
rect 3522 1468 3526 1471
rect 3518 1462 3521 1468
rect 3550 1462 3553 1538
rect 3566 1462 3569 1538
rect 3582 1492 3585 1538
rect 3574 1462 3577 1468
rect 3606 1462 3609 1468
rect 3622 1462 3625 1578
rect 3630 1462 3633 1638
rect 3646 1552 3649 1658
rect 3662 1542 3665 1728
rect 3686 1692 3689 1698
rect 3726 1682 3729 1688
rect 3702 1662 3705 1668
rect 3750 1662 3753 1728
rect 3758 1722 3761 1748
rect 3798 1732 3801 1748
rect 3806 1742 3809 1748
rect 3758 1672 3761 1678
rect 3762 1668 3766 1671
rect 3706 1658 3713 1661
rect 3690 1648 3697 1651
rect 3670 1642 3673 1648
rect 3674 1638 3681 1641
rect 3650 1488 3654 1491
rect 3662 1472 3665 1528
rect 3670 1512 3673 1548
rect 3670 1492 3673 1498
rect 3414 1362 3417 1368
rect 3438 1352 3441 1358
rect 3470 1351 3473 1418
rect 3494 1402 3497 1438
rect 3382 1342 3385 1348
rect 3502 1342 3505 1348
rect 3382 1262 3385 1288
rect 3326 1182 3329 1208
rect 3350 1152 3353 1218
rect 3374 1192 3377 1238
rect 3338 1148 3342 1151
rect 3378 1148 3382 1151
rect 3326 1122 3329 1128
rect 3358 1112 3361 1148
rect 3366 1072 3369 1088
rect 3382 1072 3385 1078
rect 3350 1063 3353 1068
rect 3314 948 3318 951
rect 3310 938 3318 941
rect 3238 872 3241 878
rect 3246 862 3249 878
rect 3254 872 3257 928
rect 3230 822 3233 858
rect 3254 782 3257 868
rect 3266 858 3270 861
rect 3278 851 3281 918
rect 3310 892 3313 938
rect 3326 932 3329 958
rect 3350 952 3353 968
rect 3362 958 3366 961
rect 3318 892 3321 898
rect 3290 868 3305 871
rect 3302 862 3305 868
rect 3290 858 3294 861
rect 3278 848 3286 851
rect 3262 792 3265 828
rect 3266 748 3270 751
rect 3214 738 3225 741
rect 3198 732 3201 738
rect 3190 672 3193 678
rect 3154 668 3158 671
rect 3166 662 3169 668
rect 3206 663 3209 668
rect 3158 658 3166 661
rect 3070 542 3073 547
rect 3086 472 3089 558
rect 3118 532 3121 588
rect 3138 548 3142 551
rect 3138 538 3142 541
rect 3096 503 3098 507
rect 3102 503 3105 507
rect 3109 503 3112 507
rect 3138 468 3142 471
rect 3014 362 3017 388
rect 2998 352 3001 358
rect 2934 251 2937 268
rect 2942 262 2945 328
rect 2974 282 2977 338
rect 2998 292 3001 348
rect 2974 272 2977 278
rect 3006 272 3009 318
rect 3022 312 3025 458
rect 3054 452 3057 458
rect 3102 442 3105 468
rect 3110 462 3113 468
rect 3150 462 3153 528
rect 3158 472 3161 658
rect 3166 552 3169 618
rect 3174 552 3177 628
rect 3182 592 3185 638
rect 3214 612 3217 738
rect 3222 612 3225 718
rect 3238 692 3241 728
rect 3278 692 3281 758
rect 3286 742 3289 798
rect 3294 792 3297 818
rect 3310 802 3313 888
rect 3374 872 3377 1038
rect 3390 1012 3393 1298
rect 3414 1292 3417 1328
rect 3422 1302 3425 1338
rect 3438 1332 3441 1338
rect 3518 1302 3521 1458
rect 3526 1362 3529 1458
rect 3570 1448 3582 1451
rect 3550 1432 3553 1438
rect 3534 1392 3537 1398
rect 3550 1391 3553 1428
rect 3546 1388 3553 1391
rect 3598 1352 3601 1418
rect 3608 1403 3610 1407
rect 3614 1403 3617 1407
rect 3621 1403 3624 1407
rect 3646 1392 3649 1448
rect 3406 1262 3409 1268
rect 3430 1262 3433 1288
rect 3446 1272 3449 1288
rect 3470 1272 3473 1278
rect 3414 1252 3417 1258
rect 3398 1192 3401 1218
rect 3438 1202 3441 1268
rect 3446 1252 3449 1258
rect 3474 1248 3478 1251
rect 3462 1182 3465 1238
rect 3494 1202 3497 1218
rect 3502 1162 3505 1168
rect 3526 1162 3529 1218
rect 3462 1151 3465 1158
rect 3506 1148 3510 1151
rect 3398 1062 3401 1108
rect 3422 1072 3425 1108
rect 3462 1092 3465 1098
rect 3478 1092 3481 1138
rect 3494 1132 3497 1138
rect 3410 1068 3414 1071
rect 3442 1068 3449 1071
rect 3430 1062 3433 1068
rect 3438 1052 3441 1058
rect 3446 1041 3449 1068
rect 3438 1038 3449 1041
rect 3398 992 3401 1038
rect 3346 868 3350 871
rect 3382 862 3385 868
rect 3326 832 3329 858
rect 3294 752 3297 788
rect 3306 758 3310 761
rect 3310 692 3313 758
rect 3330 748 3334 751
rect 3342 742 3345 838
rect 3358 772 3361 838
rect 3374 782 3377 858
rect 3338 738 3342 741
rect 3350 732 3353 758
rect 3374 742 3377 778
rect 3390 742 3393 748
rect 3362 738 3366 741
rect 3318 701 3321 718
rect 3318 698 3329 701
rect 3266 688 3270 691
rect 3310 672 3313 678
rect 3290 668 3294 671
rect 3326 663 3329 698
rect 3214 562 3217 568
rect 3198 552 3201 558
rect 3258 548 3262 551
rect 3174 542 3177 548
rect 3186 538 3190 541
rect 3174 512 3177 528
rect 3174 472 3177 478
rect 3214 472 3217 518
rect 3254 492 3257 498
rect 3190 463 3193 468
rect 3254 462 3257 488
rect 3270 482 3273 548
rect 3278 502 3281 638
rect 3310 592 3313 598
rect 3342 562 3345 588
rect 3318 558 3326 561
rect 3318 552 3321 558
rect 3330 548 3334 551
rect 3322 538 3326 541
rect 3334 532 3337 548
rect 3350 541 3353 558
rect 3358 552 3361 718
rect 3398 692 3401 958
rect 3414 952 3417 958
rect 3422 952 3425 978
rect 3426 948 3433 951
rect 3406 942 3409 948
rect 3410 878 3414 881
rect 3406 842 3409 868
rect 3418 858 3422 861
rect 3422 832 3425 838
rect 3406 762 3409 768
rect 3422 752 3425 788
rect 3430 781 3433 948
rect 3438 841 3441 1038
rect 3454 942 3457 1078
rect 3502 1072 3505 1088
rect 3482 1068 3486 1071
rect 3526 1062 3529 1088
rect 3534 1072 3537 1258
rect 3542 1152 3545 1158
rect 3550 1142 3553 1298
rect 3574 1272 3577 1348
rect 3614 1272 3617 1298
rect 3638 1262 3641 1388
rect 3654 1362 3657 1368
rect 3662 1362 3665 1468
rect 3678 1462 3681 1638
rect 3694 1492 3697 1648
rect 3710 1522 3713 1658
rect 3726 1592 3729 1638
rect 3734 1562 3737 1658
rect 3774 1652 3777 1658
rect 3790 1652 3793 1708
rect 3798 1662 3801 1678
rect 3806 1672 3809 1738
rect 3814 1722 3817 1748
rect 3838 1742 3841 1748
rect 3830 1722 3833 1728
rect 3822 1718 3830 1721
rect 3814 1672 3817 1678
rect 3806 1652 3809 1658
rect 3750 1552 3753 1578
rect 3782 1552 3785 1628
rect 3814 1622 3817 1668
rect 3822 1662 3825 1718
rect 3878 1691 3881 1868
rect 3934 1863 3937 1908
rect 3998 1872 4001 1878
rect 3978 1868 3982 1871
rect 3902 1842 3905 1858
rect 3906 1838 3913 1841
rect 3870 1688 3881 1691
rect 3910 1742 3913 1838
rect 3910 1732 3913 1738
rect 3870 1672 3873 1688
rect 3910 1672 3913 1728
rect 3918 1712 3921 1748
rect 3854 1662 3857 1668
rect 3906 1659 3910 1662
rect 3842 1638 3846 1641
rect 3790 1612 3793 1618
rect 3794 1558 3798 1561
rect 3758 1532 3761 1538
rect 3726 1522 3729 1528
rect 3766 1522 3769 1528
rect 3734 1512 3737 1518
rect 3782 1492 3785 1548
rect 3806 1522 3809 1558
rect 3822 1552 3825 1608
rect 3838 1592 3841 1628
rect 3862 1612 3865 1658
rect 3910 1592 3913 1608
rect 3874 1578 3878 1581
rect 3854 1552 3857 1558
rect 3846 1541 3849 1548
rect 3862 1542 3865 1548
rect 3918 1542 3921 1548
rect 3926 1542 3929 1688
rect 3846 1538 3857 1541
rect 3854 1522 3857 1538
rect 3846 1492 3849 1518
rect 3686 1472 3689 1488
rect 3714 1468 3718 1471
rect 3866 1468 3870 1471
rect 3714 1458 3718 1461
rect 3734 1452 3737 1458
rect 3682 1448 3686 1451
rect 3674 1358 3689 1361
rect 3686 1352 3689 1358
rect 3674 1348 3678 1351
rect 3646 1332 3649 1338
rect 3662 1292 3665 1338
rect 3686 1302 3689 1318
rect 3702 1302 3705 1448
rect 3806 1421 3809 1459
rect 3806 1418 3817 1421
rect 3718 1372 3721 1418
rect 3814 1392 3817 1418
rect 3822 1402 3825 1468
rect 3798 1362 3801 1368
rect 3822 1352 3825 1388
rect 3838 1372 3841 1468
rect 3886 1462 3889 1528
rect 3898 1468 3902 1471
rect 3910 1462 3913 1518
rect 3934 1492 3937 1548
rect 3950 1472 3953 1618
rect 3958 1561 3961 1818
rect 3966 1662 3969 1848
rect 3974 1802 3977 1818
rect 3978 1788 3982 1791
rect 3982 1752 3985 1768
rect 3990 1742 3993 1748
rect 4006 1721 4009 2118
rect 4086 2072 4089 2078
rect 4066 2068 4070 2071
rect 4018 2058 4022 2061
rect 4022 1952 4025 1958
rect 4014 1762 4017 1788
rect 4022 1782 4025 1858
rect 4014 1732 4017 1758
rect 4030 1752 4033 1988
rect 4038 1952 4041 1958
rect 4046 1952 4049 2068
rect 4078 2052 4081 2058
rect 4102 2051 4105 2148
rect 4110 2122 4113 2148
rect 4112 2103 4114 2107
rect 4118 2103 4121 2107
rect 4125 2103 4128 2107
rect 4110 2072 4113 2078
rect 4110 2062 4113 2068
rect 4102 2048 4113 2051
rect 4066 2018 4070 2021
rect 4078 2012 4081 2048
rect 4094 1952 4097 2008
rect 4102 1982 4105 2018
rect 4110 1962 4113 2048
rect 4118 1992 4121 2078
rect 4126 2062 4129 2078
rect 4134 2072 4137 2208
rect 4150 2172 4153 2318
rect 4158 2272 4161 2418
rect 4174 2411 4177 2468
rect 4170 2408 4177 2411
rect 4166 2362 4169 2408
rect 4182 2392 4185 2648
rect 4198 2572 4201 2618
rect 4206 2592 4209 2658
rect 4214 2622 4217 2748
rect 4226 2738 4230 2741
rect 4230 2672 4233 2678
rect 4238 2632 4241 2748
rect 4246 2652 4249 2798
rect 4270 2762 4273 2858
rect 4254 2732 4257 2738
rect 4254 2692 4257 2718
rect 4294 2692 4297 2728
rect 4310 2672 4313 2888
rect 4326 2722 4329 2738
rect 4318 2682 4321 2688
rect 4334 2672 4337 2938
rect 4366 2892 4369 3138
rect 4398 3111 4401 3147
rect 4470 3142 4473 3228
rect 4486 3212 4489 3298
rect 4502 3262 4505 3268
rect 4514 3258 4518 3261
rect 4486 3172 4489 3208
rect 4506 3148 4510 3151
rect 4518 3142 4521 3148
rect 4390 3108 4401 3111
rect 4390 3092 4393 3108
rect 4378 3068 4382 3071
rect 4406 3062 4409 3068
rect 4374 3042 4377 3058
rect 4414 2952 4417 3138
rect 4494 3122 4497 3128
rect 4462 3102 4465 3118
rect 4422 3082 4425 3098
rect 4430 3062 4433 3068
rect 4454 3062 4457 3068
rect 4402 2948 4406 2951
rect 4414 2942 4417 2948
rect 4382 2872 4385 2938
rect 4406 2892 4409 2938
rect 4430 2881 4433 3058
rect 4466 3048 4470 3051
rect 4446 3042 4449 3048
rect 4478 3012 4481 3058
rect 4486 3012 4489 3068
rect 4494 3062 4497 3068
rect 4510 3052 4513 3098
rect 4518 3062 4521 3068
rect 4526 3062 4529 3258
rect 4566 3232 4569 3328
rect 4590 3322 4593 3348
rect 4614 3341 4617 3388
rect 4622 3352 4625 3428
rect 4632 3403 4634 3407
rect 4638 3403 4641 3407
rect 4645 3403 4648 3407
rect 4630 3362 4633 3368
rect 4610 3338 4617 3341
rect 4578 3318 4582 3321
rect 4598 3312 4601 3338
rect 4638 3312 4641 3378
rect 4578 3278 4582 3281
rect 4578 3268 4582 3271
rect 4534 3152 4537 3188
rect 4550 3152 4553 3218
rect 4534 3122 4537 3148
rect 4494 3042 4497 3048
rect 4518 3032 4521 3058
rect 4446 2932 4449 2938
rect 4422 2878 4433 2881
rect 4422 2862 4425 2878
rect 4442 2868 4446 2871
rect 4430 2862 4433 2868
rect 4454 2862 4457 2998
rect 4526 2982 4529 3018
rect 4534 3002 4537 3118
rect 4550 3072 4553 3148
rect 4566 3142 4569 3218
rect 4558 3082 4561 3118
rect 4574 3072 4577 3268
rect 4566 3052 4569 3058
rect 4478 2952 4481 2968
rect 4526 2951 4529 2958
rect 4542 2942 4545 3038
rect 4550 2972 4553 3048
rect 4574 3022 4577 3068
rect 4582 3052 4585 3078
rect 4590 3052 4593 3258
rect 4606 3252 4609 3278
rect 4638 3272 4641 3308
rect 4626 3258 4630 3261
rect 4638 3251 4641 3258
rect 4634 3248 4641 3251
rect 4606 3072 4609 3228
rect 4632 3203 4634 3207
rect 4638 3203 4641 3207
rect 4645 3203 4648 3207
rect 4654 3162 4657 3518
rect 4662 3442 4665 3538
rect 4678 3492 4681 3538
rect 4686 3482 4689 3548
rect 4694 3492 4697 3498
rect 4670 3462 4673 3478
rect 4702 3472 4705 3548
rect 4694 3392 4697 3468
rect 4682 3348 4686 3351
rect 4702 3342 4705 3468
rect 4710 3462 4713 3518
rect 4718 3462 4721 3468
rect 4726 3392 4729 3568
rect 4734 3552 4737 3698
rect 4774 3692 4777 3718
rect 4878 3691 4881 3788
rect 4926 3752 4929 3858
rect 4966 3752 4969 3818
rect 4982 3792 4985 3818
rect 4998 3782 5001 3848
rect 4994 3778 4998 3781
rect 4994 3758 4998 3761
rect 4986 3748 4990 3751
rect 4902 3732 4905 3748
rect 4870 3688 4881 3691
rect 4750 3672 4753 3678
rect 4774 3662 4777 3678
rect 4818 3668 4822 3671
rect 4774 3592 4777 3608
rect 4798 3592 4801 3668
rect 4830 3652 4833 3688
rect 4870 3672 4873 3688
rect 4882 3678 4886 3681
rect 4898 3668 4902 3671
rect 4910 3662 4913 3668
rect 4918 3662 4921 3708
rect 4958 3692 4961 3718
rect 4926 3682 4929 3688
rect 4850 3658 4854 3661
rect 4874 3658 4878 3661
rect 4818 3648 4822 3651
rect 4838 3642 4841 3648
rect 4758 3562 4761 3568
rect 4734 3532 4737 3538
rect 4742 3521 4745 3558
rect 4754 3548 4758 3551
rect 4734 3518 4745 3521
rect 4734 3492 4737 3518
rect 4750 3472 4753 3508
rect 4746 3458 4750 3461
rect 4758 3452 4761 3548
rect 4766 3462 4769 3468
rect 4774 3462 4777 3508
rect 4798 3482 4801 3488
rect 4786 3478 4790 3481
rect 4738 3448 4742 3451
rect 4758 3432 4761 3448
rect 4758 3352 4761 3358
rect 4714 3348 4718 3351
rect 4738 3348 4742 3351
rect 4750 3342 4753 3348
rect 4662 3322 4665 3328
rect 4662 3282 4665 3288
rect 4686 3162 4689 3198
rect 4614 3092 4617 3148
rect 4686 3142 4689 3148
rect 4662 3138 4670 3141
rect 4606 3052 4609 3058
rect 4598 3022 4601 3028
rect 4606 3022 4609 3048
rect 4614 3032 4617 3048
rect 4622 3042 4625 3128
rect 4654 3072 4657 3108
rect 4678 3082 4681 3098
rect 4638 3062 4641 3068
rect 4654 3062 4657 3068
rect 4630 3052 4633 3058
rect 4686 3041 4689 3118
rect 4694 3072 4697 3188
rect 4702 3182 4705 3338
rect 4766 3312 4769 3318
rect 4766 3282 4769 3288
rect 4742 3272 4745 3278
rect 4714 3258 4718 3261
rect 4774 3212 4777 3458
rect 4782 3352 4785 3358
rect 4798 3292 4801 3438
rect 4806 3392 4809 3638
rect 4846 3552 4849 3558
rect 4854 3542 4857 3618
rect 4870 3542 4873 3588
rect 4886 3542 4889 3548
rect 4854 3472 4857 3528
rect 4894 3462 4897 3578
rect 4902 3552 4905 3558
rect 4902 3462 4905 3468
rect 4910 3462 4913 3658
rect 4942 3592 4945 3638
rect 4926 3562 4929 3568
rect 4926 3502 4929 3548
rect 4934 3532 4937 3538
rect 4966 3522 4969 3738
rect 4974 3572 4977 3718
rect 4982 3662 4985 3668
rect 4850 3458 4854 3461
rect 4922 3458 4926 3461
rect 4846 3362 4849 3368
rect 4814 3348 4822 3351
rect 4850 3348 4854 3351
rect 4890 3348 4894 3351
rect 4806 3282 4809 3318
rect 4814 3262 4817 3348
rect 4826 3338 4830 3341
rect 4822 3272 4825 3328
rect 4786 3258 4790 3261
rect 4810 3258 4814 3261
rect 4702 3152 4705 3158
rect 4726 3152 4729 3168
rect 4798 3162 4801 3218
rect 4738 3158 4742 3161
rect 4782 3152 4785 3158
rect 4754 3138 4758 3141
rect 4778 3138 4782 3141
rect 4714 3128 4718 3131
rect 4718 3092 4721 3098
rect 4798 3082 4801 3118
rect 4814 3072 4817 3228
rect 4822 3152 4825 3258
rect 4830 3172 4833 3238
rect 4838 3202 4841 3258
rect 4846 3252 4849 3318
rect 4870 3302 4873 3318
rect 4866 3288 4870 3291
rect 4886 3282 4889 3338
rect 4698 3068 4702 3071
rect 4706 3058 4710 3061
rect 4678 3038 4689 3041
rect 4730 3038 4734 3041
rect 4610 2958 4614 2961
rect 4558 2942 4561 2948
rect 4574 2922 4577 2958
rect 4582 2942 4585 2958
rect 4598 2922 4601 2948
rect 4606 2932 4609 2938
rect 4462 2862 4465 2908
rect 4470 2862 4473 2868
rect 4518 2862 4521 2868
rect 4354 2858 4358 2861
rect 4442 2858 4446 2861
rect 4546 2858 4550 2861
rect 4458 2848 4462 2851
rect 4382 2792 4385 2808
rect 4478 2782 4481 2818
rect 4494 2812 4497 2858
rect 4510 2832 4513 2858
rect 4342 2711 4345 2747
rect 4342 2708 4353 2711
rect 4350 2692 4353 2708
rect 4374 2672 4377 2738
rect 4354 2668 4358 2671
rect 4190 2542 4193 2548
rect 4198 2512 4201 2548
rect 4206 2501 4209 2588
rect 4246 2551 4249 2558
rect 4254 2542 4257 2618
rect 4310 2592 4313 2668
rect 4334 2662 4337 2668
rect 4382 2662 4385 2718
rect 4398 2702 4401 2748
rect 4422 2722 4425 2728
rect 4422 2682 4425 2688
rect 4446 2672 4449 2738
rect 4462 2692 4465 2747
rect 4494 2672 4497 2768
rect 4526 2752 4529 2818
rect 4534 2762 4537 2798
rect 4558 2742 4561 2908
rect 4590 2862 4593 2888
rect 4614 2882 4617 2918
rect 4598 2862 4601 2868
rect 4566 2832 4569 2858
rect 4606 2822 4609 2868
rect 4574 2762 4577 2818
rect 4614 2762 4617 2858
rect 4582 2742 4585 2748
rect 4530 2718 4537 2721
rect 4534 2682 4537 2718
rect 4542 2712 4545 2738
rect 4590 2732 4593 2748
rect 4610 2738 4614 2741
rect 4562 2728 4566 2731
rect 4582 2692 4585 2728
rect 4598 2722 4601 2738
rect 4606 2692 4609 2728
rect 4622 2692 4625 3018
rect 4632 3003 4634 3007
rect 4638 3003 4641 3007
rect 4645 3003 4648 3007
rect 4654 3002 4657 3018
rect 4630 2852 4633 2938
rect 4654 2932 4657 2988
rect 4678 2952 4681 3038
rect 4774 3032 4777 3058
rect 4686 3022 4689 3028
rect 4702 2962 4705 3008
rect 4798 2992 4801 3068
rect 4814 3002 4817 3058
rect 4838 3052 4841 3088
rect 4814 2992 4817 2998
rect 4714 2968 4718 2971
rect 4686 2942 4689 2958
rect 4674 2938 4678 2941
rect 4698 2938 4702 2941
rect 4662 2912 4665 2918
rect 4678 2892 4681 2898
rect 4686 2882 4689 2918
rect 4670 2872 4673 2878
rect 4638 2852 4641 2868
rect 4662 2862 4665 2868
rect 4666 2858 4670 2861
rect 4632 2803 4634 2807
rect 4638 2803 4641 2807
rect 4645 2803 4648 2807
rect 4654 2792 4657 2828
rect 4646 2752 4649 2778
rect 4662 2762 4665 2818
rect 4670 2752 4673 2808
rect 4678 2742 4681 2748
rect 4686 2742 4689 2748
rect 4522 2668 4526 2671
rect 4362 2658 4366 2661
rect 4398 2652 4401 2658
rect 4382 2582 4385 2618
rect 4214 2532 4217 2538
rect 4206 2498 4214 2501
rect 4214 2462 4217 2498
rect 4194 2458 4198 2461
rect 4198 2362 4201 2418
rect 4226 2368 4230 2371
rect 4186 2348 4190 2351
rect 4202 2348 4206 2351
rect 4174 2302 4177 2318
rect 4190 2312 4193 2338
rect 4214 2332 4217 2358
rect 4246 2352 4249 2518
rect 4254 2472 4257 2538
rect 4262 2462 4265 2488
rect 4278 2351 4281 2368
rect 4238 2342 4241 2348
rect 4262 2332 4265 2338
rect 4202 2318 4206 2321
rect 4202 2288 4209 2291
rect 4194 2258 4198 2261
rect 4174 2212 4177 2218
rect 4206 2192 4209 2288
rect 4214 2252 4217 2328
rect 4222 2322 4225 2328
rect 4238 2292 4241 2318
rect 4286 2272 4289 2288
rect 4294 2272 4297 2568
rect 4406 2552 4409 2658
rect 4438 2642 4441 2668
rect 4446 2622 4449 2668
rect 4486 2662 4489 2668
rect 4454 2642 4457 2648
rect 4478 2642 4481 2658
rect 4346 2548 4350 2551
rect 4330 2538 4334 2541
rect 4310 2522 4313 2528
rect 4310 2462 4313 2488
rect 4318 2452 4321 2518
rect 4342 2502 4345 2548
rect 4342 2478 4358 2481
rect 4342 2471 4345 2478
rect 4326 2468 4345 2471
rect 4326 2462 4329 2468
rect 4338 2458 4342 2461
rect 4334 2442 4337 2448
rect 4342 2362 4345 2368
rect 4350 2352 4353 2468
rect 4366 2462 4369 2538
rect 4374 2462 4377 2468
rect 4374 2442 4377 2448
rect 4366 2392 4369 2408
rect 4382 2402 4385 2518
rect 4382 2352 4385 2378
rect 4362 2348 4366 2351
rect 4318 2282 4321 2308
rect 4330 2288 4334 2291
rect 4294 2262 4297 2268
rect 4342 2262 4345 2298
rect 4250 2258 4254 2261
rect 4282 2258 4286 2261
rect 4214 2232 4217 2238
rect 4254 2232 4257 2258
rect 4322 2248 4326 2251
rect 4262 2242 4265 2248
rect 4294 2242 4297 2248
rect 4278 2202 4281 2218
rect 4350 2202 4353 2348
rect 4358 2318 4366 2321
rect 4358 2292 4361 2318
rect 4366 2252 4369 2298
rect 4378 2268 4382 2271
rect 4390 2222 4393 2538
rect 4398 2452 4401 2468
rect 4406 2351 4409 2548
rect 4414 2481 4417 2518
rect 4422 2492 4425 2618
rect 4466 2578 4470 2581
rect 4458 2558 4462 2561
rect 4430 2552 4433 2558
rect 4442 2538 4446 2541
rect 4414 2478 4425 2481
rect 4402 2348 4409 2351
rect 4414 2342 4417 2468
rect 4422 2462 4425 2478
rect 4446 2462 4449 2468
rect 4454 2452 4457 2518
rect 4478 2492 4481 2638
rect 4494 2532 4497 2668
rect 4582 2662 4585 2688
rect 4590 2682 4593 2688
rect 4470 2462 4473 2478
rect 4478 2472 4481 2478
rect 4486 2462 4489 2498
rect 4510 2462 4513 2658
rect 4518 2652 4521 2658
rect 4566 2652 4569 2658
rect 4550 2572 4553 2618
rect 4574 2612 4577 2658
rect 4574 2562 4577 2578
rect 4582 2562 4585 2568
rect 4526 2542 4529 2547
rect 4542 2532 4545 2538
rect 4558 2502 4561 2538
rect 4582 2532 4585 2558
rect 4590 2542 4593 2668
rect 4614 2652 4617 2678
rect 4662 2672 4665 2688
rect 4678 2672 4681 2728
rect 4674 2668 4678 2671
rect 4622 2602 4625 2658
rect 4642 2648 4646 2651
rect 4632 2603 4634 2607
rect 4638 2603 4641 2607
rect 4645 2603 4648 2607
rect 4642 2568 4646 2571
rect 4618 2548 4622 2551
rect 4598 2542 4601 2548
rect 4618 2538 4622 2541
rect 4526 2478 4553 2481
rect 4526 2462 4529 2478
rect 4550 2472 4553 2478
rect 4534 2462 4537 2468
rect 4462 2452 4465 2458
rect 4470 2392 4473 2418
rect 4446 2352 4449 2388
rect 4470 2342 4473 2388
rect 4478 2352 4481 2358
rect 4486 2342 4489 2458
rect 4494 2452 4497 2458
rect 4546 2448 4550 2451
rect 4566 2451 4569 2518
rect 4582 2472 4585 2518
rect 4626 2488 4630 2491
rect 4638 2482 4641 2548
rect 4646 2482 4649 2488
rect 4662 2472 4665 2658
rect 4670 2652 4673 2658
rect 4686 2472 4689 2618
rect 4562 2448 4569 2451
rect 4602 2458 4606 2461
rect 4574 2442 4577 2458
rect 4678 2452 4681 2459
rect 4506 2428 4510 2431
rect 4546 2428 4550 2431
rect 4518 2372 4521 2398
rect 4506 2358 4510 2361
rect 4518 2352 4521 2368
rect 4538 2358 4542 2361
rect 4526 2352 4529 2358
rect 4458 2338 4462 2341
rect 4398 2292 4401 2328
rect 4414 2322 4417 2328
rect 4430 2322 4433 2328
rect 4422 2272 4425 2308
rect 4414 2232 4417 2258
rect 4330 2188 4334 2191
rect 4154 2158 4158 2161
rect 4190 2152 4193 2158
rect 4222 2152 4225 2158
rect 4178 2148 4182 2151
rect 4142 2142 4145 2148
rect 4166 2142 4169 2148
rect 4166 2092 4169 2128
rect 4174 2092 4177 2098
rect 4166 2052 4169 2078
rect 4082 1948 4086 1951
rect 4046 1942 4049 1948
rect 4102 1932 4105 1948
rect 4126 1932 4129 1948
rect 4054 1912 4057 1918
rect 4070 1902 4073 1928
rect 4112 1903 4114 1907
rect 4118 1903 4121 1907
rect 4125 1903 4128 1907
rect 4062 1882 4065 1888
rect 4042 1818 4046 1821
rect 4078 1792 4081 1888
rect 4102 1872 4105 1898
rect 4090 1868 4094 1871
rect 4038 1752 4041 1758
rect 4054 1742 4057 1788
rect 4086 1782 4089 1858
rect 4098 1848 4102 1851
rect 4094 1802 4097 1818
rect 4062 1752 4065 1778
rect 4006 1718 4017 1721
rect 3998 1712 4001 1718
rect 3982 1692 3985 1698
rect 4014 1692 4017 1718
rect 3990 1672 3993 1678
rect 3998 1662 4001 1678
rect 4022 1672 4025 1688
rect 3970 1638 3974 1641
rect 3958 1558 3969 1561
rect 3966 1552 3969 1558
rect 3974 1552 3977 1558
rect 3990 1552 3993 1658
rect 4030 1652 4033 1728
rect 4070 1692 4073 1698
rect 4086 1682 4089 1778
rect 4102 1752 4105 1848
rect 4114 1838 4118 1841
rect 4118 1732 4121 1738
rect 4102 1692 4105 1718
rect 4112 1703 4114 1707
rect 4118 1703 4121 1707
rect 4125 1703 4128 1707
rect 4050 1658 4054 1661
rect 4014 1552 4017 1638
rect 4062 1632 4065 1668
rect 4086 1662 4089 1678
rect 4022 1592 4025 1598
rect 4054 1562 4057 1588
rect 4050 1548 4054 1551
rect 3958 1542 3961 1548
rect 3990 1542 3993 1548
rect 3966 1492 3969 1508
rect 3958 1472 3961 1478
rect 3974 1472 3977 1518
rect 3998 1492 4001 1538
rect 3986 1488 3990 1491
rect 4002 1488 4009 1491
rect 3866 1458 3870 1461
rect 3890 1458 3894 1461
rect 3938 1458 3942 1461
rect 3866 1448 3873 1451
rect 3854 1432 3857 1448
rect 3854 1392 3857 1408
rect 3830 1352 3833 1358
rect 3754 1348 3758 1351
rect 3734 1332 3737 1348
rect 3838 1342 3841 1348
rect 3766 1292 3769 1338
rect 3794 1288 3798 1291
rect 3698 1268 3702 1271
rect 3558 1242 3561 1259
rect 3602 1258 3606 1261
rect 3646 1252 3649 1258
rect 3590 1242 3593 1248
rect 3606 1242 3609 1248
rect 3550 1082 3553 1138
rect 3558 1132 3561 1198
rect 3574 1152 3577 1228
rect 3582 1192 3585 1238
rect 3608 1203 3610 1207
rect 3614 1203 3617 1207
rect 3621 1203 3624 1207
rect 3646 1192 3649 1238
rect 3634 1148 3638 1151
rect 3598 1142 3601 1148
rect 3590 1072 3593 1098
rect 3590 1062 3593 1068
rect 3446 872 3449 878
rect 3446 852 3449 868
rect 3438 838 3449 841
rect 3438 792 3441 828
rect 3446 821 3449 838
rect 3454 831 3457 938
rect 3462 882 3465 948
rect 3470 942 3473 1038
rect 3478 962 3481 988
rect 3494 952 3497 958
rect 3502 952 3505 1008
rect 3502 892 3505 948
rect 3462 862 3465 878
rect 3470 872 3473 888
rect 3490 878 3494 881
rect 3454 828 3462 831
rect 3446 818 3457 821
rect 3454 792 3457 818
rect 3470 811 3473 868
rect 3482 858 3486 861
rect 3502 842 3505 868
rect 3470 808 3481 811
rect 3478 792 3481 808
rect 3430 778 3441 781
rect 3386 688 3390 691
rect 3414 672 3417 708
rect 3422 672 3425 748
rect 3430 742 3433 768
rect 3430 692 3433 728
rect 3438 662 3441 778
rect 3470 762 3473 768
rect 3446 692 3449 728
rect 3398 602 3401 638
rect 3366 562 3369 568
rect 3382 562 3385 598
rect 3430 592 3433 618
rect 3402 588 3406 591
rect 3438 582 3441 658
rect 3454 602 3457 618
rect 3374 552 3377 558
rect 3390 551 3393 568
rect 3438 562 3441 568
rect 3454 562 3457 598
rect 3382 548 3393 551
rect 3398 552 3401 558
rect 3454 552 3457 558
rect 3426 548 3430 551
rect 3442 548 3446 551
rect 3350 538 3361 541
rect 3270 472 3273 478
rect 3294 462 3297 468
rect 3126 452 3129 458
rect 3102 422 3105 438
rect 3150 402 3153 458
rect 3038 352 3041 398
rect 3174 392 3177 428
rect 3154 388 3158 391
rect 3030 342 3033 348
rect 3046 342 3049 378
rect 3274 368 3278 371
rect 3054 301 3057 358
rect 3094 342 3097 347
rect 3190 342 3193 348
rect 3046 298 3057 301
rect 2958 262 2961 268
rect 2982 262 2985 268
rect 3014 262 3017 288
rect 3002 258 3006 261
rect 3030 252 3033 278
rect 2934 248 2942 251
rect 3002 248 3014 251
rect 2918 198 2929 201
rect 2894 152 2897 188
rect 2918 162 2921 198
rect 2934 191 2937 238
rect 2930 188 2937 191
rect 2886 142 2889 148
rect 2890 88 2894 91
rect 2902 82 2905 158
rect 2918 132 2921 158
rect 2958 151 2961 218
rect 2958 148 2966 151
rect 2934 72 2937 148
rect 2974 142 2977 228
rect 3022 142 3025 238
rect 3022 132 3025 138
rect 2982 82 2985 88
rect 2942 62 2945 68
rect 2998 62 3001 68
rect 3014 52 3017 58
rect 3022 52 3025 78
rect 3038 62 3041 228
rect 3046 72 3049 298
rect 3062 292 3065 338
rect 3078 272 3081 338
rect 3126 332 3129 338
rect 3096 303 3098 307
rect 3102 303 3105 307
rect 3109 303 3112 307
rect 3126 292 3129 298
rect 3126 282 3129 288
rect 3150 272 3153 318
rect 3066 259 3070 262
rect 3054 62 3057 68
rect 3070 62 3073 238
rect 3078 192 3081 268
rect 3158 262 3161 328
rect 3166 302 3169 328
rect 3198 262 3201 288
rect 3206 272 3209 368
rect 3310 362 3313 368
rect 3278 358 3286 361
rect 3278 352 3281 358
rect 3218 348 3222 351
rect 3290 348 3294 351
rect 3274 338 3278 341
rect 3238 322 3241 338
rect 3326 332 3329 348
rect 3334 342 3337 518
rect 3342 392 3345 528
rect 3358 482 3361 538
rect 3366 492 3369 528
rect 3374 522 3377 538
rect 3382 492 3385 548
rect 3406 542 3409 548
rect 3450 538 3454 541
rect 3414 532 3417 538
rect 3422 492 3425 508
rect 3462 502 3465 728
rect 3470 672 3473 708
rect 3470 642 3473 668
rect 3478 662 3481 698
rect 3478 622 3481 658
rect 3486 632 3489 818
rect 3494 662 3497 668
rect 3502 652 3505 688
rect 3470 562 3473 568
rect 3486 561 3489 628
rect 3494 592 3497 648
rect 3510 622 3513 938
rect 3542 872 3545 1058
rect 3586 1038 3590 1041
rect 3598 1012 3601 1058
rect 3606 1052 3609 1148
rect 3618 1088 3622 1091
rect 3618 1078 3622 1081
rect 3614 1052 3617 1058
rect 3608 1003 3610 1007
rect 3614 1003 3617 1007
rect 3621 1003 3624 1007
rect 3610 988 3614 991
rect 3550 952 3553 958
rect 3638 952 3641 1058
rect 3646 1052 3649 1058
rect 3654 992 3657 1238
rect 3670 1222 3673 1258
rect 3726 1252 3729 1258
rect 3686 1242 3689 1248
rect 3726 1232 3729 1238
rect 3686 1192 3689 1228
rect 3662 1082 3665 1138
rect 3670 1122 3673 1148
rect 3694 1112 3697 1148
rect 3670 1072 3673 1088
rect 3686 1061 3689 1108
rect 3702 1091 3705 1178
rect 3710 1152 3713 1208
rect 3734 1202 3737 1268
rect 3742 1262 3745 1268
rect 3806 1262 3809 1288
rect 3822 1282 3825 1338
rect 3862 1322 3865 1348
rect 3870 1292 3873 1448
rect 3878 1362 3881 1458
rect 3886 1432 3889 1438
rect 3894 1381 3897 1458
rect 3918 1452 3921 1458
rect 3926 1441 3929 1448
rect 3906 1438 3929 1441
rect 3910 1392 3913 1428
rect 3886 1378 3897 1381
rect 3834 1288 3838 1291
rect 3878 1282 3881 1308
rect 3842 1278 3846 1281
rect 3818 1268 3822 1271
rect 3886 1262 3889 1378
rect 3894 1362 3897 1368
rect 3902 1352 3905 1388
rect 3926 1372 3929 1398
rect 3934 1392 3937 1458
rect 3970 1448 3974 1451
rect 3894 1272 3897 1278
rect 3902 1272 3905 1338
rect 3750 1242 3753 1258
rect 3774 1242 3777 1258
rect 3822 1252 3825 1258
rect 3846 1252 3849 1258
rect 3794 1248 3798 1251
rect 3718 1192 3721 1198
rect 3854 1192 3857 1258
rect 3878 1241 3881 1258
rect 3874 1238 3881 1241
rect 3742 1162 3745 1168
rect 3710 1122 3713 1128
rect 3710 1091 3713 1108
rect 3726 1101 3729 1158
rect 3758 1152 3761 1168
rect 3770 1158 3774 1161
rect 3822 1152 3825 1158
rect 3862 1152 3865 1158
rect 3870 1152 3873 1158
rect 3778 1148 3782 1151
rect 3834 1148 3838 1151
rect 3742 1142 3745 1148
rect 3750 1122 3753 1138
rect 3782 1132 3785 1138
rect 3702 1088 3713 1091
rect 3710 1082 3713 1088
rect 3718 1098 3729 1101
rect 3686 1058 3694 1061
rect 3698 1058 3702 1061
rect 3662 1042 3665 1048
rect 3690 1038 3694 1041
rect 3662 942 3665 948
rect 3522 748 3526 751
rect 3550 742 3553 938
rect 3638 932 3641 938
rect 3670 882 3673 1008
rect 3582 872 3585 878
rect 3670 872 3673 878
rect 3614 862 3617 868
rect 3678 862 3681 1018
rect 3718 992 3721 1098
rect 3730 1088 3734 1091
rect 3734 1062 3737 1068
rect 3742 1062 3745 1078
rect 3726 952 3729 1018
rect 3734 992 3737 998
rect 3686 882 3689 938
rect 3726 932 3729 938
rect 3718 882 3721 918
rect 3558 842 3561 858
rect 3566 742 3569 858
rect 3530 688 3534 691
rect 3526 672 3529 678
rect 3486 558 3497 561
rect 3482 548 3486 551
rect 3470 512 3473 518
rect 3390 472 3393 488
rect 3466 478 3470 481
rect 3434 468 3438 471
rect 3374 412 3377 438
rect 3398 432 3401 468
rect 3406 462 3409 468
rect 3446 452 3449 478
rect 3454 462 3457 468
rect 3478 432 3481 438
rect 3446 392 3449 398
rect 3486 372 3489 498
rect 3494 472 3497 558
rect 3502 471 3505 608
rect 3518 602 3521 658
rect 3526 652 3529 668
rect 3550 642 3553 738
rect 3518 582 3521 598
rect 3534 592 3537 638
rect 3566 602 3569 738
rect 3574 592 3577 818
rect 3608 803 3610 807
rect 3614 803 3617 807
rect 3621 803 3624 807
rect 3678 792 3681 838
rect 3686 772 3689 868
rect 3734 862 3737 868
rect 3694 752 3697 798
rect 3702 762 3705 858
rect 3710 852 3713 858
rect 3734 822 3737 858
rect 3742 792 3745 1038
rect 3758 1012 3761 1068
rect 3774 1063 3777 1088
rect 3754 958 3761 961
rect 3750 892 3753 948
rect 3758 892 3761 958
rect 3766 932 3769 958
rect 3782 952 3785 1038
rect 3790 1032 3793 1148
rect 3814 1122 3817 1148
rect 3838 1092 3841 1108
rect 3862 1092 3865 1128
rect 3870 1092 3873 1148
rect 3878 1132 3881 1158
rect 3902 1152 3905 1168
rect 3910 1162 3913 1258
rect 3918 1242 3921 1298
rect 3918 1202 3921 1238
rect 3918 1152 3921 1158
rect 3926 1152 3929 1348
rect 3942 1302 3945 1418
rect 3966 1352 3969 1358
rect 3974 1332 3977 1338
rect 3950 1262 3953 1328
rect 3990 1292 3993 1448
rect 3974 1282 3977 1288
rect 3934 1152 3937 1218
rect 3942 1192 3945 1198
rect 3982 1152 3985 1158
rect 3890 1148 3894 1151
rect 3902 1132 3905 1138
rect 3934 1132 3937 1138
rect 3886 1092 3889 1118
rect 3990 1081 3993 1218
rect 3998 1092 4001 1318
rect 4006 1292 4009 1488
rect 4022 1392 4025 1408
rect 4014 1322 4017 1348
rect 4030 1342 4033 1458
rect 4038 1412 4041 1548
rect 4054 1481 4057 1518
rect 4070 1502 4073 1618
rect 4110 1592 4113 1688
rect 4118 1662 4121 1678
rect 4078 1552 4081 1558
rect 4134 1552 4137 2008
rect 4158 1952 4161 1998
rect 4166 1972 4169 2048
rect 4190 1952 4193 1958
rect 4206 1952 4209 2028
rect 4214 2012 4217 2148
rect 4230 2132 4233 2158
rect 4254 2152 4257 2158
rect 4286 2152 4289 2168
rect 4230 2062 4233 2118
rect 4254 2082 4257 2148
rect 4302 2142 4305 2158
rect 4354 2148 4358 2151
rect 4262 2102 4265 2128
rect 4342 2112 4345 2148
rect 4370 2138 4374 2141
rect 4358 2102 4361 2138
rect 4238 1962 4241 2058
rect 4242 1958 4246 1961
rect 4222 1952 4225 1958
rect 4166 1941 4169 1948
rect 4158 1938 4169 1941
rect 4198 1942 4201 1948
rect 4158 1872 4161 1938
rect 4178 1928 4182 1931
rect 4206 1872 4209 1948
rect 4254 1942 4257 1968
rect 4286 1951 4289 1978
rect 4270 1942 4273 1948
rect 4294 1922 4297 2068
rect 4306 2058 4310 2061
rect 4350 1962 4353 1968
rect 4354 1928 4358 1931
rect 4366 1931 4369 2128
rect 4382 2072 4385 2078
rect 4390 2062 4393 2088
rect 4374 1942 4377 1988
rect 4382 1952 4385 2048
rect 4390 1992 4393 2028
rect 4366 1928 4377 1931
rect 4386 1928 4390 1931
rect 4166 1862 4169 1868
rect 4142 1842 4145 1848
rect 4150 1842 4153 1848
rect 4166 1842 4169 1858
rect 4174 1852 4177 1868
rect 4142 1752 4145 1758
rect 4190 1682 4193 1818
rect 4206 1782 4209 1858
rect 4214 1842 4217 1848
rect 4218 1788 4222 1791
rect 4218 1758 4222 1761
rect 4206 1751 4209 1758
rect 4206 1748 4222 1751
rect 4234 1748 4238 1751
rect 4246 1742 4249 1788
rect 4270 1752 4273 1878
rect 4278 1863 4281 1898
rect 4294 1872 4297 1918
rect 4318 1892 4321 1928
rect 4310 1852 4313 1878
rect 4342 1872 4345 1918
rect 4366 1902 4369 1918
rect 4326 1862 4329 1868
rect 4366 1862 4369 1868
rect 4278 1792 4281 1828
rect 4318 1792 4321 1808
rect 4366 1792 4369 1798
rect 4290 1758 4294 1761
rect 4302 1752 4305 1758
rect 4246 1728 4254 1731
rect 4206 1662 4209 1688
rect 4214 1672 4217 1718
rect 4222 1672 4225 1708
rect 4230 1662 4233 1688
rect 4142 1652 4145 1658
rect 4150 1652 4153 1658
rect 4246 1652 4249 1728
rect 4286 1712 4289 1718
rect 4286 1672 4289 1708
rect 4294 1702 4297 1728
rect 4310 1712 4313 1748
rect 4274 1668 4278 1671
rect 4294 1662 4297 1698
rect 4318 1662 4321 1688
rect 4162 1638 4166 1641
rect 4182 1592 4185 1598
rect 4122 1548 4126 1551
rect 4082 1538 4086 1541
rect 4094 1522 4097 1548
rect 4054 1478 4065 1481
rect 4062 1472 4065 1478
rect 4094 1472 4097 1498
rect 4102 1492 4105 1528
rect 4112 1503 4114 1507
rect 4118 1503 4121 1507
rect 4125 1503 4128 1507
rect 4134 1502 4137 1548
rect 4142 1542 4145 1548
rect 4150 1532 4153 1558
rect 4166 1552 4169 1588
rect 4166 1511 4169 1548
rect 4174 1522 4177 1538
rect 4166 1508 4177 1511
rect 4054 1462 4057 1468
rect 4102 1392 4105 1478
rect 4122 1448 4126 1451
rect 4050 1358 4054 1361
rect 4118 1352 4121 1358
rect 4126 1352 4129 1388
rect 4050 1348 4054 1351
rect 4098 1348 4105 1351
rect 4038 1342 4041 1348
rect 4030 1272 4033 1338
rect 4054 1332 4057 1338
rect 4070 1332 4073 1348
rect 4082 1338 4086 1341
rect 4046 1262 4049 1298
rect 4070 1272 4073 1278
rect 4086 1272 4089 1288
rect 4102 1272 4105 1348
rect 4112 1303 4114 1307
rect 4118 1303 4121 1307
rect 4125 1303 4128 1307
rect 4134 1272 4137 1438
rect 4142 1282 4145 1468
rect 4158 1463 4161 1468
rect 4150 1342 4153 1418
rect 4166 1332 4169 1358
rect 4162 1288 4166 1291
rect 4006 1142 4009 1238
rect 4094 1232 4097 1258
rect 4110 1242 4113 1248
rect 3990 1078 4001 1081
rect 3842 1068 3846 1071
rect 3930 1068 3934 1071
rect 3858 1058 3862 1061
rect 3962 1058 3966 1061
rect 3814 1018 3822 1021
rect 3814 992 3817 1018
rect 3798 962 3801 978
rect 3830 962 3833 968
rect 3802 948 3806 951
rect 3822 942 3825 948
rect 3774 932 3777 938
rect 3782 902 3785 908
rect 3754 868 3758 871
rect 3762 858 3766 861
rect 3774 852 3777 868
rect 3782 862 3785 898
rect 3798 892 3801 938
rect 3810 928 3814 931
rect 3806 872 3809 898
rect 3818 888 3822 891
rect 3838 872 3841 878
rect 3758 792 3761 848
rect 3798 822 3801 848
rect 3822 842 3825 848
rect 3782 792 3785 808
rect 3822 792 3825 818
rect 3766 752 3769 778
rect 3798 752 3801 778
rect 3706 748 3710 751
rect 3722 748 3726 751
rect 3778 748 3782 751
rect 3622 691 3625 718
rect 3614 688 3625 691
rect 3614 672 3617 688
rect 3586 658 3590 661
rect 3608 603 3610 607
rect 3614 603 3617 607
rect 3621 603 3624 607
rect 3526 562 3529 588
rect 3542 562 3545 588
rect 3522 548 3526 551
rect 3510 542 3513 548
rect 3550 542 3553 568
rect 3566 542 3569 558
rect 3578 548 3582 551
rect 3590 532 3593 578
rect 3622 552 3625 568
rect 3630 542 3633 548
rect 3510 482 3513 488
rect 3502 468 3513 471
rect 3498 458 3502 461
rect 3502 372 3505 378
rect 3454 362 3457 368
rect 3402 348 3406 351
rect 3454 342 3457 348
rect 3238 282 3241 318
rect 3334 302 3337 338
rect 3110 192 3113 248
rect 3158 182 3161 258
rect 3174 252 3177 258
rect 3142 152 3145 158
rect 3090 148 3094 151
rect 3096 103 3098 107
rect 3102 103 3105 107
rect 3109 103 3112 107
rect 3106 88 3110 91
rect 3166 82 3169 208
rect 3198 172 3201 218
rect 3222 192 3225 218
rect 3174 151 3177 168
rect 3206 152 3209 158
rect 3214 152 3217 168
rect 3238 142 3241 148
rect 3198 72 3201 108
rect 3230 92 3233 98
rect 3230 82 3233 88
rect 3246 72 3249 278
rect 3254 262 3257 298
rect 3326 292 3329 298
rect 3306 288 3310 291
rect 3318 272 3321 278
rect 3310 262 3313 268
rect 3342 262 3345 278
rect 3262 142 3265 258
rect 3286 152 3289 218
rect 3342 192 3345 248
rect 3350 162 3353 328
rect 3366 322 3369 338
rect 3358 282 3361 288
rect 3422 272 3425 298
rect 3438 292 3441 318
rect 3362 268 3366 271
rect 3350 92 3353 158
rect 3366 122 3369 258
rect 3394 248 3398 251
rect 3414 232 3417 258
rect 3430 252 3433 288
rect 3446 272 3449 308
rect 3462 291 3465 368
rect 3486 362 3489 368
rect 3474 348 3478 351
rect 3482 338 3486 341
rect 3458 288 3465 291
rect 3378 218 3382 221
rect 3470 212 3473 238
rect 3502 232 3505 348
rect 3510 342 3513 468
rect 3526 422 3529 518
rect 3550 451 3553 518
rect 3542 448 3553 451
rect 3518 362 3521 368
rect 3526 352 3529 418
rect 3542 352 3545 448
rect 3550 342 3553 438
rect 3566 432 3569 458
rect 3574 392 3577 518
rect 3582 512 3585 518
rect 3590 472 3593 488
rect 3606 441 3609 538
rect 3622 472 3625 508
rect 3638 492 3641 558
rect 3654 522 3657 748
rect 3686 742 3689 748
rect 3722 738 3726 741
rect 3726 662 3729 668
rect 3678 652 3681 658
rect 3670 481 3673 618
rect 3702 552 3705 658
rect 3734 592 3737 728
rect 3742 672 3745 708
rect 3750 662 3753 728
rect 3814 692 3817 758
rect 3822 692 3825 748
rect 3830 742 3833 758
rect 3838 742 3841 748
rect 3798 672 3801 678
rect 3846 672 3849 808
rect 3854 682 3857 758
rect 3742 622 3745 658
rect 3774 652 3777 658
rect 3750 642 3753 648
rect 3742 592 3745 608
rect 3734 572 3737 588
rect 3790 581 3793 658
rect 3786 578 3793 581
rect 3770 568 3774 571
rect 3758 562 3761 568
rect 3782 552 3785 578
rect 3790 562 3793 568
rect 3678 542 3681 548
rect 3790 542 3793 548
rect 3750 501 3753 528
rect 3782 512 3785 538
rect 3798 512 3801 668
rect 3846 662 3849 668
rect 3806 552 3809 608
rect 3814 592 3817 658
rect 3814 542 3817 568
rect 3822 552 3825 578
rect 3830 572 3833 578
rect 3838 571 3841 658
rect 3854 592 3857 658
rect 3862 642 3865 1038
rect 3870 862 3873 898
rect 3870 692 3873 838
rect 3878 792 3881 1058
rect 3902 1002 3905 1058
rect 3990 1052 3993 1068
rect 3918 1042 3921 1048
rect 3918 992 3921 1038
rect 3926 982 3929 1018
rect 3950 1012 3953 1018
rect 3942 962 3945 988
rect 3974 971 3977 1038
rect 3990 1002 3993 1048
rect 3998 992 4001 1078
rect 4014 1062 4017 1078
rect 4022 1062 4025 1158
rect 4038 1142 4041 1208
rect 4094 1192 4097 1228
rect 4082 1188 4086 1191
rect 4050 1158 4054 1161
rect 4106 1158 4110 1161
rect 4054 1142 4057 1148
rect 4070 1142 4073 1148
rect 4094 1132 4097 1148
rect 4126 1142 4129 1228
rect 4142 1182 4145 1218
rect 4142 1152 4145 1168
rect 4150 1162 4153 1248
rect 4174 1172 4177 1508
rect 4190 1482 4193 1648
rect 4246 1602 4249 1648
rect 4286 1642 4289 1658
rect 4270 1592 4273 1618
rect 4230 1392 4233 1558
rect 4246 1551 4249 1588
rect 4278 1542 4281 1618
rect 4286 1582 4289 1638
rect 4286 1552 4289 1578
rect 4302 1562 4305 1658
rect 4310 1571 4313 1638
rect 4318 1571 4321 1578
rect 4310 1568 4321 1571
rect 4310 1552 4313 1558
rect 4282 1538 4286 1541
rect 4238 1502 4241 1538
rect 4238 1492 4241 1498
rect 4262 1482 4265 1538
rect 4318 1531 4321 1568
rect 4314 1528 4321 1531
rect 4286 1492 4289 1528
rect 4250 1478 4254 1481
rect 4318 1472 4321 1498
rect 4326 1472 4329 1788
rect 4334 1752 4337 1788
rect 4350 1752 4353 1778
rect 4350 1662 4353 1748
rect 4366 1662 4369 1668
rect 4350 1562 4353 1588
rect 4358 1552 4361 1648
rect 4374 1592 4377 1928
rect 4398 1912 4401 2218
rect 4422 2212 4425 2268
rect 4430 2252 4433 2318
rect 4490 2288 4494 2291
rect 4470 2278 4478 2281
rect 4470 2262 4473 2278
rect 4502 2272 4505 2318
rect 4510 2292 4513 2338
rect 4538 2318 4542 2321
rect 4574 2292 4577 2438
rect 4590 2432 4593 2448
rect 4606 2442 4609 2448
rect 4632 2403 4634 2407
rect 4638 2403 4641 2407
rect 4645 2403 4648 2407
rect 4598 2342 4601 2348
rect 4478 2262 4481 2268
rect 4510 2262 4513 2288
rect 4590 2282 4593 2338
rect 4622 2332 4625 2338
rect 4650 2318 4654 2321
rect 4686 2282 4689 2458
rect 4462 2252 4465 2258
rect 4414 2132 4417 2138
rect 4406 2052 4409 2068
rect 4414 2052 4417 2088
rect 4414 2032 4417 2048
rect 4422 2012 4425 2208
rect 4438 2172 4441 2248
rect 4462 2232 4465 2238
rect 4502 2232 4505 2258
rect 4582 2242 4585 2258
rect 4446 2151 4449 2158
rect 4494 2152 4497 2158
rect 4526 2152 4529 2158
rect 4522 2148 4526 2151
rect 4462 2142 4465 2148
rect 4430 2072 4433 2098
rect 4438 2072 4441 2078
rect 4442 2058 4446 2061
rect 4446 2042 4449 2048
rect 4454 2002 4457 2088
rect 4470 2072 4473 2078
rect 4478 2062 4481 2148
rect 4486 2142 4489 2148
rect 4486 2072 4489 2138
rect 4506 2128 4510 2131
rect 4526 2128 4534 2131
rect 4518 2092 4521 2108
rect 4526 2072 4529 2128
rect 4538 2118 4545 2121
rect 4542 2072 4545 2118
rect 4582 2092 4585 2148
rect 4590 2142 4593 2278
rect 4686 2272 4689 2278
rect 4634 2258 4638 2261
rect 4646 2232 4649 2258
rect 4614 2092 4617 2228
rect 4632 2203 4634 2207
rect 4638 2203 4641 2207
rect 4645 2203 4648 2207
rect 4586 2068 4590 2071
rect 4470 1972 4473 1978
rect 4454 1962 4457 1968
rect 4438 1952 4441 1958
rect 4470 1952 4473 1958
rect 4418 1948 4422 1951
rect 4406 1912 4409 1938
rect 4382 1812 4385 1858
rect 4382 1752 4385 1758
rect 4382 1642 4385 1698
rect 4390 1692 4393 1898
rect 4422 1892 4425 1928
rect 4430 1922 4433 1928
rect 4430 1872 4433 1918
rect 4438 1902 4441 1938
rect 4462 1932 4465 1938
rect 4478 1892 4481 2058
rect 4486 1902 4489 2048
rect 4494 2042 4497 2068
rect 4502 2002 4505 2058
rect 4518 1992 4521 2038
rect 4494 1952 4497 1958
rect 4518 1952 4521 1988
rect 4450 1868 4454 1871
rect 4482 1868 4486 1871
rect 4430 1852 4433 1858
rect 4486 1852 4489 1858
rect 4458 1848 4462 1851
rect 4406 1742 4409 1828
rect 4414 1742 4417 1748
rect 4394 1668 4398 1671
rect 4390 1612 4393 1618
rect 4406 1581 4409 1738
rect 4414 1722 4417 1738
rect 4422 1732 4425 1748
rect 4414 1662 4417 1688
rect 4422 1632 4425 1638
rect 4430 1622 4433 1848
rect 4474 1768 4478 1771
rect 4438 1762 4441 1768
rect 4466 1758 4470 1761
rect 4494 1752 4497 1858
rect 4502 1792 4505 1818
rect 4470 1748 4478 1751
rect 4462 1702 4465 1748
rect 4470 1742 4473 1748
rect 4510 1702 4513 1938
rect 4526 1922 4529 2068
rect 4542 2052 4545 2068
rect 4566 2062 4569 2068
rect 4594 2058 4598 2061
rect 4566 1992 4569 2058
rect 4606 2052 4609 2068
rect 4622 2052 4625 2078
rect 4638 2032 4641 2158
rect 4662 2152 4665 2218
rect 4670 2152 4673 2258
rect 4686 2202 4689 2268
rect 4694 2262 4697 2898
rect 4718 2892 4721 2958
rect 4726 2862 4729 2978
rect 4766 2952 4769 2988
rect 4774 2892 4777 2968
rect 4790 2942 4793 2988
rect 4846 2952 4849 3178
rect 4854 3082 4857 3268
rect 4866 3248 4870 3251
rect 4878 3242 4881 3268
rect 4894 3262 4897 3338
rect 4902 3271 4905 3458
rect 4918 3442 4921 3448
rect 4950 3382 4953 3418
rect 4982 3381 4985 3498
rect 4990 3392 4993 3698
rect 5006 3672 5009 4018
rect 5014 3982 5017 4268
rect 5022 4242 5025 4248
rect 5070 4242 5073 4258
rect 5054 4172 5057 4178
rect 5082 4158 5086 4161
rect 5046 4142 5049 4158
rect 5058 4148 5062 4151
rect 5070 4151 5073 4158
rect 5070 4148 5081 4151
rect 5030 4132 5033 4138
rect 5030 4082 5033 4128
rect 5062 4121 5065 4148
rect 5062 4118 5073 4121
rect 5014 3951 5017 3958
rect 5030 3942 5033 4078
rect 5062 4072 5065 4098
rect 5070 4052 5073 4118
rect 5078 4092 5081 4148
rect 5086 4132 5089 4148
rect 5102 4142 5105 4268
rect 5118 4151 5121 4168
rect 5174 4142 5177 4218
rect 5182 4152 5185 4168
rect 5086 4052 5089 4068
rect 5046 3942 5049 3968
rect 5066 3948 5070 3951
rect 5054 3942 5057 3948
rect 5022 3872 5025 3908
rect 5014 3862 5017 3868
rect 5014 3762 5017 3818
rect 5030 3752 5033 3938
rect 5038 3752 5041 3758
rect 5038 3692 5041 3728
rect 5046 3672 5049 3938
rect 5070 3932 5073 3938
rect 5070 3861 5073 3928
rect 5078 3892 5081 3958
rect 5086 3872 5089 3978
rect 5094 3962 5097 4018
rect 5094 3922 5097 3948
rect 5102 3942 5105 4088
rect 5174 4072 5177 4138
rect 5110 3992 5113 3998
rect 5146 3958 5150 3961
rect 5094 3872 5097 3918
rect 5102 3912 5105 3938
rect 5118 3932 5121 3958
rect 5126 3942 5129 3948
rect 5134 3922 5137 3948
rect 5158 3942 5161 4059
rect 5174 3932 5177 3948
rect 5190 3942 5193 4508
rect 5086 3862 5089 3868
rect 5070 3858 5078 3861
rect 5054 3842 5057 3848
rect 5070 3822 5073 3858
rect 5078 3842 5081 3848
rect 5090 3828 5094 3831
rect 5090 3768 5094 3771
rect 5126 3762 5129 3858
rect 5150 3852 5153 3858
rect 5126 3752 5129 3758
rect 5078 3742 5081 3748
rect 5102 3692 5105 3738
rect 5054 3682 5057 3688
rect 5134 3682 5137 3768
rect 5158 3711 5161 3747
rect 5190 3712 5193 3938
rect 5158 3708 5169 3711
rect 5166 3692 5169 3708
rect 5022 3662 5025 3668
rect 5030 3662 5033 3668
rect 5054 3572 5057 3678
rect 5106 3668 5110 3671
rect 5170 3668 5174 3671
rect 5066 3658 5070 3661
rect 5078 3622 5081 3668
rect 5086 3662 5089 3668
rect 5150 3662 5153 3668
rect 5190 3662 5193 3708
rect 5014 3552 5017 3558
rect 5110 3552 5113 3658
rect 5014 3482 5017 3538
rect 5054 3482 5057 3548
rect 5062 3492 5065 3518
rect 5030 3462 5033 3468
rect 5006 3452 5009 3458
rect 4982 3378 4993 3381
rect 4934 3372 4937 3378
rect 4910 3362 4913 3368
rect 4938 3358 4942 3361
rect 4962 3358 4966 3361
rect 4918 3352 4921 3358
rect 4954 3348 4958 3351
rect 4918 3322 4921 3338
rect 4934 3281 4937 3318
rect 4930 3278 4937 3281
rect 4902 3268 4910 3271
rect 4910 3252 4913 3268
rect 4926 3262 4929 3268
rect 4934 3252 4937 3258
rect 4890 3248 4894 3251
rect 4886 3202 4889 3218
rect 4894 3152 4897 3248
rect 4910 3192 4913 3248
rect 4918 3172 4921 3178
rect 4934 3162 4937 3168
rect 4870 3142 4873 3148
rect 4918 3142 4921 3148
rect 4862 3062 4865 3118
rect 4874 3088 4878 3091
rect 4870 3062 4873 3068
rect 4862 3052 4865 3058
rect 4862 3032 4865 3038
rect 4870 2952 4873 2968
rect 4826 2948 4830 2951
rect 4838 2942 4841 2948
rect 4846 2942 4849 2948
rect 4866 2928 4870 2931
rect 4750 2882 4753 2888
rect 4738 2868 4742 2871
rect 4706 2858 4710 2861
rect 4726 2852 4729 2858
rect 4758 2802 4761 2878
rect 4798 2872 4801 2888
rect 4814 2862 4817 2868
rect 4854 2863 4857 2918
rect 4790 2842 4793 2858
rect 4742 2792 4745 2798
rect 4798 2752 4801 2758
rect 4738 2748 4742 2751
rect 4730 2738 4734 2741
rect 4806 2732 4809 2858
rect 4822 2852 4825 2858
rect 4838 2752 4841 2828
rect 4846 2792 4849 2818
rect 4878 2792 4881 3078
rect 4886 2992 4889 3088
rect 4894 3042 4897 3138
rect 4910 3112 4913 3138
rect 4942 3092 4945 3138
rect 4950 3122 4953 3348
rect 4962 3338 4966 3341
rect 4974 3292 4977 3358
rect 4990 3352 4993 3378
rect 5002 3368 5006 3371
rect 4958 3172 4961 3218
rect 4966 3162 4969 3198
rect 4982 3162 4985 3168
rect 4978 3148 4982 3151
rect 4990 3151 4993 3348
rect 4998 3342 5001 3348
rect 5046 3332 5049 3418
rect 5058 3348 5062 3351
rect 5062 3272 5065 3338
rect 5070 3332 5073 3538
rect 5078 3522 5081 3548
rect 5110 3542 5113 3548
rect 5090 3538 5094 3541
rect 5126 3532 5129 3638
rect 5134 3592 5137 3618
rect 5150 3602 5153 3658
rect 5150 3532 5153 3558
rect 5162 3538 5166 3541
rect 5086 3342 5089 3468
rect 5094 3462 5097 3518
rect 5126 3502 5129 3528
rect 5118 3362 5121 3488
rect 5134 3472 5137 3518
rect 5142 3362 5145 3528
rect 5150 3492 5153 3498
rect 5158 3482 5161 3518
rect 5154 3468 5158 3471
rect 5166 3462 5169 3528
rect 5158 3392 5161 3448
rect 5166 3432 5169 3458
rect 5178 3448 5182 3451
rect 5166 3372 5169 3418
rect 5174 3382 5177 3388
rect 5162 3358 5166 3361
rect 5110 3352 5113 3358
rect 5134 3342 5137 3348
rect 5106 3338 5110 3341
rect 4986 3148 4993 3151
rect 4998 3262 5001 3268
rect 5010 3258 5014 3261
rect 5090 3258 5094 3261
rect 4998 3152 5001 3258
rect 5094 3192 5097 3198
rect 5054 3152 5057 3158
rect 5030 3142 5033 3148
rect 4994 3138 4998 3141
rect 4994 3118 4998 3121
rect 4898 2948 4902 2951
rect 4902 2932 4905 2938
rect 4886 2882 4889 2918
rect 4910 2872 4913 3058
rect 4926 3042 4929 3058
rect 4958 3052 4961 3118
rect 5006 3092 5009 3138
rect 4990 3062 4993 3088
rect 5014 3082 5017 3118
rect 5046 3092 5049 3148
rect 5002 3068 5006 3071
rect 4974 3052 4977 3058
rect 4982 3012 4985 3058
rect 4990 2972 4993 2988
rect 4942 2942 4945 2968
rect 4966 2942 4969 2958
rect 4918 2892 4921 2928
rect 4886 2862 4889 2868
rect 4822 2742 4825 2748
rect 4838 2732 4841 2738
rect 4702 2672 4705 2728
rect 4862 2722 4865 2758
rect 4886 2742 4889 2858
rect 4910 2792 4913 2808
rect 4894 2752 4897 2758
rect 4902 2742 4905 2778
rect 4910 2732 4913 2748
rect 4718 2712 4721 2718
rect 4750 2662 4753 2708
rect 4774 2672 4777 2678
rect 4702 2261 4705 2558
rect 4710 2552 4713 2558
rect 4734 2542 4737 2658
rect 4790 2642 4793 2658
rect 4806 2622 4809 2628
rect 4826 2618 4830 2621
rect 4750 2552 4753 2608
rect 4766 2582 4769 2588
rect 4782 2552 4785 2558
rect 4754 2548 4758 2551
rect 4734 2532 4737 2538
rect 4782 2532 4785 2548
rect 4806 2542 4809 2548
rect 4814 2542 4817 2548
rect 4794 2538 4798 2541
rect 4838 2532 4841 2618
rect 4862 2592 4865 2658
rect 4738 2488 4742 2491
rect 4750 2472 4753 2498
rect 4750 2352 4753 2448
rect 4758 2432 4761 2458
rect 4758 2352 4761 2418
rect 4766 2392 4769 2518
rect 4814 2492 4817 2528
rect 4830 2491 4833 2528
rect 4846 2522 4849 2528
rect 4830 2488 4838 2491
rect 4782 2482 4785 2488
rect 4778 2448 4782 2451
rect 4770 2378 4774 2381
rect 4782 2352 4785 2358
rect 4710 2342 4713 2348
rect 4734 2332 4737 2338
rect 4734 2272 4737 2318
rect 4750 2272 4753 2338
rect 4790 2302 4793 2438
rect 4798 2422 4801 2458
rect 4822 2422 4825 2468
rect 4830 2462 4833 2478
rect 4838 2452 4841 2488
rect 4862 2482 4865 2548
rect 4850 2468 4854 2471
rect 4862 2462 4865 2468
rect 4870 2462 4873 2668
rect 4878 2572 4881 2718
rect 4918 2672 4921 2878
rect 4926 2802 4929 2818
rect 4926 2782 4929 2798
rect 4934 2761 4937 2918
rect 4950 2902 4953 2938
rect 4970 2918 4974 2921
rect 4958 2852 4961 2918
rect 5022 2902 5025 3068
rect 5062 3062 5065 3188
rect 5070 3072 5073 3078
rect 5078 3072 5081 3128
rect 5094 3072 5097 3178
rect 5062 3052 5065 3058
rect 5042 3048 5046 3051
rect 5090 3048 5094 3051
rect 5070 2982 5073 3048
rect 5070 2962 5073 2978
rect 5030 2952 5033 2958
rect 5054 2942 5057 2948
rect 5038 2882 5041 2888
rect 5050 2878 5054 2881
rect 5022 2872 5025 2878
rect 5070 2871 5073 2958
rect 5090 2948 5094 2951
rect 5090 2938 5097 2941
rect 5062 2868 5073 2871
rect 4974 2858 4982 2861
rect 4942 2782 4945 2788
rect 4930 2758 4937 2761
rect 4958 2732 4961 2748
rect 4966 2742 4969 2798
rect 4974 2792 4977 2858
rect 4982 2758 4990 2761
rect 4926 2692 4929 2718
rect 4942 2682 4945 2718
rect 4958 2702 4961 2728
rect 4966 2672 4969 2678
rect 4918 2622 4921 2668
rect 4934 2572 4937 2648
rect 4942 2632 4945 2668
rect 4974 2662 4977 2748
rect 4982 2692 4985 2758
rect 5022 2751 5025 2758
rect 4990 2692 4993 2738
rect 5022 2672 5025 2678
rect 5030 2662 5033 2758
rect 5054 2752 5057 2868
rect 5062 2862 5065 2868
rect 5070 2852 5073 2858
rect 5078 2852 5081 2918
rect 5086 2882 5089 2888
rect 5062 2682 5065 2708
rect 5070 2672 5073 2748
rect 5086 2712 5089 2718
rect 5058 2668 5062 2671
rect 5074 2668 5078 2671
rect 5002 2658 5006 2661
rect 5026 2658 5030 2661
rect 4958 2652 4961 2658
rect 4966 2641 4969 2658
rect 4982 2652 4985 2658
rect 5086 2652 5089 2668
rect 5034 2648 5038 2651
rect 5050 2648 5054 2651
rect 5066 2648 5070 2651
rect 4990 2641 4993 2648
rect 4966 2638 4993 2641
rect 4922 2568 4926 2571
rect 4878 2492 4881 2558
rect 4910 2552 4913 2558
rect 4886 2511 4889 2528
rect 4894 2522 4897 2528
rect 4886 2508 4897 2511
rect 4894 2492 4897 2508
rect 4878 2452 4881 2478
rect 4886 2472 4889 2478
rect 4850 2448 4854 2451
rect 4878 2442 4881 2448
rect 4854 2392 4857 2408
rect 4806 2362 4809 2368
rect 4826 2358 4830 2361
rect 4854 2352 4857 2378
rect 4886 2371 4889 2468
rect 4902 2462 4905 2538
rect 4910 2482 4913 2488
rect 4966 2462 4969 2518
rect 4974 2482 4977 2538
rect 4982 2502 4985 2547
rect 5046 2502 5049 2548
rect 5002 2488 5006 2491
rect 5054 2472 5057 2538
rect 5062 2462 5065 2548
rect 4902 2422 4905 2458
rect 4942 2452 4945 2458
rect 4878 2368 4889 2371
rect 4930 2368 4934 2371
rect 4878 2362 4881 2368
rect 4890 2358 4894 2361
rect 4802 2348 4806 2351
rect 4870 2342 4873 2358
rect 4894 2342 4897 2348
rect 4902 2342 4905 2358
rect 4982 2342 4985 2398
rect 5086 2372 5089 2648
rect 5094 2532 5097 2938
rect 5102 2792 5105 3328
rect 5110 3202 5113 3328
rect 5142 3322 5145 3338
rect 5150 3172 5153 3338
rect 5158 3292 5161 3318
rect 5166 3262 5169 3358
rect 5182 3332 5185 3438
rect 5186 3258 5190 3261
rect 5166 3192 5169 3258
rect 5186 3248 5190 3251
rect 5146 3148 5150 3151
rect 5126 3062 5129 3068
rect 5118 3052 5121 3058
rect 5118 2872 5121 2878
rect 5118 2732 5121 2748
rect 5126 2742 5129 2938
rect 5134 2872 5137 3148
rect 5142 3082 5145 3098
rect 5162 3058 5166 3061
rect 5142 2912 5145 3058
rect 5154 3048 5158 3051
rect 5174 3042 5177 3068
rect 5166 2942 5169 2948
rect 5174 2942 5177 2968
rect 5154 2938 5158 2941
rect 5138 2858 5142 2861
rect 5102 2602 5105 2718
rect 5110 2662 5113 2688
rect 5118 2582 5121 2618
rect 5126 2592 5129 2738
rect 5134 2672 5137 2688
rect 5158 2682 5161 2818
rect 5166 2692 5169 2928
rect 5182 2892 5185 2918
rect 5182 2792 5185 2868
rect 5182 2672 5185 2768
rect 5142 2652 5145 2658
rect 5166 2642 5169 2648
rect 5146 2618 5150 2621
rect 5102 2482 5105 2568
rect 5110 2562 5113 2568
rect 5126 2552 5129 2558
rect 5110 2542 5113 2548
rect 5150 2542 5153 2558
rect 5158 2552 5161 2558
rect 5134 2532 5137 2538
rect 5174 2532 5177 2568
rect 5146 2518 5150 2521
rect 5118 2482 5121 2518
rect 5138 2488 5142 2491
rect 5142 2462 5145 2468
rect 5150 2462 5153 2508
rect 5182 2502 5185 2658
rect 5190 2552 5193 2928
rect 5174 2492 5177 2498
rect 4990 2351 4993 2358
rect 4914 2338 4918 2341
rect 4798 2312 4801 2338
rect 4826 2318 4830 2321
rect 4838 2291 4841 2328
rect 4834 2288 4841 2291
rect 4834 2278 4838 2281
rect 4702 2258 4713 2261
rect 4698 2248 4702 2251
rect 4690 2178 4694 2181
rect 4710 2152 4713 2258
rect 4726 2252 4729 2258
rect 4726 2212 4729 2218
rect 4766 2212 4769 2259
rect 4734 2162 4737 2168
rect 4758 2152 4761 2168
rect 4658 2138 4662 2141
rect 4702 2122 4705 2148
rect 4646 2052 4649 2118
rect 4710 2092 4713 2148
rect 4750 2142 4753 2148
rect 4766 2142 4769 2148
rect 4774 2142 4777 2268
rect 4846 2262 4849 2338
rect 4854 2262 4857 2268
rect 4798 2242 4801 2258
rect 4790 2162 4793 2238
rect 4798 2221 4801 2228
rect 4798 2218 4809 2221
rect 4806 2192 4809 2218
rect 4802 2148 4806 2151
rect 4794 2138 4798 2141
rect 4718 2132 4721 2138
rect 4666 2068 4670 2071
rect 4662 2042 4665 2048
rect 4670 2032 4673 2058
rect 4702 2052 4705 2059
rect 4632 2003 4634 2007
rect 4638 2003 4641 2007
rect 4645 2003 4648 2007
rect 4542 1892 4545 1908
rect 4518 1842 4521 1858
rect 4526 1692 4529 1878
rect 4534 1862 4537 1868
rect 4550 1852 4553 1868
rect 4558 1822 4561 1848
rect 4566 1812 4569 1938
rect 4574 1862 4577 1928
rect 4582 1872 4585 1978
rect 4590 1872 4593 1968
rect 4650 1958 4654 1961
rect 4598 1951 4601 1958
rect 4638 1942 4641 1948
rect 4654 1942 4657 1948
rect 4614 1922 4617 1938
rect 4618 1878 4622 1881
rect 4574 1852 4577 1858
rect 4574 1832 4577 1838
rect 4566 1771 4569 1808
rect 4558 1768 4569 1771
rect 4534 1752 4537 1758
rect 4558 1742 4561 1768
rect 4574 1732 4577 1738
rect 4582 1722 4585 1818
rect 4598 1772 4601 1818
rect 4590 1762 4593 1768
rect 4606 1752 4609 1848
rect 4614 1752 4617 1758
rect 4606 1732 4609 1738
rect 4566 1692 4569 1718
rect 4474 1688 4478 1691
rect 4610 1688 4614 1691
rect 4446 1662 4449 1668
rect 4454 1662 4457 1668
rect 4502 1662 4505 1678
rect 4510 1662 4513 1678
rect 4534 1662 4537 1688
rect 4622 1672 4625 1878
rect 4632 1803 4634 1807
rect 4638 1803 4641 1807
rect 4645 1803 4648 1807
rect 4634 1778 4638 1781
rect 4642 1678 4646 1681
rect 4554 1668 4558 1671
rect 4602 1668 4606 1671
rect 4634 1668 4638 1671
rect 4654 1662 4657 1888
rect 4662 1802 4665 2028
rect 4678 1962 4681 2028
rect 4718 1992 4721 2118
rect 4734 2062 4737 2088
rect 4778 2068 4782 2071
rect 4726 2058 4734 2061
rect 4678 1942 4681 1958
rect 4710 1952 4713 1958
rect 4694 1942 4697 1948
rect 4702 1932 4705 1948
rect 4726 1922 4729 2058
rect 4790 2052 4793 2118
rect 4822 2092 4825 2258
rect 4830 2142 4833 2188
rect 4802 2058 4806 2061
rect 4810 2048 4814 2051
rect 4786 1968 4790 1971
rect 4734 1952 4737 1968
rect 4822 1962 4825 1968
rect 4770 1958 4774 1961
rect 4774 1942 4777 1948
rect 4750 1932 4753 1938
rect 4726 1872 4729 1918
rect 4742 1872 4745 1878
rect 4490 1658 4494 1661
rect 4570 1658 4574 1661
rect 4586 1658 4590 1661
rect 4438 1652 4441 1658
rect 4398 1578 4409 1581
rect 4346 1548 4350 1551
rect 4370 1548 4374 1551
rect 4334 1492 4337 1548
rect 4250 1468 4254 1471
rect 4326 1462 4329 1468
rect 4282 1458 4289 1461
rect 4254 1392 4257 1408
rect 4190 1362 4193 1368
rect 4230 1352 4233 1388
rect 4254 1362 4257 1388
rect 4186 1348 4190 1351
rect 4198 1342 4201 1348
rect 4206 1342 4209 1348
rect 4206 1292 4209 1328
rect 4246 1292 4249 1318
rect 4222 1263 4225 1288
rect 4238 1272 4241 1278
rect 4254 1262 4257 1308
rect 4262 1302 4265 1448
rect 4274 1338 4278 1341
rect 4270 1292 4273 1318
rect 4278 1302 4281 1318
rect 4262 1252 4265 1258
rect 4198 1162 4201 1178
rect 4214 1162 4217 1168
rect 4150 1148 4158 1151
rect 4210 1148 4214 1151
rect 4050 1118 4054 1121
rect 4034 1068 4038 1071
rect 4066 1068 4070 1071
rect 4050 1058 4054 1061
rect 4058 1048 4062 1051
rect 3966 968 3977 971
rect 3946 958 3953 961
rect 3886 952 3889 958
rect 3926 942 3929 948
rect 3886 872 3889 938
rect 3934 922 3937 938
rect 3922 888 3926 891
rect 3934 872 3937 918
rect 3878 752 3881 758
rect 3886 712 3889 868
rect 3894 662 3897 798
rect 3910 752 3913 768
rect 3902 682 3905 688
rect 3886 641 3889 658
rect 3910 651 3913 728
rect 3918 672 3921 868
rect 3934 862 3937 868
rect 3926 852 3929 858
rect 3942 772 3945 918
rect 3950 912 3953 958
rect 3950 872 3953 898
rect 3958 872 3961 918
rect 3966 892 3969 968
rect 3974 952 3977 958
rect 3982 932 3985 958
rect 3966 881 3969 888
rect 3966 878 3974 881
rect 3954 858 3958 861
rect 3982 832 3985 858
rect 3990 792 3993 978
rect 3998 892 4001 968
rect 4006 952 4009 958
rect 4014 952 4017 958
rect 3998 822 4001 828
rect 3982 752 3985 788
rect 4006 782 4009 948
rect 4022 941 4025 968
rect 4086 952 4089 1008
rect 4094 962 4097 968
rect 4074 948 4078 951
rect 4090 948 4097 951
rect 4018 938 4025 941
rect 4030 932 4033 938
rect 4038 932 4041 948
rect 4054 942 4057 948
rect 4074 938 4078 941
rect 4018 928 4022 931
rect 4078 882 4081 888
rect 4026 868 4030 871
rect 4054 862 4057 878
rect 4086 862 4089 908
rect 4014 832 4017 848
rect 4030 792 4033 858
rect 4014 752 4017 758
rect 4054 752 4057 818
rect 4062 762 4065 768
rect 4086 752 4089 858
rect 3930 748 3934 751
rect 3954 748 3958 751
rect 4066 748 4070 751
rect 3930 738 3934 741
rect 4022 741 4025 748
rect 4014 738 4025 741
rect 3930 728 3934 731
rect 3954 728 3958 731
rect 4002 728 4006 731
rect 3918 662 3921 668
rect 3910 648 3921 651
rect 3886 638 3897 641
rect 3862 592 3865 598
rect 3886 592 3889 628
rect 3846 571 3849 578
rect 3838 568 3849 571
rect 3846 562 3849 568
rect 3878 562 3881 568
rect 3862 542 3865 548
rect 3750 498 3761 501
rect 3662 478 3673 481
rect 3678 482 3681 488
rect 3598 438 3609 441
rect 3598 391 3601 438
rect 3608 403 3610 407
rect 3614 403 3617 407
rect 3621 403 3624 407
rect 3598 388 3606 391
rect 3574 352 3577 378
rect 3510 272 3513 338
rect 3554 328 3558 331
rect 3590 322 3593 358
rect 3630 351 3633 458
rect 3638 452 3641 478
rect 3638 392 3641 398
rect 3646 362 3649 468
rect 3654 462 3657 468
rect 3654 362 3657 398
rect 3630 348 3638 351
rect 3518 263 3521 318
rect 3598 292 3601 328
rect 3630 292 3633 338
rect 3630 282 3633 288
rect 3550 272 3553 278
rect 3534 242 3537 268
rect 3374 152 3377 198
rect 3526 192 3529 218
rect 3534 192 3537 238
rect 3558 232 3561 258
rect 3590 252 3593 258
rect 3418 158 3422 161
rect 3386 138 3390 141
rect 3398 102 3401 158
rect 3438 152 3441 188
rect 3454 152 3457 158
rect 3470 142 3473 178
rect 3494 172 3497 178
rect 3490 148 3494 151
rect 3410 138 3414 141
rect 3450 138 3454 141
rect 3258 88 3262 91
rect 3082 68 3086 71
rect 3210 68 3214 71
rect 3034 58 3038 61
rect 3198 62 3201 68
rect 3166 52 3169 59
rect 3050 48 3054 51
rect 3038 42 3041 48
rect 3214 32 3217 68
rect 3246 62 3249 68
rect 3318 63 3321 78
rect 3226 58 3230 61
rect 3382 62 3385 68
rect 3406 52 3409 58
rect 3422 52 3425 118
rect 3438 92 3441 98
rect 3446 82 3449 88
rect 3478 82 3481 88
rect 3474 68 3478 71
rect 3494 62 3497 108
rect 3502 72 3505 148
rect 3518 132 3521 168
rect 3466 58 3470 61
rect 3502 52 3505 58
rect 3510 52 3513 98
rect 3526 62 3529 188
rect 3534 72 3537 178
rect 3590 152 3593 228
rect 3598 142 3601 278
rect 3630 242 3633 258
rect 3638 232 3641 348
rect 3662 342 3665 478
rect 3742 472 3745 478
rect 3670 462 3673 468
rect 3734 462 3737 468
rect 3694 392 3697 398
rect 3686 362 3689 368
rect 3682 348 3686 351
rect 3730 348 3734 351
rect 3670 342 3673 348
rect 3742 342 3745 468
rect 3738 338 3742 341
rect 3670 302 3673 338
rect 3678 272 3681 338
rect 3662 263 3665 268
rect 3694 262 3697 268
rect 3710 262 3713 298
rect 3718 272 3721 278
rect 3726 272 3729 288
rect 3742 282 3745 338
rect 3750 302 3753 408
rect 3694 242 3697 248
rect 3608 203 3610 207
rect 3614 203 3617 207
rect 3621 203 3624 207
rect 3710 192 3713 258
rect 3726 222 3729 258
rect 3734 242 3737 248
rect 3638 162 3641 168
rect 3662 152 3665 188
rect 3674 168 3678 171
rect 3650 138 3654 141
rect 3590 132 3593 138
rect 3662 112 3665 148
rect 3670 122 3673 138
rect 3670 112 3673 118
rect 3634 88 3638 91
rect 3654 72 3657 78
rect 3662 62 3665 68
rect 3670 62 3673 68
rect 3578 58 3582 61
rect 3598 52 3601 58
rect 3686 52 3689 88
rect 3710 72 3713 178
rect 3726 142 3729 148
rect 3742 142 3745 278
rect 3750 262 3753 298
rect 3758 292 3761 498
rect 3806 472 3809 538
rect 3814 522 3817 538
rect 3822 512 3825 538
rect 3854 522 3857 538
rect 3886 512 3889 548
rect 3894 502 3897 638
rect 3906 578 3910 581
rect 3902 532 3905 538
rect 3846 472 3849 478
rect 3778 468 3782 471
rect 3774 452 3777 458
rect 3790 422 3793 458
rect 3790 342 3793 388
rect 3798 381 3801 468
rect 3806 392 3809 468
rect 3826 458 3830 461
rect 3866 459 3870 462
rect 3814 412 3817 458
rect 3830 432 3833 448
rect 3862 392 3865 428
rect 3798 378 3809 381
rect 3798 342 3801 348
rect 3786 288 3790 291
rect 3758 262 3761 268
rect 3778 258 3782 261
rect 3754 248 3758 251
rect 3778 248 3782 251
rect 3782 192 3785 238
rect 3798 152 3801 338
rect 3806 272 3809 378
rect 3834 368 3838 371
rect 3814 362 3817 368
rect 3846 362 3849 368
rect 3878 362 3881 498
rect 3814 342 3817 348
rect 3822 342 3825 358
rect 3858 348 3862 351
rect 3814 152 3817 158
rect 3790 142 3793 148
rect 3822 142 3825 338
rect 3830 222 3833 348
rect 3878 342 3881 348
rect 3854 322 3857 338
rect 3838 282 3841 308
rect 3838 272 3841 278
rect 3842 258 3846 261
rect 3830 152 3833 218
rect 3854 182 3857 318
rect 3886 262 3889 388
rect 3918 372 3921 648
rect 3926 542 3929 728
rect 3974 722 3977 728
rect 3942 692 3945 718
rect 3966 672 3969 708
rect 3938 668 3942 671
rect 3934 652 3937 658
rect 3926 522 3929 538
rect 3926 492 3929 498
rect 3934 482 3937 488
rect 3942 371 3945 668
rect 3950 662 3953 668
rect 3958 552 3961 598
rect 3966 542 3969 668
rect 3982 652 3985 659
rect 4014 592 4017 738
rect 4046 692 4049 698
rect 4070 692 4073 718
rect 4054 672 4057 688
rect 4078 682 4081 688
rect 4070 642 4073 648
rect 4086 632 4089 748
rect 4094 632 4097 948
rect 4102 851 4105 1138
rect 4112 1103 4114 1107
rect 4118 1103 4121 1107
rect 4125 1103 4128 1107
rect 4138 1058 4142 1061
rect 4112 903 4114 907
rect 4118 903 4121 907
rect 4125 903 4128 907
rect 4130 888 4134 891
rect 4122 858 4126 861
rect 4102 848 4110 851
rect 4134 751 4137 758
rect 4102 732 4105 738
rect 4112 703 4114 707
rect 4118 703 4121 707
rect 4125 703 4128 707
rect 4134 662 4137 728
rect 4070 572 4073 578
rect 4094 572 4097 618
rect 4106 558 4110 561
rect 4010 548 4014 551
rect 4006 521 4009 538
rect 3998 518 4009 521
rect 3986 488 3990 491
rect 3950 462 3953 478
rect 3974 472 3977 478
rect 3962 468 3966 471
rect 3982 442 3985 458
rect 3934 368 3945 371
rect 3934 352 3937 368
rect 3966 351 3969 358
rect 3894 272 3897 278
rect 3902 272 3905 318
rect 3910 282 3913 338
rect 3918 332 3921 338
rect 3918 292 3921 328
rect 3934 282 3937 348
rect 3950 312 3953 338
rect 3998 312 4001 518
rect 4030 512 4033 558
rect 4042 548 4046 551
rect 4054 532 4057 548
rect 4062 542 4065 548
rect 4090 538 4094 541
rect 4054 522 4057 528
rect 4046 482 4049 518
rect 4094 492 4097 508
rect 4112 503 4114 507
rect 4118 503 4121 507
rect 4125 503 4128 507
rect 4038 462 4041 468
rect 4030 392 4033 398
rect 4034 348 4038 351
rect 3910 252 3913 258
rect 3858 168 3862 171
rect 3842 148 3846 151
rect 3814 132 3817 138
rect 3774 102 3777 128
rect 3822 102 3825 138
rect 3706 58 3710 61
rect 3718 52 3721 58
rect 3442 48 3446 51
rect 3482 48 3486 51
rect 3790 32 3793 68
rect 3854 62 3857 68
rect 3870 62 3873 68
rect 3886 52 3889 148
rect 3910 142 3913 148
rect 3950 142 3953 258
rect 3958 192 3961 308
rect 4014 272 4017 328
rect 4046 292 4049 478
rect 4086 472 4089 478
rect 4134 472 4137 658
rect 4142 551 4145 998
rect 4150 592 4153 1148
rect 4166 1132 4169 1138
rect 4190 1092 4193 1148
rect 4174 1072 4177 1078
rect 4222 1071 4225 1138
rect 4218 1068 4225 1071
rect 4206 1062 4209 1068
rect 4230 1062 4233 1188
rect 4246 1092 4249 1218
rect 4218 1058 4222 1061
rect 4238 1048 4246 1051
rect 4190 1042 4193 1048
rect 4214 952 4217 968
rect 4162 948 4166 951
rect 4214 942 4217 948
rect 4190 922 4193 938
rect 4214 872 4217 918
rect 4238 892 4241 1048
rect 4254 1022 4257 1068
rect 4262 892 4265 1238
rect 4286 1132 4289 1458
rect 4302 1452 4305 1458
rect 4310 1432 4313 1458
rect 4326 1442 4329 1448
rect 4294 1262 4297 1288
rect 4302 1282 4305 1298
rect 4310 1182 4313 1428
rect 4334 1422 4337 1488
rect 4350 1452 4353 1458
rect 4342 1392 4345 1448
rect 4358 1372 4361 1548
rect 4390 1532 4393 1548
rect 4398 1542 4401 1578
rect 4414 1571 4417 1578
rect 4410 1568 4417 1571
rect 4398 1502 4401 1538
rect 4386 1488 4390 1491
rect 4366 1472 4369 1478
rect 4390 1452 4393 1468
rect 4398 1462 4401 1498
rect 4406 1472 4409 1488
rect 4390 1382 4393 1448
rect 4326 1282 4329 1338
rect 4334 1292 4337 1348
rect 4374 1292 4377 1318
rect 4358 1282 4361 1288
rect 4390 1282 4393 1288
rect 4318 1232 4321 1258
rect 4302 1152 4305 1158
rect 4326 1142 4329 1278
rect 4342 1232 4345 1268
rect 4354 1258 4358 1261
rect 4378 1258 4382 1261
rect 4354 1248 4358 1251
rect 4382 1192 4385 1198
rect 4342 1162 4345 1168
rect 4354 1158 4361 1161
rect 4310 1092 4313 1128
rect 4310 1082 4313 1088
rect 4326 1072 4329 1078
rect 4342 1071 4345 1158
rect 4358 1142 4361 1158
rect 4366 1152 4369 1188
rect 4406 1152 4409 1268
rect 4414 1252 4417 1258
rect 4414 1152 4417 1248
rect 4422 1222 4425 1378
rect 4430 1292 4433 1348
rect 4438 1342 4441 1458
rect 4446 1402 4449 1658
rect 4462 1632 4465 1658
rect 4558 1648 4566 1651
rect 4578 1648 4582 1651
rect 4462 1552 4465 1558
rect 4462 1462 4465 1488
rect 4486 1482 4489 1538
rect 4486 1472 4489 1478
rect 4502 1472 4505 1518
rect 4526 1492 4529 1548
rect 4510 1412 4513 1458
rect 4534 1452 4537 1618
rect 4550 1472 4553 1568
rect 4558 1492 4561 1648
rect 4570 1548 4574 1551
rect 4562 1488 4566 1491
rect 4574 1472 4577 1538
rect 4534 1412 4537 1448
rect 4542 1432 4545 1458
rect 4574 1442 4577 1468
rect 4438 1272 4441 1298
rect 4462 1272 4465 1318
rect 4470 1292 4473 1328
rect 4478 1292 4481 1388
rect 4518 1352 4521 1378
rect 4542 1362 4545 1428
rect 4486 1332 4489 1348
rect 4522 1338 4526 1341
rect 4510 1332 4513 1338
rect 4486 1292 4489 1298
rect 4450 1248 4454 1251
rect 4422 1152 4425 1218
rect 4462 1192 4465 1268
rect 4502 1262 4505 1318
rect 4542 1271 4545 1318
rect 4574 1311 4577 1328
rect 4582 1322 4585 1348
rect 4566 1308 4577 1311
rect 4598 1312 4601 1648
rect 4606 1592 4609 1648
rect 4646 1642 4649 1658
rect 4654 1642 4657 1648
rect 4632 1603 4634 1607
rect 4638 1603 4641 1607
rect 4645 1603 4648 1607
rect 4614 1542 4617 1568
rect 4634 1558 4638 1561
rect 4614 1462 4617 1478
rect 4622 1472 4625 1518
rect 4622 1372 4625 1468
rect 4632 1403 4634 1407
rect 4638 1403 4641 1407
rect 4645 1403 4648 1407
rect 4654 1402 4657 1588
rect 4662 1562 4665 1798
rect 4678 1711 4681 1868
rect 4710 1842 4713 1859
rect 4718 1732 4721 1748
rect 4726 1742 4729 1868
rect 4750 1852 4753 1858
rect 4766 1852 4769 1918
rect 4782 1912 4785 1948
rect 4806 1942 4809 1948
rect 4826 1938 4830 1941
rect 4798 1882 4801 1898
rect 4778 1868 4782 1871
rect 4750 1832 4753 1838
rect 4774 1812 4777 1868
rect 4774 1772 4777 1778
rect 4758 1762 4761 1768
rect 4782 1761 4785 1818
rect 4790 1811 4793 1848
rect 4806 1822 4809 1938
rect 4838 1882 4841 2218
rect 4850 2158 4854 2161
rect 4850 2138 4854 2141
rect 4862 2132 4865 2258
rect 4878 2092 4881 2218
rect 4886 2172 4889 2238
rect 4918 2152 4921 2158
rect 4926 2131 4929 2338
rect 4934 2272 4937 2278
rect 4946 2268 4950 2271
rect 4934 2262 4937 2268
rect 4966 2252 4969 2258
rect 4966 2152 4969 2248
rect 4950 2132 4953 2138
rect 4926 2128 4937 2131
rect 4918 2072 4921 2078
rect 4934 2072 4937 2128
rect 4966 2122 4969 2138
rect 4958 2118 4966 2121
rect 4958 2082 4961 2118
rect 4974 2072 4977 2218
rect 4982 2172 4985 2338
rect 5038 2332 5041 2368
rect 5110 2362 5113 2438
rect 5070 2352 5073 2358
rect 5054 2342 5057 2348
rect 5102 2342 5105 2348
rect 5090 2338 5094 2341
rect 5050 2328 5054 2331
rect 5082 2328 5086 2331
rect 5110 2331 5113 2358
rect 5118 2352 5121 2458
rect 5158 2452 5161 2458
rect 5102 2328 5113 2331
rect 5126 2342 5129 2448
rect 5134 2362 5137 2368
rect 5126 2332 5129 2338
rect 5022 2292 5025 2328
rect 5070 2321 5073 2328
rect 5070 2318 5081 2321
rect 5030 2312 5033 2318
rect 5006 2262 5009 2278
rect 5054 2272 5057 2288
rect 4998 2132 5001 2148
rect 4990 2092 4993 2108
rect 4894 2052 4897 2058
rect 4934 2022 4937 2068
rect 4974 2062 4977 2068
rect 4942 2042 4945 2048
rect 4950 2032 4953 2048
rect 4890 1978 4894 1981
rect 4850 1958 4854 1961
rect 4874 1958 4878 1961
rect 4866 1948 4870 1951
rect 4854 1892 4857 1898
rect 4934 1872 4937 1938
rect 4814 1852 4817 1858
rect 4838 1852 4841 1868
rect 4950 1862 4953 2018
rect 4958 1952 4961 1958
rect 4982 1942 4985 2078
rect 4994 2068 4998 2071
rect 5006 2062 5009 2248
rect 5030 2232 5033 2258
rect 5014 2072 5017 2168
rect 5022 2112 5025 2148
rect 5030 2082 5033 2228
rect 5054 2092 5057 2118
rect 5062 2102 5065 2318
rect 5070 2272 5073 2308
rect 5078 2302 5081 2318
rect 5078 2262 5081 2288
rect 5086 2272 5089 2278
rect 5094 2252 5097 2298
rect 5102 2292 5105 2328
rect 5134 2322 5137 2338
rect 5110 2302 5113 2318
rect 5102 2252 5105 2278
rect 5114 2268 5118 2271
rect 5082 2148 5086 2151
rect 5070 2072 5073 2118
rect 5038 2062 5041 2068
rect 5046 2062 5049 2068
rect 5066 2058 5070 2061
rect 5006 2022 5009 2058
rect 5022 2012 5025 2018
rect 5022 1972 5025 1978
rect 4958 1872 4961 1918
rect 4966 1892 4969 1908
rect 4982 1891 4985 1938
rect 4998 1922 5001 1948
rect 5006 1892 5009 1918
rect 4982 1888 4993 1891
rect 4974 1882 4977 1888
rect 4990 1872 4993 1888
rect 4846 1852 4849 1858
rect 4822 1832 4825 1838
rect 4838 1832 4841 1848
rect 4790 1808 4801 1811
rect 4782 1758 4790 1761
rect 4726 1732 4729 1738
rect 4782 1722 4785 1738
rect 4678 1708 4689 1711
rect 4686 1692 4689 1708
rect 4678 1672 4681 1678
rect 4670 1662 4673 1668
rect 4702 1662 4705 1688
rect 4710 1672 4713 1718
rect 4718 1662 4721 1668
rect 4758 1662 4761 1708
rect 4766 1662 4769 1668
rect 4754 1658 4758 1661
rect 4734 1652 4737 1658
rect 4790 1652 4793 1748
rect 4798 1712 4801 1808
rect 4810 1758 4814 1761
rect 4806 1712 4809 1748
rect 4818 1738 4822 1741
rect 4814 1702 4817 1738
rect 4830 1732 4833 1778
rect 4862 1751 4865 1768
rect 4846 1732 4849 1738
rect 4826 1718 4830 1721
rect 4762 1648 4766 1651
rect 4686 1632 4689 1648
rect 4734 1622 4737 1648
rect 4674 1558 4678 1561
rect 4662 1551 4665 1558
rect 4662 1548 4670 1551
rect 4710 1551 4713 1558
rect 4678 1542 4681 1548
rect 4694 1522 4697 1538
rect 4694 1482 4697 1488
rect 4674 1468 4678 1471
rect 4686 1452 4689 1458
rect 4710 1452 4713 1458
rect 4686 1442 4689 1448
rect 4662 1351 4665 1438
rect 4670 1362 4673 1368
rect 4678 1361 4681 1418
rect 4678 1358 4686 1361
rect 4662 1348 4670 1351
rect 4658 1338 4662 1341
rect 4566 1272 4569 1308
rect 4606 1292 4609 1318
rect 4638 1282 4641 1318
rect 4582 1272 4585 1278
rect 4542 1268 4553 1271
rect 4538 1258 4542 1261
rect 4470 1162 4473 1168
rect 4478 1152 4481 1238
rect 4550 1192 4553 1268
rect 4566 1262 4569 1268
rect 4622 1252 4625 1258
rect 4594 1248 4598 1251
rect 4632 1203 4634 1207
rect 4638 1203 4641 1207
rect 4645 1203 4648 1207
rect 4662 1192 4665 1238
rect 4490 1158 4494 1161
rect 4510 1152 4513 1158
rect 4518 1152 4521 1158
rect 4442 1148 4446 1151
rect 4498 1148 4502 1151
rect 4530 1148 4534 1151
rect 4374 1142 4377 1148
rect 4334 1068 4345 1071
rect 4334 1062 4337 1068
rect 4326 1058 4334 1061
rect 4326 962 4329 1058
rect 4342 1052 4345 1058
rect 4350 1052 4353 1118
rect 4398 1102 4401 1148
rect 4406 1122 4409 1148
rect 4422 1142 4425 1148
rect 4462 1132 4465 1148
rect 4362 1068 4366 1071
rect 4390 992 4393 1088
rect 4414 992 4417 1128
rect 4422 1062 4425 1068
rect 4430 1062 4433 1118
rect 4470 1092 4473 1148
rect 4482 1138 4486 1141
rect 4454 1072 4457 1078
rect 4390 962 4393 968
rect 4398 962 4401 978
rect 4346 958 4350 961
rect 4326 952 4329 958
rect 4350 952 4353 958
rect 4414 952 4417 958
rect 4454 952 4457 978
rect 4478 961 4481 1118
rect 4518 1112 4521 1138
rect 4546 1128 4550 1131
rect 4574 1092 4577 1158
rect 4598 1152 4601 1168
rect 4626 1158 4630 1161
rect 4646 1152 4649 1178
rect 4670 1162 4673 1348
rect 4718 1342 4721 1538
rect 4742 1502 4745 1538
rect 4726 1482 4729 1488
rect 4734 1452 4737 1468
rect 4742 1462 4745 1498
rect 4766 1492 4769 1508
rect 4750 1462 4753 1478
rect 4758 1452 4761 1458
rect 4774 1411 4777 1628
rect 4786 1548 4790 1551
rect 4798 1472 4801 1698
rect 4806 1622 4809 1678
rect 4870 1672 4873 1848
rect 4910 1842 4913 1858
rect 4950 1852 4953 1858
rect 4958 1832 4961 1868
rect 5014 1862 5017 1868
rect 4886 1672 4889 1788
rect 4922 1778 4926 1781
rect 4930 1758 4934 1761
rect 4894 1692 4897 1758
rect 4950 1752 4953 1768
rect 5018 1748 5022 1751
rect 4934 1742 4937 1748
rect 4962 1738 4966 1741
rect 4910 1692 4913 1738
rect 4962 1718 4966 1721
rect 4918 1682 4921 1718
rect 4950 1672 4953 1688
rect 4958 1672 4961 1688
rect 4974 1682 4977 1728
rect 5014 1672 5017 1738
rect 4842 1658 4846 1661
rect 4806 1552 4809 1618
rect 4838 1592 4841 1638
rect 4846 1562 4849 1648
rect 4870 1602 4873 1668
rect 4934 1658 4942 1661
rect 4806 1462 4809 1548
rect 4814 1532 4817 1538
rect 4822 1522 4825 1558
rect 4846 1552 4849 1558
rect 4854 1552 4857 1588
rect 4878 1582 4881 1588
rect 4894 1572 4897 1598
rect 4902 1592 4905 1648
rect 4926 1642 4929 1648
rect 4830 1542 4833 1548
rect 4830 1472 4833 1538
rect 4846 1472 4849 1498
rect 4862 1492 4865 1518
rect 4886 1492 4889 1508
rect 4878 1482 4881 1488
rect 4894 1472 4897 1548
rect 4910 1492 4913 1608
rect 4934 1562 4937 1658
rect 4942 1642 4945 1648
rect 5002 1548 5006 1551
rect 4934 1512 4937 1548
rect 4974 1542 4977 1548
rect 4982 1542 4985 1548
rect 4858 1468 4862 1471
rect 4902 1462 4905 1468
rect 4926 1462 4929 1478
rect 4934 1472 4937 1478
rect 4942 1472 4945 1478
rect 4958 1472 4961 1538
rect 4798 1458 4806 1461
rect 4782 1422 4785 1458
rect 4798 1412 4801 1458
rect 4810 1448 4814 1451
rect 4850 1448 4854 1451
rect 4822 1442 4825 1448
rect 4830 1432 4833 1448
rect 4774 1408 4785 1411
rect 4734 1351 4737 1358
rect 4698 1338 4702 1341
rect 4702 1322 4705 1328
rect 4710 1292 4713 1298
rect 4734 1292 4737 1308
rect 4758 1292 4761 1398
rect 4702 1272 4705 1278
rect 4750 1272 4753 1278
rect 4766 1272 4769 1408
rect 4782 1292 4785 1408
rect 4814 1352 4817 1428
rect 4838 1361 4841 1418
rect 4834 1358 4841 1361
rect 4826 1348 4830 1351
rect 4806 1342 4809 1348
rect 4794 1318 4798 1321
rect 4722 1268 4726 1271
rect 4682 1258 4686 1261
rect 4698 1248 4702 1251
rect 4746 1248 4750 1251
rect 4790 1242 4793 1248
rect 4726 1232 4729 1238
rect 4678 1152 4681 1218
rect 4586 1148 4590 1151
rect 4634 1148 4638 1151
rect 4658 1148 4662 1151
rect 4694 1151 4697 1158
rect 4710 1152 4713 1158
rect 4694 1148 4702 1151
rect 4602 1138 4606 1141
rect 4698 1138 4702 1141
rect 4662 1082 4665 1088
rect 4626 1078 4630 1081
rect 4566 1072 4569 1078
rect 4514 1058 4518 1061
rect 4474 958 4481 961
rect 4282 947 4286 950
rect 4338 948 4342 951
rect 4450 948 4454 951
rect 4466 948 4470 951
rect 4362 938 4366 941
rect 4378 938 4382 941
rect 4278 892 4281 928
rect 4302 922 4305 938
rect 4318 932 4321 938
rect 4442 928 4446 931
rect 4478 922 4481 928
rect 4230 872 4233 878
rect 4246 872 4249 878
rect 4302 872 4305 898
rect 4310 882 4313 888
rect 4310 862 4313 878
rect 4186 858 4190 861
rect 4254 852 4257 858
rect 4282 848 4289 851
rect 4190 692 4193 848
rect 4254 762 4257 838
rect 4270 761 4273 848
rect 4286 792 4289 848
rect 4294 822 4297 858
rect 4350 792 4353 888
rect 4374 882 4377 918
rect 4374 852 4377 859
rect 4282 768 4289 771
rect 4270 758 4281 761
rect 4214 732 4217 758
rect 4254 752 4257 758
rect 4234 748 4238 751
rect 4210 728 4214 731
rect 4206 662 4209 688
rect 4222 682 4225 738
rect 4270 732 4273 738
rect 4246 702 4249 718
rect 4250 678 4254 681
rect 4222 671 4225 678
rect 4218 668 4225 671
rect 4158 642 4161 659
rect 4218 658 4222 661
rect 4194 648 4198 651
rect 4182 592 4185 638
rect 4190 582 4193 628
rect 4206 592 4209 648
rect 4278 632 4281 758
rect 4238 612 4241 618
rect 4286 591 4289 768
rect 4330 758 4334 761
rect 4294 752 4297 758
rect 4306 748 4310 751
rect 4294 712 4297 738
rect 4310 692 4313 748
rect 4318 662 4321 698
rect 4326 672 4329 708
rect 4350 682 4353 778
rect 4374 752 4377 788
rect 4390 761 4393 918
rect 4414 872 4417 908
rect 4406 862 4409 868
rect 4438 862 4441 908
rect 4474 888 4478 891
rect 4450 878 4454 881
rect 4458 868 4462 871
rect 4486 862 4489 988
rect 4514 948 4518 951
rect 4526 942 4529 1068
rect 4578 1058 4582 1061
rect 4590 1051 4593 1078
rect 4586 1048 4593 1051
rect 4598 1062 4601 1068
rect 4634 1058 4638 1061
rect 4526 922 4529 938
rect 4542 892 4545 968
rect 4574 942 4577 1018
rect 4494 862 4497 878
rect 4526 872 4529 888
rect 4558 872 4561 938
rect 4566 862 4569 888
rect 4578 878 4582 881
rect 4554 858 4558 861
rect 4422 852 4425 858
rect 4438 782 4441 858
rect 4474 848 4478 851
rect 4502 812 4505 818
rect 4526 792 4529 858
rect 4590 852 4593 858
rect 4386 758 4393 761
rect 4398 752 4401 758
rect 4362 748 4366 751
rect 4386 748 4390 751
rect 4438 751 4441 758
rect 4510 752 4513 768
rect 4398 732 4401 748
rect 4374 692 4377 728
rect 4366 672 4369 678
rect 4406 672 4409 738
rect 4414 692 4417 718
rect 4422 712 4425 738
rect 4518 722 4521 748
rect 4502 712 4505 718
rect 4466 688 4470 691
rect 4282 588 4289 591
rect 4166 562 4169 568
rect 4142 548 4150 551
rect 4162 538 4169 541
rect 4070 412 4073 468
rect 4158 462 4161 508
rect 4166 452 4169 538
rect 4182 482 4185 548
rect 4190 542 4193 578
rect 4190 502 4193 538
rect 4198 482 4201 558
rect 4270 552 4273 588
rect 4234 548 4238 551
rect 4262 542 4265 548
rect 4206 538 4214 541
rect 4222 491 4225 528
rect 4254 512 4257 518
rect 4218 488 4225 491
rect 4222 462 4225 468
rect 4074 368 4078 371
rect 4062 342 4065 348
rect 4062 322 4065 338
rect 4070 292 4073 348
rect 4102 322 4105 448
rect 4182 412 4185 458
rect 4230 442 4233 498
rect 4254 492 4257 498
rect 4238 482 4241 488
rect 4262 472 4265 478
rect 4258 468 4262 471
rect 4270 462 4273 548
rect 4278 492 4281 518
rect 4318 502 4321 548
rect 4326 542 4329 668
rect 4390 662 4393 668
rect 4422 662 4425 678
rect 4438 672 4441 688
rect 4478 682 4481 708
rect 4486 692 4489 698
rect 4454 672 4457 678
rect 4542 672 4545 688
rect 4434 668 4438 671
rect 4446 662 4449 668
rect 4402 658 4406 661
rect 4382 642 4385 648
rect 4374 542 4377 598
rect 4414 592 4417 658
rect 4534 652 4537 658
rect 4466 648 4470 651
rect 4390 562 4393 568
rect 4402 558 4409 561
rect 4450 558 4454 561
rect 4310 462 4313 468
rect 4334 462 4337 538
rect 4370 488 4374 491
rect 4374 462 4377 468
rect 4134 351 4137 358
rect 4150 342 4153 408
rect 4170 368 4174 371
rect 4198 362 4201 368
rect 4210 358 4214 361
rect 4194 348 4198 351
rect 4210 348 4214 351
rect 4112 303 4114 307
rect 4118 303 4121 307
rect 4125 303 4128 307
rect 4046 272 4049 288
rect 4026 268 4030 271
rect 4014 262 4017 268
rect 4046 262 4049 268
rect 3974 252 3977 258
rect 4014 192 4017 258
rect 4054 251 4057 268
rect 4126 262 4129 268
rect 4106 258 4110 261
rect 4042 248 4057 251
rect 4054 192 4057 198
rect 3974 142 3977 148
rect 3998 132 4001 148
rect 3950 92 3953 128
rect 3982 82 3985 108
rect 3982 72 3985 78
rect 3906 58 3910 61
rect 3958 52 3961 68
rect 3990 62 3993 68
rect 4006 62 4009 88
rect 4014 72 4017 98
rect 4022 72 4025 98
rect 4022 62 4025 68
rect 4030 62 4033 98
rect 4046 72 4049 148
rect 4062 142 4065 188
rect 4070 152 4073 178
rect 4094 172 4097 198
rect 4142 172 4145 188
rect 4166 172 4169 348
rect 4202 338 4206 341
rect 4230 341 4233 438
rect 4238 352 4241 418
rect 4230 338 4238 341
rect 4242 318 4246 321
rect 4186 278 4190 281
rect 4194 268 4198 271
rect 4178 248 4182 251
rect 4198 172 4201 258
rect 4206 232 4209 268
rect 4230 252 4233 318
rect 4238 292 4241 308
rect 4262 272 4265 428
rect 4270 402 4273 458
rect 4334 412 4337 458
rect 4362 438 4369 441
rect 4342 352 4345 358
rect 4286 312 4289 348
rect 4294 282 4297 338
rect 4214 242 4217 248
rect 4238 242 4241 248
rect 4214 192 4217 218
rect 4142 152 4145 168
rect 4070 102 4073 148
rect 4110 142 4113 148
rect 4118 142 4121 148
rect 4166 142 4169 168
rect 4194 158 4198 161
rect 4174 142 4177 158
rect 4230 152 4233 228
rect 4254 182 4257 258
rect 4262 212 4265 268
rect 4278 262 4281 268
rect 4254 172 4257 178
rect 4238 152 4241 168
rect 4254 152 4257 158
rect 4294 152 4297 278
rect 4302 262 4305 308
rect 4326 151 4329 158
rect 4214 142 4217 148
rect 4230 142 4233 148
rect 4246 142 4249 148
rect 4162 138 4166 141
rect 4078 132 4081 138
rect 4222 132 4225 138
rect 4112 103 4114 107
rect 4118 103 4121 107
rect 4125 103 4128 107
rect 4190 92 4193 118
rect 4050 68 4054 71
rect 4062 62 4065 88
rect 4190 72 4193 88
rect 4198 82 4201 108
rect 4230 102 4233 128
rect 4342 112 4345 348
rect 4350 342 4353 348
rect 4350 292 4353 338
rect 4358 312 4361 318
rect 4358 292 4361 298
rect 4366 292 4369 438
rect 4374 332 4377 448
rect 4382 422 4385 518
rect 4390 472 4393 538
rect 4398 472 4401 518
rect 4406 492 4409 558
rect 4414 542 4417 548
rect 4422 542 4425 548
rect 4446 542 4449 548
rect 4430 532 4433 538
rect 4442 468 4446 471
rect 4430 462 4433 468
rect 4454 462 4457 468
rect 4450 458 4454 461
rect 4422 452 4425 458
rect 4406 392 4409 448
rect 4414 442 4417 448
rect 4410 368 4414 371
rect 4390 332 4393 368
rect 4402 348 4406 351
rect 4374 292 4377 328
rect 4406 312 4409 348
rect 4422 332 4425 448
rect 4430 372 4433 408
rect 4366 252 4369 278
rect 4390 268 4398 271
rect 4382 262 4385 268
rect 4390 232 4393 268
rect 4406 262 4409 298
rect 4462 292 4465 638
rect 4478 542 4481 548
rect 4470 482 4473 488
rect 4478 472 4481 518
rect 4486 492 4489 648
rect 4494 532 4497 548
rect 4526 511 4529 547
rect 4542 542 4545 668
rect 4518 508 4529 511
rect 4550 522 4553 838
rect 4590 792 4593 838
rect 4586 748 4590 751
rect 4558 732 4561 748
rect 4574 742 4577 748
rect 4598 742 4601 1058
rect 4614 1042 4617 1048
rect 4694 1042 4697 1058
rect 4710 1042 4713 1148
rect 4726 1112 4729 1118
rect 4718 1052 4721 1058
rect 4606 862 4609 868
rect 4614 862 4617 908
rect 4622 872 4625 1008
rect 4632 1003 4634 1007
rect 4638 1003 4641 1007
rect 4645 1003 4648 1007
rect 4634 988 4638 991
rect 4654 872 4657 1038
rect 4678 992 4681 1028
rect 4702 952 4705 998
rect 4734 962 4737 988
rect 4742 962 4745 1188
rect 4774 1132 4777 1238
rect 4794 1228 4798 1231
rect 4806 1172 4809 1338
rect 4814 1262 4817 1348
rect 4834 1338 4838 1341
rect 4870 1312 4873 1438
rect 4902 1352 4905 1458
rect 4914 1448 4918 1451
rect 4942 1372 4945 1468
rect 4990 1463 4993 1518
rect 4950 1442 4953 1448
rect 4958 1432 4961 1448
rect 4950 1352 4953 1358
rect 4890 1348 4894 1351
rect 4894 1292 4897 1308
rect 4878 1272 4881 1278
rect 4934 1272 4937 1338
rect 4814 1191 4817 1238
rect 4814 1188 4825 1191
rect 4798 1142 4801 1148
rect 4822 1142 4825 1188
rect 4758 1062 4761 1068
rect 4718 952 4721 958
rect 4674 948 4678 951
rect 4730 948 4734 951
rect 4694 942 4697 948
rect 4714 938 4718 941
rect 4726 882 4729 888
rect 4702 872 4705 878
rect 4750 872 4753 1038
rect 4774 1022 4777 1028
rect 4790 1012 4793 1068
rect 4806 1052 4809 1078
rect 4822 1071 4825 1138
rect 4838 1132 4841 1228
rect 4854 1152 4857 1218
rect 4862 1192 4865 1259
rect 4950 1222 4953 1338
rect 4966 1301 4969 1318
rect 4982 1312 4985 1328
rect 4958 1298 4969 1301
rect 4958 1263 4961 1298
rect 4974 1272 4977 1278
rect 4990 1272 4993 1358
rect 4998 1352 5001 1508
rect 5014 1472 5017 1668
rect 5022 1663 5025 1708
rect 5030 1702 5033 2038
rect 5046 1992 5049 2058
rect 5078 1962 5081 2148
rect 5086 2118 5094 2121
rect 5086 2082 5089 2118
rect 5086 2062 5089 2078
rect 5094 2072 5097 2078
rect 5102 2022 5105 2248
rect 5110 2082 5113 2218
rect 5118 2082 5121 2088
rect 5126 2061 5129 2288
rect 5142 2252 5145 2448
rect 5150 2372 5153 2428
rect 5166 2422 5169 2468
rect 5174 2352 5177 2468
rect 5150 2292 5153 2348
rect 5182 2341 5185 2478
rect 5174 2338 5185 2341
rect 5134 2222 5137 2228
rect 5134 2152 5137 2218
rect 5158 2182 5161 2338
rect 5118 2058 5129 2061
rect 5134 2062 5137 2128
rect 5150 2122 5153 2148
rect 5146 2068 5150 2071
rect 5110 2052 5113 2058
rect 5054 1872 5057 1948
rect 5078 1912 5081 1948
rect 5086 1892 5089 2018
rect 5118 1952 5121 2058
rect 5102 1872 5105 1878
rect 5054 1842 5057 1868
rect 5118 1862 5121 1948
rect 5126 1942 5129 1988
rect 5134 1862 5137 1918
rect 5142 1892 5145 2058
rect 5150 2042 5153 2048
rect 5150 1952 5153 1988
rect 5166 1942 5169 2098
rect 5174 2092 5177 2338
rect 5182 2212 5185 2328
rect 5190 2262 5193 2268
rect 5178 2068 5182 2071
rect 5174 2052 5177 2058
rect 5182 1992 5185 2038
rect 5174 1932 5177 1938
rect 5166 1882 5169 1928
rect 5062 1742 5065 1808
rect 5078 1762 5081 1798
rect 5102 1792 5105 1848
rect 5102 1752 5105 1758
rect 5166 1752 5169 1858
rect 5134 1742 5137 1748
rect 5114 1738 5118 1741
rect 5154 1738 5158 1741
rect 5114 1728 5118 1731
rect 5078 1682 5081 1688
rect 5054 1672 5057 1678
rect 5070 1652 5073 1658
rect 5054 1552 5057 1648
rect 5062 1562 5065 1618
rect 5074 1558 5078 1561
rect 5074 1548 5078 1551
rect 5022 1532 5025 1548
rect 5058 1538 5062 1541
rect 5090 1538 5094 1541
rect 5046 1532 5049 1538
rect 5022 1492 5025 1528
rect 5034 1518 5038 1521
rect 5050 1488 5054 1491
rect 5058 1468 5062 1471
rect 5070 1462 5073 1528
rect 5134 1512 5137 1738
rect 5174 1732 5177 1908
rect 5182 1792 5185 1978
rect 5190 1972 5193 2078
rect 5190 1892 5193 1958
rect 5186 1748 5190 1751
rect 5150 1712 5153 1718
rect 5150 1642 5153 1658
rect 5146 1548 5150 1551
rect 5158 1542 5161 1668
rect 5090 1488 5094 1491
rect 5158 1482 5161 1538
rect 5086 1462 5089 1468
rect 5066 1458 5070 1461
rect 5138 1458 5142 1461
rect 5022 1442 5025 1458
rect 5090 1448 5094 1451
rect 5126 1442 5129 1458
rect 5086 1392 5089 1428
rect 5006 1352 5009 1358
rect 4998 1342 5001 1348
rect 5030 1342 5033 1378
rect 5058 1358 5062 1361
rect 5038 1352 5041 1358
rect 5126 1352 5129 1438
rect 5138 1348 5142 1351
rect 5054 1342 5057 1348
rect 5018 1338 5022 1341
rect 5014 1332 5017 1338
rect 5034 1328 5038 1331
rect 5014 1292 5017 1298
rect 5030 1262 5033 1268
rect 5038 1262 5041 1268
rect 4990 1152 4993 1258
rect 5006 1252 5009 1258
rect 5014 1252 5017 1258
rect 4998 1161 5001 1218
rect 4998 1158 5006 1161
rect 4922 1148 4926 1151
rect 4970 1148 4974 1151
rect 5002 1148 5006 1151
rect 4878 1142 4881 1148
rect 4886 1142 4889 1148
rect 4934 1142 4937 1148
rect 4982 1142 4985 1148
rect 4906 1138 4910 1141
rect 5010 1138 5014 1141
rect 4894 1122 4897 1128
rect 4918 1122 4921 1138
rect 4830 1092 4833 1098
rect 4870 1092 4873 1118
rect 4882 1088 4886 1091
rect 4862 1082 4865 1088
rect 4902 1072 4905 1118
rect 4822 1068 4833 1071
rect 4814 1062 4817 1068
rect 4798 992 4801 1018
rect 4758 962 4761 968
rect 4762 948 4766 951
rect 4770 938 4774 941
rect 4782 932 4785 968
rect 4814 951 4817 958
rect 4762 888 4766 891
rect 4638 862 4641 868
rect 4606 792 4609 858
rect 4622 848 4630 851
rect 4558 702 4561 728
rect 4566 682 4569 718
rect 4582 672 4585 678
rect 4598 662 4601 728
rect 4606 672 4609 738
rect 4622 692 4625 848
rect 4632 803 4634 807
rect 4638 803 4641 807
rect 4645 803 4648 807
rect 4654 772 4657 868
rect 4662 842 4665 858
rect 4678 752 4681 868
rect 4738 858 4742 861
rect 4686 842 4689 848
rect 4710 842 4713 858
rect 4750 842 4753 868
rect 4750 772 4753 838
rect 4758 832 4761 858
rect 4798 752 4801 948
rect 4814 872 4817 928
rect 4822 922 4825 1058
rect 4830 882 4833 1068
rect 4850 1058 4854 1061
rect 4878 1052 4881 1058
rect 4926 1052 4929 1138
rect 4874 968 4878 971
rect 4890 958 4894 961
rect 4898 948 4902 951
rect 4886 942 4889 948
rect 4910 942 4913 958
rect 4926 952 4929 1048
rect 4870 892 4873 908
rect 4862 872 4865 878
rect 4818 858 4822 861
rect 4806 752 4809 828
rect 4762 748 4766 751
rect 4734 742 4737 748
rect 4798 742 4801 748
rect 4862 742 4865 748
rect 4678 692 4681 738
rect 4654 672 4657 678
rect 4618 668 4622 671
rect 4586 658 4590 661
rect 4606 622 4609 658
rect 4646 622 4649 648
rect 4632 603 4634 607
rect 4638 603 4641 607
rect 4645 603 4648 607
rect 4558 532 4561 548
rect 4598 542 4601 578
rect 4670 572 4673 648
rect 4686 592 4689 738
rect 4694 662 4697 708
rect 4710 692 4713 698
rect 4742 682 4745 718
rect 4758 702 4761 728
rect 4734 672 4737 678
rect 4766 672 4769 738
rect 4790 732 4793 738
rect 4774 722 4777 728
rect 4810 718 4814 721
rect 4862 692 4865 698
rect 4782 672 4785 688
rect 4870 672 4873 758
rect 4702 642 4705 668
rect 4730 658 4734 661
rect 4762 658 4766 661
rect 4750 652 4753 658
rect 4714 648 4718 651
rect 4654 562 4657 568
rect 4626 558 4630 561
rect 4650 548 4654 551
rect 4606 542 4609 548
rect 4642 538 4646 541
rect 4518 492 4521 508
rect 4550 482 4553 518
rect 4510 472 4513 478
rect 4534 462 4537 478
rect 4582 472 4585 528
rect 4590 512 4593 518
rect 4622 512 4625 518
rect 4502 452 4505 458
rect 4494 442 4497 448
rect 4510 362 4513 368
rect 4526 362 4529 368
rect 4538 358 4542 361
rect 4478 351 4481 358
rect 4558 352 4561 418
rect 4582 362 4585 468
rect 4598 462 4601 508
rect 4654 482 4657 528
rect 4670 491 4673 568
rect 4666 488 4673 491
rect 4522 348 4526 351
rect 4538 348 4542 351
rect 4466 288 4470 291
rect 4454 272 4457 278
rect 4446 262 4449 268
rect 4398 192 4401 258
rect 4494 242 4497 338
rect 4518 322 4521 348
rect 4558 342 4561 348
rect 4530 338 4534 341
rect 4566 332 4569 338
rect 4518 302 4521 318
rect 4574 302 4577 328
rect 4582 282 4585 358
rect 4590 352 4593 458
rect 4632 403 4634 407
rect 4638 403 4641 407
rect 4645 403 4648 407
rect 4622 352 4625 398
rect 4654 391 4657 478
rect 4710 472 4713 478
rect 4650 388 4657 391
rect 4590 312 4593 348
rect 4422 202 4425 238
rect 4406 192 4409 198
rect 4358 152 4361 158
rect 4366 152 4369 158
rect 4374 152 4377 168
rect 4446 152 4449 218
rect 4382 142 4385 148
rect 4438 142 4441 148
rect 4198 72 4201 78
rect 4230 72 4233 98
rect 4238 92 4241 98
rect 3978 58 3982 61
rect 3966 52 3969 58
rect 4014 52 4017 58
rect 4038 51 4041 58
rect 4094 52 4097 68
rect 4110 52 4113 68
rect 4206 62 4209 68
rect 4222 62 4225 68
rect 4238 62 4241 88
rect 4298 78 4302 81
rect 4342 72 4345 88
rect 4358 72 4361 128
rect 4366 72 4369 98
rect 4318 62 4321 68
rect 4366 62 4369 68
rect 4126 52 4129 59
rect 4382 52 4385 98
rect 4390 82 4393 128
rect 4462 92 4465 218
rect 4502 152 4505 188
rect 4510 152 4513 268
rect 4590 262 4593 298
rect 4606 262 4609 318
rect 4614 312 4617 338
rect 4622 312 4625 348
rect 4650 288 4654 291
rect 4662 272 4665 468
rect 4686 462 4689 468
rect 4718 462 4721 498
rect 4726 492 4729 648
rect 4750 592 4753 638
rect 4758 582 4761 658
rect 4798 652 4801 659
rect 4742 542 4745 548
rect 4782 542 4785 548
rect 4814 542 4817 548
rect 4802 538 4806 541
rect 4754 528 4758 531
rect 4766 492 4769 528
rect 4754 488 4758 491
rect 4738 468 4742 471
rect 4782 462 4785 538
rect 4806 532 4809 538
rect 4814 521 4817 538
rect 4806 518 4817 521
rect 4822 532 4825 628
rect 4862 552 4865 668
rect 4878 552 4881 848
rect 4894 742 4897 868
rect 4894 732 4897 738
rect 4910 732 4913 788
rect 4886 692 4889 698
rect 4910 692 4913 728
rect 4918 712 4921 948
rect 4926 942 4929 948
rect 4934 931 4937 1138
rect 4954 1128 4958 1131
rect 4942 1092 4945 1118
rect 4966 1072 4969 1078
rect 5006 1072 5009 1138
rect 5014 1092 5017 1128
rect 4942 1062 4945 1068
rect 5030 1062 5033 1258
rect 5046 1252 5049 1318
rect 5054 1242 5057 1338
rect 5062 1332 5065 1338
rect 5086 1282 5089 1288
rect 5166 1282 5169 1338
rect 5178 1288 5182 1291
rect 5102 1272 5105 1278
rect 5062 1262 5065 1268
rect 5074 1258 5078 1261
rect 5062 1242 5065 1248
rect 5102 1221 5105 1268
rect 5118 1252 5121 1259
rect 5102 1218 5113 1221
rect 5082 1148 5086 1151
rect 5110 1142 5113 1218
rect 5182 1192 5185 1278
rect 5046 1072 5049 1078
rect 5054 1062 5057 1088
rect 5078 1082 5081 1138
rect 5110 1072 5113 1138
rect 4986 1058 4990 1061
rect 5002 1058 5006 1061
rect 4982 992 4985 1048
rect 5126 1032 5129 1138
rect 5174 1032 5177 1068
rect 4998 962 5001 978
rect 4946 948 4950 951
rect 4926 928 4937 931
rect 4966 932 4969 948
rect 4926 782 4929 928
rect 4934 862 4937 918
rect 4974 892 4977 948
rect 4990 942 4993 948
rect 4982 872 4985 898
rect 4986 868 4990 871
rect 4998 861 5001 958
rect 5030 942 5033 958
rect 5102 951 5105 958
rect 5118 942 5121 1018
rect 5154 948 5158 951
rect 5134 942 5137 948
rect 5034 938 5038 941
rect 5014 932 5017 938
rect 5142 932 5145 948
rect 5162 938 5166 941
rect 5182 932 5185 958
rect 4994 858 5001 861
rect 5006 852 5009 918
rect 5126 892 5129 918
rect 5018 868 5022 871
rect 5078 852 5081 858
rect 4990 842 4993 848
rect 5050 788 5054 791
rect 4926 752 4929 778
rect 4950 742 4953 778
rect 4958 752 4961 758
rect 4898 688 4902 691
rect 4942 662 4945 718
rect 4974 672 4977 738
rect 4998 672 5001 778
rect 5022 752 5025 758
rect 5006 692 5009 748
rect 5038 682 5041 728
rect 5042 668 5046 671
rect 4886 572 4889 648
rect 4910 552 4913 558
rect 4926 552 4929 658
rect 4974 571 4977 668
rect 4990 662 4993 668
rect 4998 662 5001 668
rect 5054 662 5057 768
rect 5062 762 5065 768
rect 5094 752 5097 868
rect 5138 858 5142 861
rect 5118 752 5121 798
rect 5094 742 5097 748
rect 5074 738 5078 741
rect 5018 658 5022 661
rect 5062 652 5065 658
rect 5070 652 5073 718
rect 5082 668 5086 671
rect 4966 568 4977 571
rect 4934 552 4937 568
rect 4966 552 4969 568
rect 4974 552 4977 558
rect 5030 552 5033 588
rect 5082 568 5086 571
rect 4842 548 4846 551
rect 5050 548 5054 551
rect 4862 542 4865 548
rect 4870 542 4873 548
rect 4878 532 4881 548
rect 4894 532 4897 548
rect 5042 538 5046 541
rect 4918 532 4921 538
rect 4798 462 4801 518
rect 4678 352 4681 358
rect 4694 352 4697 418
rect 4662 262 4665 268
rect 4670 262 4673 308
rect 4526 252 4529 259
rect 4518 102 4521 118
rect 4510 92 4513 98
rect 4406 62 4409 78
rect 4462 72 4465 88
rect 4518 72 4521 98
rect 4526 92 4529 208
rect 4542 192 4545 238
rect 4550 92 4553 238
rect 4414 62 4417 68
rect 4542 62 4545 68
rect 4566 62 4569 128
rect 4590 92 4593 248
rect 4632 203 4634 207
rect 4638 203 4641 207
rect 4645 203 4648 207
rect 4670 202 4673 258
rect 4642 168 4646 171
rect 4678 152 4681 348
rect 4686 292 4689 298
rect 4726 292 4729 448
rect 4742 352 4745 358
rect 4774 352 4777 358
rect 4790 352 4793 458
rect 4806 432 4809 518
rect 4822 502 4825 528
rect 4846 492 4849 498
rect 4830 462 4833 468
rect 4854 462 4857 518
rect 4946 488 4950 491
rect 4878 472 4881 478
rect 4998 472 5001 528
rect 5038 482 5041 488
rect 4898 458 4902 461
rect 4814 392 4817 448
rect 4850 388 4854 391
rect 4798 352 4801 368
rect 4862 352 4865 378
rect 4926 372 4929 468
rect 5006 463 5009 468
rect 4942 442 4945 448
rect 4966 352 4969 358
rect 5006 352 5009 358
rect 4810 348 4817 351
rect 4782 342 4785 348
rect 4758 332 4761 338
rect 4750 322 4753 328
rect 4766 322 4769 328
rect 4702 282 4705 288
rect 4722 268 4726 271
rect 4714 258 4718 261
rect 4726 182 4729 268
rect 4734 262 4737 318
rect 4778 268 4782 271
rect 4790 262 4793 338
rect 4798 292 4801 318
rect 4806 282 4809 298
rect 4786 258 4790 261
rect 4774 252 4777 258
rect 4602 148 4606 151
rect 4702 151 4705 158
rect 4734 142 4737 198
rect 4750 192 4753 238
rect 4746 158 4750 161
rect 4746 148 4750 151
rect 4602 138 4606 141
rect 4598 82 4601 108
rect 4574 72 4577 78
rect 4582 62 4585 68
rect 4446 52 4449 59
rect 4034 48 4041 51
rect 4050 48 4054 51
rect 4226 48 4230 51
rect 4554 48 4558 51
rect 3990 42 3993 48
rect 4062 42 4065 48
rect 4238 42 4241 48
rect 4366 42 4369 48
rect 4390 42 4393 48
rect 4406 42 4409 48
rect 3954 38 3958 41
rect 4606 32 4609 138
rect 4622 92 4625 128
rect 4702 72 4705 108
rect 4758 72 4761 208
rect 4774 202 4777 218
rect 4814 192 4817 348
rect 4830 322 4833 348
rect 4870 332 4873 348
rect 4854 252 4857 328
rect 4882 318 4886 321
rect 4894 292 4897 348
rect 5014 342 5017 348
rect 5046 342 5049 538
rect 5062 532 5065 568
rect 5078 542 5081 548
rect 5054 472 5057 528
rect 5094 472 5097 728
rect 5126 712 5129 848
rect 5158 792 5161 868
rect 5166 862 5169 928
rect 5166 772 5169 858
rect 5174 802 5177 858
rect 5182 852 5185 858
rect 5178 788 5182 791
rect 5102 492 5105 708
rect 5142 672 5145 748
rect 5190 722 5193 728
rect 5178 718 5182 721
rect 5146 658 5150 661
rect 5126 552 5129 658
rect 5138 548 5142 551
rect 5126 492 5129 548
rect 5074 468 5078 471
rect 5054 462 5057 468
rect 5062 462 5065 468
rect 5054 352 5057 458
rect 5086 372 5089 458
rect 5062 352 5065 368
rect 5094 342 5097 348
rect 5066 338 5070 341
rect 5110 332 5113 448
rect 5182 422 5185 468
rect 5182 342 5185 418
rect 4910 322 4913 328
rect 4914 288 4918 291
rect 4974 282 4977 328
rect 5022 301 5025 318
rect 5014 298 5025 301
rect 4894 262 4897 268
rect 4942 262 4945 268
rect 4974 263 4977 268
rect 4866 258 4870 261
rect 5014 262 5017 298
rect 5038 292 5041 328
rect 5062 262 5065 298
rect 5078 262 5081 318
rect 5110 292 5113 328
rect 5126 302 5129 318
rect 5098 288 5102 291
rect 5186 288 5190 291
rect 5110 272 5113 278
rect 5042 258 5046 261
rect 4830 222 4833 238
rect 4870 182 4873 248
rect 4906 188 4910 191
rect 4766 162 4769 168
rect 4782 102 4785 148
rect 4790 142 4793 178
rect 4798 122 4801 148
rect 4806 92 4809 118
rect 4814 92 4817 168
rect 4838 152 4841 158
rect 4830 92 4833 148
rect 4846 142 4849 178
rect 4870 172 4873 178
rect 4894 162 4897 168
rect 4942 152 4945 258
rect 4966 152 4969 198
rect 5002 178 5006 181
rect 4854 102 4857 148
rect 4894 132 4897 148
rect 4902 142 4905 148
rect 5022 92 5025 218
rect 5054 152 5057 158
rect 5062 142 5065 258
rect 5110 212 5113 268
rect 5130 258 5134 261
rect 5106 188 5110 191
rect 5166 151 5169 158
rect 5054 92 5057 138
rect 5010 88 5014 91
rect 4838 72 4841 78
rect 4906 68 4910 71
rect 4686 63 4689 68
rect 4950 62 4953 78
rect 4958 72 4961 88
rect 5038 62 5041 78
rect 5122 68 5126 71
rect 5134 62 5137 148
rect 5174 92 5177 108
rect 4754 58 4758 61
rect 4826 58 4830 61
rect 4854 52 4857 58
rect 4818 48 4822 51
rect 536 3 538 7
rect 542 3 545 7
rect 549 3 552 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1573 3 1576 7
rect 2094 -18 2097 18
rect 2584 3 2586 7
rect 2590 3 2593 7
rect 2597 3 2600 7
rect 3254 -18 3257 8
rect 3608 3 3610 7
rect 3614 3 3617 7
rect 3621 3 3624 7
rect 4632 3 4634 7
rect 4638 3 4641 7
rect 4645 3 4648 7
rect 2094 -22 2098 -18
rect 3254 -22 3258 -18
<< m3contact >>
rect 1050 4903 1054 4907
rect 1057 4903 1061 4907
rect 846 4888 850 4892
rect 966 4888 970 4892
rect 1254 4888 1258 4892
rect 230 4878 234 4882
rect 286 4878 290 4882
rect 422 4878 426 4882
rect 454 4878 458 4882
rect 598 4878 602 4882
rect 838 4878 842 4882
rect 870 4878 874 4882
rect 1190 4878 1194 4882
rect 182 4868 186 4872
rect 214 4868 218 4872
rect 246 4868 250 4872
rect 134 4858 138 4862
rect 254 4858 258 4862
rect 190 4848 194 4852
rect 78 4828 82 4832
rect 158 4818 162 4822
rect 246 4838 250 4842
rect 206 4818 210 4822
rect 102 4768 106 4772
rect 134 4758 138 4762
rect 46 4748 50 4752
rect 118 4738 122 4742
rect 158 4748 162 4752
rect 190 4748 194 4752
rect 166 4738 170 4742
rect 182 4738 186 4742
rect 134 4728 138 4732
rect 158 4728 162 4732
rect 110 4718 114 4722
rect 54 4708 58 4712
rect 102 4708 106 4712
rect 174 4708 178 4712
rect 38 4668 42 4672
rect 6 4588 10 4592
rect 46 4588 50 4592
rect 94 4698 98 4702
rect 134 4688 138 4692
rect 182 4688 186 4692
rect 102 4678 106 4682
rect 246 4738 250 4742
rect 270 4818 274 4822
rect 374 4828 378 4832
rect 382 4818 386 4822
rect 342 4808 346 4812
rect 366 4808 370 4812
rect 366 4788 370 4792
rect 310 4758 314 4762
rect 310 4748 314 4752
rect 262 4718 266 4722
rect 310 4718 314 4722
rect 206 4698 210 4702
rect 126 4668 130 4672
rect 190 4668 194 4672
rect 110 4658 114 4662
rect 142 4658 146 4662
rect 102 4648 106 4652
rect 94 4558 98 4562
rect 70 4548 74 4552
rect 14 4538 18 4542
rect 22 4498 26 4502
rect 94 4498 98 4502
rect 102 4478 106 4482
rect 246 4658 250 4662
rect 310 4708 314 4712
rect 310 4688 314 4692
rect 342 4738 346 4742
rect 350 4718 354 4722
rect 326 4688 330 4692
rect 318 4678 322 4682
rect 302 4668 306 4672
rect 254 4648 258 4652
rect 262 4648 266 4652
rect 190 4638 194 4642
rect 262 4628 266 4632
rect 190 4568 194 4572
rect 286 4658 290 4662
rect 278 4578 282 4582
rect 270 4558 274 4562
rect 334 4668 338 4672
rect 318 4568 322 4572
rect 686 4868 690 4872
rect 710 4868 714 4872
rect 742 4868 746 4872
rect 990 4868 994 4872
rect 1070 4868 1074 4872
rect 566 4858 570 4862
rect 582 4858 586 4862
rect 382 4728 386 4732
rect 366 4668 370 4672
rect 702 4858 706 4862
rect 582 4848 586 4852
rect 614 4848 618 4852
rect 638 4848 642 4852
rect 502 4818 506 4822
rect 526 4818 530 4822
rect 538 4803 542 4807
rect 545 4803 549 4807
rect 574 4798 578 4802
rect 614 4758 618 4762
rect 694 4838 698 4842
rect 710 4838 714 4842
rect 678 4798 682 4802
rect 678 4778 682 4782
rect 686 4768 690 4772
rect 726 4778 730 4782
rect 678 4748 682 4752
rect 702 4748 706 4752
rect 470 4728 474 4732
rect 430 4708 434 4712
rect 470 4698 474 4702
rect 526 4728 530 4732
rect 478 4688 482 4692
rect 430 4668 434 4672
rect 446 4668 450 4672
rect 462 4668 466 4672
rect 390 4658 394 4662
rect 422 4658 426 4662
rect 446 4648 450 4652
rect 374 4638 378 4642
rect 382 4578 386 4582
rect 374 4558 378 4562
rect 118 4548 122 4552
rect 166 4548 170 4552
rect 278 4548 282 4552
rect 302 4548 306 4552
rect 310 4548 314 4552
rect 326 4548 330 4552
rect 110 4458 114 4462
rect 126 4458 130 4462
rect 54 4418 58 4422
rect 102 4418 106 4422
rect 54 4368 58 4372
rect 6 4358 10 4362
rect 46 4358 50 4362
rect 30 4348 34 4352
rect 86 4358 90 4362
rect 22 4318 26 4322
rect 70 4268 74 4272
rect 62 4258 66 4262
rect 22 4188 26 4192
rect 214 4468 218 4472
rect 166 4458 170 4462
rect 158 4368 162 4372
rect 150 4358 154 4362
rect 190 4448 194 4452
rect 318 4528 322 4532
rect 334 4528 338 4532
rect 294 4488 298 4492
rect 318 4488 322 4492
rect 254 4458 258 4462
rect 278 4458 282 4462
rect 286 4448 290 4452
rect 262 4438 266 4442
rect 182 4358 186 4362
rect 238 4348 242 4352
rect 142 4318 146 4322
rect 142 4278 146 4282
rect 190 4328 194 4332
rect 166 4268 170 4272
rect 126 4228 130 4232
rect 94 4208 98 4212
rect 94 4198 98 4202
rect 86 4188 90 4192
rect 62 4158 66 4162
rect 430 4568 434 4572
rect 366 4538 370 4542
rect 414 4538 418 4542
rect 422 4538 426 4542
rect 398 4528 402 4532
rect 350 4518 354 4522
rect 382 4488 386 4492
rect 398 4478 402 4482
rect 422 4478 426 4482
rect 326 4468 330 4472
rect 350 4468 354 4472
rect 414 4468 418 4472
rect 502 4658 506 4662
rect 518 4658 522 4662
rect 510 4648 514 4652
rect 550 4718 554 4722
rect 726 4748 730 4752
rect 718 4738 722 4742
rect 566 4708 570 4712
rect 686 4708 690 4712
rect 710 4708 714 4712
rect 558 4698 562 4702
rect 582 4688 586 4692
rect 734 4688 738 4692
rect 542 4668 546 4672
rect 526 4638 530 4642
rect 486 4628 490 4632
rect 518 4628 522 4632
rect 462 4558 466 4562
rect 494 4548 498 4552
rect 502 4538 506 4542
rect 518 4538 522 4542
rect 538 4603 542 4607
rect 545 4603 549 4607
rect 678 4678 682 4682
rect 782 4858 786 4862
rect 814 4858 818 4862
rect 846 4858 850 4862
rect 766 4848 770 4852
rect 782 4798 786 4802
rect 758 4748 762 4752
rect 766 4748 770 4752
rect 774 4738 778 4742
rect 750 4698 754 4702
rect 806 4768 810 4772
rect 798 4758 802 4762
rect 798 4748 802 4752
rect 798 4728 802 4732
rect 798 4708 802 4712
rect 798 4688 802 4692
rect 750 4678 754 4682
rect 806 4678 810 4682
rect 878 4858 882 4862
rect 1046 4858 1050 4862
rect 878 4848 882 4852
rect 894 4848 898 4852
rect 910 4848 914 4852
rect 830 4828 834 4832
rect 862 4828 866 4832
rect 822 4758 826 4762
rect 854 4758 858 4762
rect 822 4738 826 4742
rect 598 4658 602 4662
rect 582 4618 586 4622
rect 654 4618 658 4622
rect 526 4528 530 4532
rect 470 4518 474 4522
rect 438 4458 442 4462
rect 446 4458 450 4462
rect 302 4358 306 4362
rect 374 4358 378 4362
rect 398 4358 402 4362
rect 278 4348 282 4352
rect 254 4338 258 4342
rect 238 4328 242 4332
rect 206 4188 210 4192
rect 262 4278 266 4282
rect 246 4268 250 4272
rect 286 4268 290 4272
rect 286 4248 290 4252
rect 270 4208 274 4212
rect 222 4178 226 4182
rect 214 4168 218 4172
rect 222 4158 226 4162
rect 246 4158 250 4162
rect 302 4158 306 4162
rect 142 4148 146 4152
rect 206 4148 210 4152
rect 38 4068 42 4072
rect 134 4138 138 4142
rect 238 4138 242 4142
rect 102 4088 106 4092
rect 150 4088 154 4092
rect 166 4078 170 4082
rect 118 4068 122 4072
rect 142 4068 146 4072
rect 102 4048 106 4052
rect 102 3968 106 3972
rect 294 4148 298 4152
rect 270 4138 274 4142
rect 286 4128 290 4132
rect 278 4078 282 4082
rect 334 4328 338 4332
rect 398 4338 402 4342
rect 486 4458 490 4462
rect 446 4348 450 4352
rect 470 4358 474 4362
rect 518 4468 522 4472
rect 538 4403 542 4407
rect 545 4403 549 4407
rect 710 4668 714 4672
rect 766 4668 770 4672
rect 774 4668 778 4672
rect 670 4658 674 4662
rect 742 4658 746 4662
rect 662 4608 666 4612
rect 702 4638 706 4642
rect 654 4578 658 4582
rect 638 4568 642 4572
rect 662 4568 666 4572
rect 590 4538 594 4542
rect 646 4528 650 4532
rect 638 4478 642 4482
rect 614 4468 618 4472
rect 590 4448 594 4452
rect 630 4448 634 4452
rect 598 4438 602 4442
rect 614 4438 618 4442
rect 574 4408 578 4412
rect 598 4408 602 4412
rect 566 4388 570 4392
rect 574 4368 578 4372
rect 622 4398 626 4402
rect 582 4348 586 4352
rect 598 4348 602 4352
rect 462 4338 466 4342
rect 614 4338 618 4342
rect 638 4338 642 4342
rect 430 4328 434 4332
rect 414 4318 418 4322
rect 422 4318 426 4322
rect 366 4268 370 4272
rect 366 4258 370 4262
rect 374 4258 378 4262
rect 390 4258 394 4262
rect 326 4238 330 4242
rect 350 4238 354 4242
rect 366 4238 370 4242
rect 326 4218 330 4222
rect 382 4198 386 4202
rect 574 4288 578 4292
rect 606 4288 610 4292
rect 422 4268 426 4272
rect 414 4188 418 4192
rect 438 4248 442 4252
rect 558 4258 562 4262
rect 598 4268 602 4272
rect 454 4228 458 4232
rect 550 4228 554 4232
rect 430 4178 434 4182
rect 318 4158 322 4162
rect 374 4148 378 4152
rect 430 4148 434 4152
rect 390 4138 394 4142
rect 422 4138 426 4142
rect 342 4128 346 4132
rect 342 4118 346 4122
rect 310 4068 314 4072
rect 334 4068 338 4072
rect 246 4058 250 4062
rect 270 4058 274 4062
rect 302 4058 306 4062
rect 190 4048 194 4052
rect 150 3968 154 3972
rect 94 3948 98 3952
rect 110 3948 114 3952
rect 142 3948 146 3952
rect 38 3938 42 3942
rect 38 3918 42 3922
rect 118 3938 122 3942
rect 166 3948 170 3952
rect 246 3958 250 3962
rect 190 3938 194 3942
rect 166 3928 170 3932
rect 174 3928 178 3932
rect 94 3898 98 3902
rect 206 3898 210 3902
rect 110 3888 114 3892
rect 198 3888 202 3892
rect 278 4038 282 4042
rect 326 4048 330 4052
rect 318 4028 322 4032
rect 310 4008 314 4012
rect 374 4118 378 4122
rect 494 4178 498 4182
rect 470 4158 474 4162
rect 538 4203 542 4207
rect 545 4203 549 4207
rect 510 4158 514 4162
rect 566 4158 570 4162
rect 478 4138 482 4142
rect 462 4108 466 4112
rect 510 4118 514 4122
rect 478 4088 482 4092
rect 486 4088 490 4092
rect 494 4088 498 4092
rect 422 4078 426 4082
rect 382 4068 386 4072
rect 334 3938 338 3942
rect 310 3918 314 3922
rect 334 3918 338 3922
rect 270 3888 274 3892
rect 182 3878 186 3882
rect 262 3878 266 3882
rect 230 3858 234 3862
rect 246 3858 250 3862
rect 262 3858 266 3862
rect 278 3858 282 3862
rect 166 3848 170 3852
rect 206 3838 210 3842
rect 222 3838 226 3842
rect 342 3898 346 3902
rect 326 3858 330 3862
rect 318 3848 322 3852
rect 302 3818 306 3822
rect 334 3818 338 3822
rect 246 3798 250 3802
rect 134 3778 138 3782
rect 454 4068 458 4072
rect 454 4058 458 4062
rect 462 4058 466 4062
rect 438 4038 442 4042
rect 374 4008 378 4012
rect 382 3978 386 3982
rect 406 3988 410 3992
rect 526 4148 530 4152
rect 582 4148 586 4152
rect 526 4118 530 4122
rect 590 4088 594 4092
rect 494 4078 498 4082
rect 686 4558 690 4562
rect 678 4548 682 4552
rect 678 4528 682 4532
rect 678 4468 682 4472
rect 846 4708 850 4712
rect 854 4678 858 4682
rect 798 4658 802 4662
rect 814 4658 818 4662
rect 838 4658 842 4662
rect 758 4598 762 4602
rect 766 4578 770 4582
rect 718 4568 722 4572
rect 726 4568 730 4572
rect 790 4568 794 4572
rect 702 4548 706 4552
rect 750 4538 754 4542
rect 734 4528 738 4532
rect 750 4528 754 4532
rect 750 4518 754 4522
rect 758 4518 762 4522
rect 702 4478 706 4482
rect 702 4458 706 4462
rect 718 4458 722 4462
rect 774 4548 778 4552
rect 790 4548 794 4552
rect 846 4648 850 4652
rect 854 4638 858 4642
rect 910 4768 914 4772
rect 1014 4758 1018 4762
rect 886 4688 890 4692
rect 870 4648 874 4652
rect 862 4628 866 4632
rect 822 4618 826 4622
rect 902 4618 906 4622
rect 806 4578 810 4582
rect 806 4538 810 4542
rect 790 4528 794 4532
rect 766 4498 770 4502
rect 798 4488 802 4492
rect 758 4478 762 4482
rect 782 4478 786 4482
rect 734 4458 738 4462
rect 694 4438 698 4442
rect 694 4398 698 4402
rect 694 4348 698 4352
rect 662 4298 666 4302
rect 694 4288 698 4292
rect 654 4268 658 4272
rect 734 4378 738 4382
rect 758 4398 762 4402
rect 742 4328 746 4332
rect 726 4278 730 4282
rect 710 4248 714 4252
rect 750 4308 754 4312
rect 734 4258 738 4262
rect 814 4518 818 4522
rect 806 4468 810 4472
rect 814 4438 818 4442
rect 806 4428 810 4432
rect 766 4358 770 4362
rect 798 4378 802 4382
rect 806 4348 810 4352
rect 774 4338 778 4342
rect 766 4288 770 4292
rect 838 4568 842 4572
rect 1254 4868 1258 4872
rect 1150 4858 1154 4862
rect 1230 4858 1234 4862
rect 1238 4838 1242 4842
rect 1070 4818 1074 4822
rect 1286 4868 1290 4872
rect 2074 4903 2078 4907
rect 2081 4903 2085 4907
rect 3098 4903 3102 4907
rect 3105 4903 3109 4907
rect 2270 4888 2274 4892
rect 2310 4888 2314 4892
rect 2398 4888 2402 4892
rect 1502 4878 1506 4882
rect 1774 4878 1778 4882
rect 1806 4878 1810 4882
rect 1838 4878 1842 4882
rect 1958 4878 1962 4882
rect 1974 4878 1978 4882
rect 2174 4878 2178 4882
rect 2382 4878 2386 4882
rect 1550 4868 1554 4872
rect 1598 4868 1602 4872
rect 1686 4868 1690 4872
rect 1758 4868 1762 4872
rect 1790 4868 1794 4872
rect 1334 4858 1338 4862
rect 1358 4859 1362 4863
rect 1478 4859 1482 4863
rect 1270 4838 1274 4842
rect 1246 4828 1250 4832
rect 1174 4758 1178 4762
rect 1182 4758 1186 4762
rect 1150 4738 1154 4742
rect 1086 4728 1090 4732
rect 1126 4728 1130 4732
rect 1070 4708 1074 4712
rect 1050 4703 1054 4707
rect 1057 4703 1061 4707
rect 966 4688 970 4692
rect 1126 4698 1130 4702
rect 1166 4688 1170 4692
rect 1190 4748 1194 4752
rect 1294 4848 1298 4852
rect 1294 4828 1298 4832
rect 1310 4828 1314 4832
rect 1326 4808 1330 4812
rect 1286 4748 1290 4752
rect 1318 4748 1322 4752
rect 1182 4738 1186 4742
rect 1206 4728 1210 4732
rect 1190 4718 1194 4722
rect 1270 4738 1274 4742
rect 1286 4738 1290 4742
rect 1262 4708 1266 4712
rect 1278 4698 1282 4702
rect 1238 4688 1242 4692
rect 1246 4688 1250 4692
rect 1158 4678 1162 4682
rect 1182 4678 1186 4682
rect 934 4668 938 4672
rect 1006 4668 1010 4672
rect 1134 4668 1138 4672
rect 1158 4668 1162 4672
rect 1190 4668 1194 4672
rect 1014 4658 1018 4662
rect 990 4638 994 4642
rect 950 4568 954 4572
rect 902 4558 906 4562
rect 918 4558 922 4562
rect 958 4558 962 4562
rect 1022 4628 1026 4632
rect 846 4548 850 4552
rect 966 4548 970 4552
rect 990 4548 994 4552
rect 838 4538 842 4542
rect 894 4538 898 4542
rect 862 4528 866 4532
rect 942 4498 946 4502
rect 878 4478 882 4482
rect 894 4478 898 4482
rect 862 4448 866 4452
rect 886 4428 890 4432
rect 878 4418 882 4422
rect 838 4388 842 4392
rect 870 4388 874 4392
rect 822 4358 826 4362
rect 838 4338 842 4342
rect 870 4328 874 4332
rect 854 4318 858 4322
rect 934 4468 938 4472
rect 982 4528 986 4532
rect 902 4448 906 4452
rect 982 4508 986 4512
rect 990 4508 994 4512
rect 1022 4468 1026 4472
rect 934 4448 938 4452
rect 974 4448 978 4452
rect 998 4448 1002 4452
rect 982 4438 986 4442
rect 1014 4418 1018 4422
rect 1086 4658 1090 4662
rect 1206 4658 1210 4662
rect 1222 4658 1226 4662
rect 1134 4648 1138 4652
rect 1142 4648 1146 4652
rect 1254 4668 1258 4672
rect 1254 4658 1258 4662
rect 1230 4638 1234 4642
rect 1246 4618 1250 4622
rect 1142 4608 1146 4612
rect 1182 4608 1186 4612
rect 1198 4608 1202 4612
rect 1050 4503 1054 4507
rect 1057 4503 1061 4507
rect 1038 4398 1042 4402
rect 1038 4388 1042 4392
rect 958 4368 962 4372
rect 1022 4368 1026 4372
rect 990 4358 994 4362
rect 998 4358 1002 4362
rect 990 4348 994 4352
rect 1014 4348 1018 4352
rect 958 4328 962 4332
rect 998 4338 1002 4342
rect 990 4328 994 4332
rect 918 4318 922 4322
rect 966 4318 970 4322
rect 846 4278 850 4282
rect 894 4278 898 4282
rect 902 4278 906 4282
rect 830 4268 834 4272
rect 782 4258 786 4262
rect 798 4258 802 4262
rect 814 4258 818 4262
rect 878 4258 882 4262
rect 782 4248 786 4252
rect 774 4238 778 4242
rect 734 4208 738 4212
rect 758 4198 762 4202
rect 854 4248 858 4252
rect 870 4248 874 4252
rect 822 4228 826 4232
rect 806 4188 810 4192
rect 742 4168 746 4172
rect 766 4168 770 4172
rect 718 4158 722 4162
rect 678 4148 682 4152
rect 638 4138 642 4142
rect 630 4088 634 4092
rect 486 4068 490 4072
rect 542 4068 546 4072
rect 582 4068 586 4072
rect 614 4068 618 4072
rect 518 4058 522 4062
rect 494 4048 498 4052
rect 526 4048 530 4052
rect 470 4038 474 4042
rect 574 4038 578 4042
rect 538 4003 542 4007
rect 545 4003 549 4007
rect 366 3958 370 3962
rect 398 3958 402 3962
rect 454 3958 458 3962
rect 542 3958 546 3962
rect 366 3948 370 3952
rect 406 3948 410 3952
rect 446 3948 450 3952
rect 694 4098 698 4102
rect 750 4138 754 4142
rect 838 4158 842 4162
rect 902 4268 906 4272
rect 966 4278 970 4282
rect 998 4318 1002 4322
rect 934 4268 938 4272
rect 950 4268 954 4272
rect 958 4268 962 4272
rect 998 4268 1002 4272
rect 918 4258 922 4262
rect 910 4198 914 4202
rect 934 4238 938 4242
rect 990 4238 994 4242
rect 942 4208 946 4212
rect 926 4188 930 4192
rect 790 4148 794 4152
rect 822 4148 826 4152
rect 846 4148 850 4152
rect 926 4148 930 4152
rect 830 4128 834 4132
rect 886 4128 890 4132
rect 918 4128 922 4132
rect 662 4088 666 4092
rect 710 4078 714 4082
rect 670 4068 674 4072
rect 686 4068 690 4072
rect 646 4048 650 4052
rect 734 4048 738 4052
rect 774 4088 778 4092
rect 798 4068 802 4072
rect 718 4038 722 4042
rect 742 4038 746 4042
rect 750 4038 754 4042
rect 638 4018 642 4022
rect 598 3958 602 3962
rect 678 3958 682 3962
rect 758 4028 762 4032
rect 742 3988 746 3992
rect 462 3948 466 3952
rect 590 3948 594 3952
rect 614 3948 618 3952
rect 862 4088 866 4092
rect 878 4088 882 4092
rect 854 4068 858 4072
rect 862 4068 866 4072
rect 902 4068 906 4072
rect 918 4068 922 4072
rect 918 4048 922 4052
rect 950 4168 954 4172
rect 1014 4248 1018 4252
rect 950 4158 954 4162
rect 982 4158 986 4162
rect 1126 4518 1130 4522
rect 1102 4478 1106 4482
rect 1094 4458 1098 4462
rect 1086 4398 1090 4402
rect 1102 4348 1106 4352
rect 1126 4388 1130 4392
rect 1158 4558 1162 4562
rect 1222 4578 1226 4582
rect 1198 4568 1202 4572
rect 1214 4568 1218 4572
rect 1246 4568 1250 4572
rect 1238 4548 1242 4552
rect 1190 4508 1194 4512
rect 1158 4488 1162 4492
rect 1174 4468 1178 4472
rect 1190 4458 1194 4462
rect 1198 4448 1202 4452
rect 1166 4428 1170 4432
rect 1206 4398 1210 4402
rect 1190 4388 1194 4392
rect 1174 4358 1178 4362
rect 1166 4338 1170 4342
rect 1142 4328 1146 4332
rect 1158 4328 1162 4332
rect 1238 4528 1242 4532
rect 1230 4518 1234 4522
rect 1222 4468 1226 4472
rect 1238 4478 1242 4482
rect 1230 4448 1234 4452
rect 1270 4448 1274 4452
rect 1214 4388 1218 4392
rect 1222 4358 1226 4362
rect 1230 4348 1234 4352
rect 1214 4338 1218 4342
rect 1262 4338 1266 4342
rect 1110 4318 1114 4322
rect 1182 4318 1186 4322
rect 1094 4308 1098 4312
rect 1050 4303 1054 4307
rect 1057 4303 1061 4307
rect 1054 4268 1058 4272
rect 1038 4258 1042 4262
rect 1102 4259 1106 4263
rect 1166 4288 1170 4292
rect 1190 4278 1194 4282
rect 1174 4268 1178 4272
rect 1150 4258 1154 4262
rect 1030 4248 1034 4252
rect 1054 4248 1058 4252
rect 1166 4248 1170 4252
rect 1190 4248 1194 4252
rect 1150 4238 1154 4242
rect 1174 4188 1178 4192
rect 1206 4248 1210 4252
rect 1206 4238 1210 4242
rect 1046 4168 1050 4172
rect 1182 4168 1186 4172
rect 1110 4158 1114 4162
rect 982 4148 986 4152
rect 1174 4148 1178 4152
rect 990 4138 994 4142
rect 1014 4138 1018 4142
rect 1166 4138 1170 4142
rect 950 4128 954 4132
rect 950 4108 954 4112
rect 886 4038 890 4042
rect 942 4038 946 4042
rect 822 3988 826 3992
rect 846 3988 850 3992
rect 790 3948 794 3952
rect 374 3938 378 3942
rect 414 3938 418 3942
rect 422 3938 426 3942
rect 590 3938 594 3942
rect 734 3938 738 3942
rect 398 3928 402 3932
rect 366 3878 370 3882
rect 374 3868 378 3872
rect 406 3878 410 3882
rect 406 3848 410 3852
rect 390 3828 394 3832
rect 366 3818 370 3822
rect 374 3808 378 3812
rect 310 3758 314 3762
rect 350 3758 354 3762
rect 206 3738 210 3742
rect 6 3688 10 3692
rect 94 3678 98 3682
rect 174 3678 178 3682
rect 54 3668 58 3672
rect 30 3658 34 3662
rect 46 3658 50 3662
rect 6 3598 10 3602
rect 158 3668 162 3672
rect 222 3668 226 3672
rect 150 3648 154 3652
rect 118 3628 122 3632
rect 6 3448 10 3452
rect 110 3488 114 3492
rect 70 3468 74 3472
rect 150 3548 154 3552
rect 190 3648 194 3652
rect 166 3628 170 3632
rect 190 3608 194 3612
rect 198 3558 202 3562
rect 182 3548 186 3552
rect 158 3538 162 3542
rect 166 3528 170 3532
rect 198 3528 202 3532
rect 174 3518 178 3522
rect 126 3498 130 3502
rect 166 3478 170 3482
rect 150 3468 154 3472
rect 190 3478 194 3482
rect 110 3458 114 3462
rect 102 3438 106 3442
rect 134 3448 138 3452
rect 150 3428 154 3432
rect 158 3428 162 3432
rect 118 3418 122 3422
rect 94 3338 98 3342
rect 118 3338 122 3342
rect 14 3298 18 3302
rect 6 3258 10 3262
rect 78 3308 82 3312
rect 78 3298 82 3302
rect 62 3268 66 3272
rect 230 3658 234 3662
rect 270 3718 274 3722
rect 294 3718 298 3722
rect 302 3708 306 3712
rect 438 3918 442 3922
rect 566 3928 570 3932
rect 670 3928 674 3932
rect 478 3918 482 3922
rect 470 3908 474 3912
rect 742 3918 746 3922
rect 662 3898 666 3902
rect 494 3868 498 3872
rect 566 3868 570 3872
rect 486 3858 490 3862
rect 422 3818 426 3822
rect 462 3818 466 3822
rect 478 3818 482 3822
rect 430 3798 434 3802
rect 406 3788 410 3792
rect 414 3788 418 3792
rect 422 3758 426 3762
rect 414 3748 418 3752
rect 350 3738 354 3742
rect 382 3738 386 3742
rect 310 3678 314 3682
rect 254 3658 258 3662
rect 222 3498 226 3502
rect 222 3478 226 3482
rect 238 3478 242 3482
rect 246 3478 250 3482
rect 214 3468 218 3472
rect 230 3468 234 3472
rect 206 3438 210 3442
rect 246 3438 250 3442
rect 214 3428 218 3432
rect 230 3378 234 3382
rect 238 3368 242 3372
rect 174 3358 178 3362
rect 230 3348 234 3352
rect 166 3328 170 3332
rect 230 3328 234 3332
rect 238 3328 242 3332
rect 126 3298 130 3302
rect 118 3288 122 3292
rect 134 3278 138 3282
rect 222 3298 226 3302
rect 182 3288 186 3292
rect 110 3258 114 3262
rect 118 3258 122 3262
rect 166 3258 170 3262
rect 70 3248 74 3252
rect 86 3248 90 3252
rect 110 3248 114 3252
rect 62 3168 66 3172
rect 70 3158 74 3162
rect 110 3168 114 3172
rect 22 3138 26 3142
rect 54 3138 58 3142
rect 6 3078 10 3082
rect 14 2978 18 2982
rect 14 2948 18 2952
rect 14 2928 18 2932
rect 102 3138 106 3142
rect 94 3128 98 3132
rect 118 3138 122 3142
rect 118 3128 122 3132
rect 126 3078 130 3082
rect 158 3078 162 3082
rect 174 3078 178 3082
rect 86 3058 90 3062
rect 118 3058 122 3062
rect 174 3058 178 3062
rect 62 3038 66 3042
rect 70 2958 74 2962
rect 102 2978 106 2982
rect 150 2978 154 2982
rect 54 2918 58 2922
rect 70 2898 74 2902
rect 14 2888 18 2892
rect 214 3278 218 3282
rect 198 3158 202 3162
rect 214 3108 218 3112
rect 206 3068 210 3072
rect 206 3038 210 3042
rect 126 2948 130 2952
rect 182 2948 186 2952
rect 198 2948 202 2952
rect 150 2938 154 2942
rect 118 2918 122 2922
rect 142 2918 146 2922
rect 190 2898 194 2902
rect 134 2888 138 2892
rect 158 2888 162 2892
rect 182 2888 186 2892
rect 86 2878 90 2882
rect 102 2868 106 2872
rect 158 2878 162 2882
rect 6 2748 10 2752
rect 70 2738 74 2742
rect 38 2668 42 2672
rect 142 2838 146 2842
rect 134 2738 138 2742
rect 126 2698 130 2702
rect 158 2748 162 2752
rect 182 2738 186 2742
rect 182 2688 186 2692
rect 118 2668 122 2672
rect 150 2668 154 2672
rect 190 2678 194 2682
rect 398 3728 402 3732
rect 350 3718 354 3722
rect 334 3698 338 3702
rect 358 3698 362 3702
rect 366 3698 370 3702
rect 374 3688 378 3692
rect 406 3688 410 3692
rect 318 3658 322 3662
rect 358 3658 362 3662
rect 278 3648 282 3652
rect 278 3598 282 3602
rect 318 3578 322 3582
rect 294 3568 298 3572
rect 262 3558 266 3562
rect 302 3558 306 3562
rect 326 3558 330 3562
rect 286 3548 290 3552
rect 270 3528 274 3532
rect 278 3518 282 3522
rect 278 3478 282 3482
rect 302 3468 306 3472
rect 262 3458 266 3462
rect 262 3438 266 3442
rect 326 3478 330 3482
rect 278 3428 282 3432
rect 318 3428 322 3432
rect 262 3378 266 3382
rect 254 3298 258 3302
rect 254 3288 258 3292
rect 326 3358 330 3362
rect 262 3278 266 3282
rect 302 3338 306 3342
rect 286 3318 290 3322
rect 286 3288 290 3292
rect 318 3298 322 3302
rect 430 3748 434 3752
rect 446 3728 450 3732
rect 446 3668 450 3672
rect 454 3648 458 3652
rect 538 3803 542 3807
rect 545 3803 549 3807
rect 510 3698 514 3702
rect 542 3698 546 3702
rect 486 3668 490 3672
rect 470 3658 474 3662
rect 398 3638 402 3642
rect 438 3638 442 3642
rect 390 3628 394 3632
rect 374 3608 378 3612
rect 358 3558 362 3562
rect 358 3538 362 3542
rect 382 3568 386 3572
rect 454 3628 458 3632
rect 414 3618 418 3622
rect 486 3588 490 3592
rect 454 3578 458 3582
rect 446 3568 450 3572
rect 406 3558 410 3562
rect 430 3558 434 3562
rect 742 3898 746 3902
rect 726 3868 730 3872
rect 774 3868 778 3872
rect 846 3978 850 3982
rect 838 3958 842 3962
rect 870 3968 874 3972
rect 854 3958 858 3962
rect 870 3948 874 3952
rect 854 3938 858 3942
rect 838 3908 842 3912
rect 838 3878 842 3882
rect 878 3868 882 3872
rect 606 3858 610 3862
rect 718 3858 722 3862
rect 782 3858 786 3862
rect 870 3858 874 3862
rect 822 3848 826 3852
rect 702 3828 706 3832
rect 686 3818 690 3822
rect 742 3788 746 3792
rect 654 3768 658 3772
rect 590 3758 594 3762
rect 766 3778 770 3782
rect 750 3758 754 3762
rect 710 3748 714 3752
rect 686 3738 690 3742
rect 630 3698 634 3702
rect 574 3668 578 3672
rect 566 3658 570 3662
rect 606 3658 610 3662
rect 526 3638 530 3642
rect 538 3603 542 3607
rect 545 3603 549 3607
rect 646 3668 650 3672
rect 598 3588 602 3592
rect 510 3568 514 3572
rect 582 3548 586 3552
rect 398 3538 402 3542
rect 366 3518 370 3522
rect 390 3468 394 3472
rect 382 3458 386 3462
rect 398 3458 402 3462
rect 342 3288 346 3292
rect 286 3268 290 3272
rect 294 3268 298 3272
rect 326 3268 330 3272
rect 238 3258 242 3262
rect 254 3258 258 3262
rect 246 3238 250 3242
rect 270 3228 274 3232
rect 278 3228 282 3232
rect 230 3188 234 3192
rect 278 3168 282 3172
rect 310 3238 314 3242
rect 286 3098 290 3102
rect 270 3078 274 3082
rect 238 3068 242 3072
rect 286 3068 290 3072
rect 310 3068 314 3072
rect 294 3058 298 3062
rect 278 2958 282 2962
rect 222 2938 226 2942
rect 230 2938 234 2942
rect 214 2908 218 2912
rect 222 2848 226 2852
rect 214 2698 218 2702
rect 206 2668 210 2672
rect 126 2658 130 2662
rect 142 2658 146 2662
rect 158 2648 162 2652
rect 190 2648 194 2652
rect 190 2598 194 2602
rect 62 2568 66 2572
rect 166 2568 170 2572
rect 126 2558 130 2562
rect 46 2548 50 2552
rect 102 2548 106 2552
rect 222 2678 226 2682
rect 238 2928 242 2932
rect 246 2908 250 2912
rect 238 2898 242 2902
rect 350 3258 354 3262
rect 358 3248 362 3252
rect 422 3518 426 3522
rect 414 3478 418 3482
rect 478 3538 482 3542
rect 494 3538 498 3542
rect 526 3528 530 3532
rect 454 3508 458 3512
rect 470 3498 474 3502
rect 454 3468 458 3472
rect 462 3468 466 3472
rect 582 3538 586 3542
rect 566 3518 570 3522
rect 542 3508 546 3512
rect 622 3558 626 3562
rect 614 3548 618 3552
rect 614 3528 618 3532
rect 438 3458 442 3462
rect 534 3458 538 3462
rect 406 3448 410 3452
rect 422 3438 426 3442
rect 406 3388 410 3392
rect 390 3368 394 3372
rect 406 3368 410 3372
rect 398 3348 402 3352
rect 422 3358 426 3362
rect 446 3358 450 3362
rect 510 3368 514 3372
rect 566 3448 570 3452
rect 574 3438 578 3442
rect 558 3408 562 3412
rect 538 3403 542 3407
rect 545 3403 549 3407
rect 542 3368 546 3372
rect 510 3358 514 3362
rect 526 3358 530 3362
rect 526 3348 530 3352
rect 646 3648 650 3652
rect 670 3728 674 3732
rect 670 3708 674 3712
rect 718 3718 722 3722
rect 726 3698 730 3702
rect 894 3978 898 3982
rect 942 3968 946 3972
rect 942 3938 946 3942
rect 950 3938 954 3942
rect 918 3908 922 3912
rect 966 4068 970 4072
rect 1006 4068 1010 4072
rect 1014 4058 1018 4062
rect 974 4038 978 4042
rect 982 3988 986 3992
rect 958 3908 962 3912
rect 902 3878 906 3882
rect 926 3868 930 3872
rect 966 3868 970 3872
rect 926 3838 930 3842
rect 974 3838 978 3842
rect 918 3828 922 3832
rect 886 3798 890 3802
rect 910 3798 914 3802
rect 894 3788 898 3792
rect 806 3778 810 3782
rect 774 3768 778 3772
rect 902 3768 906 3772
rect 814 3758 818 3762
rect 774 3728 778 3732
rect 798 3738 802 3742
rect 790 3698 794 3702
rect 822 3698 826 3702
rect 782 3688 786 3692
rect 934 3808 938 3812
rect 934 3798 938 3802
rect 950 3778 954 3782
rect 950 3758 954 3762
rect 966 3758 970 3762
rect 1006 4048 1010 4052
rect 998 4008 1002 4012
rect 1022 4008 1026 4012
rect 1022 3968 1026 3972
rect 1050 4103 1054 4107
rect 1057 4103 1061 4107
rect 1142 4088 1146 4092
rect 1062 4068 1066 4072
rect 1126 4068 1130 4072
rect 1158 4068 1162 4072
rect 1158 4058 1162 4062
rect 1054 3988 1058 3992
rect 1102 3968 1106 3972
rect 1182 4088 1186 4092
rect 1166 4018 1170 4022
rect 1150 3978 1154 3982
rect 1174 3978 1178 3982
rect 1142 3968 1146 3972
rect 998 3928 1002 3932
rect 998 3868 1002 3872
rect 1006 3858 1010 3862
rect 1046 3948 1050 3952
rect 1110 3948 1114 3952
rect 1062 3938 1066 3942
rect 1050 3903 1054 3907
rect 1057 3903 1061 3907
rect 1030 3868 1034 3872
rect 1062 3868 1066 3872
rect 1022 3858 1026 3862
rect 998 3848 1002 3852
rect 1014 3848 1018 3852
rect 1054 3848 1058 3852
rect 1062 3848 1066 3852
rect 1030 3828 1034 3832
rect 1022 3768 1026 3772
rect 1006 3758 1010 3762
rect 982 3748 986 3752
rect 990 3748 994 3752
rect 894 3738 898 3742
rect 942 3738 946 3742
rect 974 3738 978 3742
rect 862 3718 866 3722
rect 990 3718 994 3722
rect 838 3688 842 3692
rect 814 3678 818 3682
rect 854 3678 858 3682
rect 934 3678 938 3682
rect 678 3668 682 3672
rect 758 3668 762 3672
rect 910 3668 914 3672
rect 950 3668 954 3672
rect 974 3678 978 3682
rect 718 3658 722 3662
rect 766 3658 770 3662
rect 886 3658 890 3662
rect 958 3658 962 3662
rect 974 3658 978 3662
rect 686 3638 690 3642
rect 654 3628 658 3632
rect 646 3588 650 3592
rect 654 3568 658 3572
rect 638 3528 642 3532
rect 686 3548 690 3552
rect 646 3508 650 3512
rect 646 3488 650 3492
rect 638 3478 642 3482
rect 670 3458 674 3462
rect 598 3448 602 3452
rect 614 3448 618 3452
rect 678 3448 682 3452
rect 726 3578 730 3582
rect 798 3578 802 3582
rect 654 3438 658 3442
rect 686 3438 690 3442
rect 654 3418 658 3422
rect 598 3348 602 3352
rect 526 3338 530 3342
rect 574 3338 578 3342
rect 494 3328 498 3332
rect 582 3318 586 3322
rect 398 3308 402 3312
rect 390 3298 394 3302
rect 382 3278 386 3282
rect 374 3238 378 3242
rect 374 3228 378 3232
rect 326 3208 330 3212
rect 342 3198 346 3202
rect 350 3188 354 3192
rect 342 3178 346 3182
rect 326 3158 330 3162
rect 422 3298 426 3302
rect 414 3288 418 3292
rect 350 3148 354 3152
rect 606 3298 610 3302
rect 494 3288 498 3292
rect 598 3288 602 3292
rect 598 3278 602 3282
rect 526 3258 530 3262
rect 582 3238 586 3242
rect 526 3228 530 3232
rect 454 3208 458 3212
rect 478 3208 482 3212
rect 454 3178 458 3182
rect 470 3158 474 3162
rect 538 3203 542 3207
rect 545 3203 549 3207
rect 566 3168 570 3172
rect 422 3148 426 3152
rect 494 3148 498 3152
rect 526 3148 530 3152
rect 406 3138 410 3142
rect 486 3138 490 3142
rect 382 3128 386 3132
rect 390 3128 394 3132
rect 358 3118 362 3122
rect 390 3118 394 3122
rect 406 3108 410 3112
rect 470 3128 474 3132
rect 414 3098 418 3102
rect 422 3098 426 3102
rect 390 3078 394 3082
rect 342 3058 346 3062
rect 326 3038 330 3042
rect 462 3078 466 3082
rect 422 3068 426 3072
rect 414 3058 418 3062
rect 374 3048 378 3052
rect 406 3048 410 3052
rect 358 3028 362 3032
rect 390 3018 394 3022
rect 342 2988 346 2992
rect 358 2988 362 2992
rect 318 2918 322 2922
rect 342 2968 346 2972
rect 430 3028 434 3032
rect 430 2978 434 2982
rect 406 2968 410 2972
rect 374 2958 378 2962
rect 390 2958 394 2962
rect 358 2948 362 2952
rect 366 2938 370 2942
rect 342 2898 346 2902
rect 326 2888 330 2892
rect 478 3118 482 3122
rect 470 2958 474 2962
rect 422 2938 426 2942
rect 526 3108 530 3112
rect 518 3088 522 3092
rect 502 3078 506 3082
rect 486 3068 490 3072
rect 486 2968 490 2972
rect 494 2968 498 2972
rect 518 2968 522 2972
rect 582 3128 586 3132
rect 734 3558 738 3562
rect 806 3548 810 3552
rect 838 3548 842 3552
rect 878 3648 882 3652
rect 926 3648 930 3652
rect 942 3648 946 3652
rect 990 3648 994 3652
rect 870 3628 874 3632
rect 894 3628 898 3632
rect 846 3538 850 3542
rect 798 3528 802 3532
rect 790 3508 794 3512
rect 742 3448 746 3452
rect 734 3428 738 3432
rect 694 3378 698 3382
rect 710 3378 714 3382
rect 662 3358 666 3362
rect 646 3348 650 3352
rect 686 3348 690 3352
rect 646 3338 650 3342
rect 630 3298 634 3302
rect 622 3288 626 3292
rect 614 3268 618 3272
rect 678 3328 682 3332
rect 710 3328 714 3332
rect 654 3308 658 3312
rect 686 3308 690 3312
rect 686 3288 690 3292
rect 726 3398 730 3402
rect 742 3378 746 3382
rect 902 3618 906 3622
rect 878 3568 882 3572
rect 918 3568 922 3572
rect 1094 3938 1098 3942
rect 1102 3928 1106 3932
rect 1078 3908 1082 3912
rect 1118 3908 1122 3912
rect 1102 3888 1106 3892
rect 1118 3888 1122 3892
rect 1198 4168 1202 4172
rect 1222 4328 1226 4332
rect 1230 4318 1234 4322
rect 1246 4308 1250 4312
rect 1262 4278 1266 4282
rect 1222 4258 1226 4262
rect 1246 4258 1250 4262
rect 1222 4248 1226 4252
rect 1230 4208 1234 4212
rect 1222 4188 1226 4192
rect 1222 4158 1226 4162
rect 1214 4148 1218 4152
rect 1222 4128 1226 4132
rect 1190 4058 1194 4062
rect 1158 3968 1162 3972
rect 1166 3968 1170 3972
rect 1182 3968 1186 3972
rect 1150 3898 1154 3902
rect 1142 3888 1146 3892
rect 1174 3928 1178 3932
rect 1158 3878 1162 3882
rect 1166 3878 1170 3882
rect 1358 4758 1362 4762
rect 1414 4808 1418 4812
rect 1350 4748 1354 4752
rect 1374 4748 1378 4752
rect 1398 4738 1402 4742
rect 1318 4718 1322 4722
rect 1302 4698 1306 4702
rect 1302 4678 1306 4682
rect 1334 4678 1338 4682
rect 1302 4658 1306 4662
rect 1318 4658 1322 4662
rect 1286 4558 1290 4562
rect 1294 4538 1298 4542
rect 1286 4358 1290 4362
rect 1374 4668 1378 4672
rect 1382 4658 1386 4662
rect 1534 4858 1538 4862
rect 1502 4768 1506 4772
rect 1422 4758 1426 4762
rect 1502 4748 1506 4752
rect 1454 4698 1458 4702
rect 1430 4678 1434 4682
rect 1470 4678 1474 4682
rect 1454 4658 1458 4662
rect 1446 4648 1450 4652
rect 1422 4638 1426 4642
rect 1430 4638 1434 4642
rect 1446 4638 1450 4642
rect 1414 4578 1418 4582
rect 1342 4548 1346 4552
rect 1358 4548 1362 4552
rect 1374 4548 1378 4552
rect 1454 4548 1458 4552
rect 1502 4658 1506 4662
rect 1526 4788 1530 4792
rect 1622 4828 1626 4832
rect 1654 4808 1658 4812
rect 1562 4803 1566 4807
rect 1569 4803 1573 4807
rect 1542 4778 1546 4782
rect 1566 4778 1570 4782
rect 1518 4768 1522 4772
rect 1558 4768 1562 4772
rect 1574 4758 1578 4762
rect 1606 4758 1610 4762
rect 1518 4728 1522 4732
rect 1510 4618 1514 4622
rect 1502 4548 1506 4552
rect 1366 4538 1370 4542
rect 1398 4538 1402 4542
rect 1446 4538 1450 4542
rect 1342 4508 1346 4512
rect 1310 4498 1314 4502
rect 1342 4478 1346 4482
rect 1398 4508 1402 4512
rect 1358 4468 1362 4472
rect 1438 4498 1442 4502
rect 1422 4478 1426 4482
rect 1510 4478 1514 4482
rect 1494 4468 1498 4472
rect 1502 4458 1506 4462
rect 1430 4448 1434 4452
rect 1494 4448 1498 4452
rect 1414 4438 1418 4442
rect 1478 4438 1482 4442
rect 1294 4338 1298 4342
rect 1334 4408 1338 4412
rect 1366 4388 1370 4392
rect 1334 4358 1338 4362
rect 1366 4348 1370 4352
rect 1310 4268 1314 4272
rect 1326 4268 1330 4272
rect 1286 4258 1290 4262
rect 1318 4258 1322 4262
rect 1246 4128 1250 4132
rect 1310 4248 1314 4252
rect 1326 4208 1330 4212
rect 1390 4338 1394 4342
rect 1342 4328 1346 4332
rect 1374 4298 1378 4302
rect 1342 4288 1346 4292
rect 1358 4268 1362 4272
rect 1470 4378 1474 4382
rect 1486 4368 1490 4372
rect 1478 4358 1482 4362
rect 1470 4348 1474 4352
rect 1454 4318 1458 4322
rect 1406 4288 1410 4292
rect 1430 4288 1434 4292
rect 1382 4248 1386 4252
rect 1382 4238 1386 4242
rect 1334 4178 1338 4182
rect 1510 4388 1514 4392
rect 1486 4338 1490 4342
rect 1470 4298 1474 4302
rect 1438 4258 1442 4262
rect 1502 4258 1506 4262
rect 1558 4628 1562 4632
rect 1598 4748 1602 4752
rect 1630 4748 1634 4752
rect 1678 4858 1682 4862
rect 1670 4808 1674 4812
rect 1702 4838 1706 4842
rect 1734 4838 1738 4842
rect 1790 4838 1794 4842
rect 1694 4808 1698 4812
rect 1710 4828 1714 4832
rect 1678 4748 1682 4752
rect 1606 4738 1610 4742
rect 1622 4738 1626 4742
rect 1638 4738 1642 4742
rect 1694 4738 1698 4742
rect 1702 4738 1706 4742
rect 1598 4718 1602 4722
rect 1662 4728 1666 4732
rect 1638 4698 1642 4702
rect 1574 4678 1578 4682
rect 1646 4678 1650 4682
rect 1590 4658 1594 4662
rect 1582 4648 1586 4652
rect 1622 4648 1626 4652
rect 1606 4638 1610 4642
rect 1558 4618 1562 4622
rect 1566 4618 1570 4622
rect 1582 4618 1586 4622
rect 1562 4603 1566 4607
rect 1569 4603 1573 4607
rect 1550 4588 1554 4592
rect 1622 4628 1626 4632
rect 1590 4588 1594 4592
rect 1630 4588 1634 4592
rect 1598 4548 1602 4552
rect 1638 4548 1642 4552
rect 1598 4528 1602 4532
rect 1614 4528 1618 4532
rect 1550 4508 1554 4512
rect 1614 4518 1618 4522
rect 1558 4468 1562 4472
rect 1590 4468 1594 4472
rect 1622 4478 1626 4482
rect 1622 4448 1626 4452
rect 1566 4428 1570 4432
rect 1582 4418 1586 4422
rect 1562 4403 1566 4407
rect 1569 4403 1573 4407
rect 1598 4338 1602 4342
rect 1534 4328 1538 4332
rect 1574 4308 1578 4312
rect 1582 4288 1586 4292
rect 1310 4148 1314 4152
rect 1262 4118 1266 4122
rect 1294 4118 1298 4122
rect 1358 4138 1362 4142
rect 1326 4128 1330 4132
rect 1342 4128 1346 4132
rect 1358 4128 1362 4132
rect 1302 4108 1306 4112
rect 1310 4108 1314 4112
rect 1286 4098 1290 4102
rect 1222 4088 1226 4092
rect 1230 4088 1234 4092
rect 1262 4068 1266 4072
rect 1246 4058 1250 4062
rect 1230 4008 1234 4012
rect 1198 3988 1202 3992
rect 1238 3988 1242 3992
rect 1230 3978 1234 3982
rect 1198 3968 1202 3972
rect 1214 3968 1218 3972
rect 1198 3958 1202 3962
rect 1206 3958 1210 3962
rect 1190 3948 1194 3952
rect 1294 4038 1298 4042
rect 1310 4038 1314 4042
rect 1254 4028 1258 4032
rect 1294 4018 1298 4022
rect 1278 3998 1282 4002
rect 1254 3978 1258 3982
rect 1190 3888 1194 3892
rect 1198 3878 1202 3882
rect 1142 3868 1146 3872
rect 1094 3858 1098 3862
rect 1110 3858 1114 3862
rect 1070 3838 1074 3842
rect 1014 3718 1018 3722
rect 1006 3688 1010 3692
rect 1070 3738 1074 3742
rect 1030 3698 1034 3702
rect 1022 3688 1026 3692
rect 1070 3708 1074 3712
rect 1050 3703 1054 3707
rect 1057 3703 1061 3707
rect 1094 3808 1098 3812
rect 1102 3768 1106 3772
rect 1158 3848 1162 3852
rect 1150 3838 1154 3842
rect 1142 3798 1146 3802
rect 1118 3758 1122 3762
rect 1134 3758 1138 3762
rect 1206 3848 1210 3852
rect 1174 3838 1178 3842
rect 1166 3808 1170 3812
rect 1214 3808 1218 3812
rect 1150 3748 1154 3752
rect 1142 3728 1146 3732
rect 1110 3718 1114 3722
rect 1126 3718 1130 3722
rect 1118 3698 1122 3702
rect 1102 3678 1106 3682
rect 1038 3668 1042 3672
rect 1078 3668 1082 3672
rect 1094 3668 1098 3672
rect 1174 3738 1178 3742
rect 1278 3938 1282 3942
rect 1262 3928 1266 3932
rect 1238 3918 1242 3922
rect 1238 3888 1242 3892
rect 1262 3888 1266 3892
rect 1302 3948 1306 3952
rect 1318 3948 1322 3952
rect 1318 3908 1322 3912
rect 1310 3898 1314 3902
rect 1398 4138 1402 4142
rect 1382 4118 1386 4122
rect 1398 4118 1402 4122
rect 1382 4088 1386 4092
rect 1366 4068 1370 4072
rect 1422 4108 1426 4112
rect 1406 4078 1410 4082
rect 1454 4158 1458 4162
rect 1494 4158 1498 4162
rect 1454 4148 1458 4152
rect 1462 4098 1466 4102
rect 1414 4068 1418 4072
rect 1430 4068 1434 4072
rect 1406 4058 1410 4062
rect 1510 4128 1514 4132
rect 1510 4118 1514 4122
rect 1550 4248 1554 4252
rect 1654 4508 1658 4512
rect 1646 4488 1650 4492
rect 1646 4458 1650 4462
rect 1638 4448 1642 4452
rect 1630 4348 1634 4352
rect 1638 4348 1642 4352
rect 1646 4338 1650 4342
rect 1630 4328 1634 4332
rect 1646 4298 1650 4302
rect 1614 4278 1618 4282
rect 1590 4268 1594 4272
rect 1614 4248 1618 4252
rect 1574 4218 1578 4222
rect 1582 4218 1586 4222
rect 1562 4203 1566 4207
rect 1569 4203 1573 4207
rect 1526 4168 1530 4172
rect 1526 4148 1530 4152
rect 1518 4078 1522 4082
rect 1518 4068 1522 4072
rect 1494 4058 1498 4062
rect 1382 4038 1386 4042
rect 1350 3908 1354 3912
rect 1342 3898 1346 3902
rect 1334 3878 1338 3882
rect 1302 3868 1306 3872
rect 1390 3938 1394 3942
rect 1390 3928 1394 3932
rect 1366 3898 1370 3902
rect 1374 3888 1378 3892
rect 1398 3898 1402 3902
rect 1366 3868 1370 3872
rect 1358 3858 1362 3862
rect 1326 3848 1330 3852
rect 1358 3848 1362 3852
rect 1350 3838 1354 3842
rect 1334 3828 1338 3832
rect 1302 3778 1306 3782
rect 1326 3768 1330 3772
rect 1302 3758 1306 3762
rect 1302 3748 1306 3752
rect 1310 3738 1314 3742
rect 1230 3728 1234 3732
rect 1166 3678 1170 3682
rect 1014 3658 1018 3662
rect 1038 3658 1042 3662
rect 1118 3658 1122 3662
rect 1126 3658 1130 3662
rect 1014 3648 1018 3652
rect 1086 3648 1090 3652
rect 1150 3648 1154 3652
rect 1182 3648 1186 3652
rect 998 3638 1002 3642
rect 934 3628 938 3632
rect 1006 3588 1010 3592
rect 918 3558 922 3562
rect 886 3548 890 3552
rect 902 3548 906 3552
rect 822 3528 826 3532
rect 870 3528 874 3532
rect 854 3508 858 3512
rect 862 3508 866 3512
rect 846 3488 850 3492
rect 846 3458 850 3462
rect 862 3458 866 3462
rect 830 3448 834 3452
rect 838 3448 842 3452
rect 806 3368 810 3372
rect 782 3358 786 3362
rect 798 3348 802 3352
rect 726 3338 730 3342
rect 726 3298 730 3302
rect 750 3338 754 3342
rect 718 3288 722 3292
rect 654 3278 658 3282
rect 670 3258 674 3262
rect 702 3258 706 3262
rect 630 3248 634 3252
rect 662 3248 666 3252
rect 702 3228 706 3232
rect 670 3218 674 3222
rect 646 3168 650 3172
rect 638 3148 642 3152
rect 598 3118 602 3122
rect 574 3108 578 3112
rect 614 3108 618 3112
rect 550 3098 554 3102
rect 542 3088 546 3092
rect 538 3003 542 3007
rect 545 3003 549 3007
rect 606 3078 610 3082
rect 630 3078 634 3082
rect 558 2988 562 2992
rect 566 2978 570 2982
rect 606 3038 610 3042
rect 558 2958 562 2962
rect 574 2958 578 2962
rect 486 2948 490 2952
rect 462 2928 466 2932
rect 414 2918 418 2922
rect 278 2868 282 2872
rect 366 2868 370 2872
rect 398 2868 402 2872
rect 254 2848 258 2852
rect 350 2838 354 2842
rect 374 2838 378 2842
rect 430 2848 434 2852
rect 414 2788 418 2792
rect 246 2768 250 2772
rect 262 2768 266 2772
rect 366 2768 370 2772
rect 246 2738 250 2742
rect 278 2748 282 2752
rect 302 2747 306 2751
rect 382 2748 386 2752
rect 398 2748 402 2752
rect 430 2748 434 2752
rect 326 2738 330 2742
rect 310 2718 314 2722
rect 262 2668 266 2672
rect 238 2658 242 2662
rect 270 2658 274 2662
rect 294 2658 298 2662
rect 230 2648 234 2652
rect 254 2588 258 2592
rect 318 2588 322 2592
rect 294 2578 298 2582
rect 294 2568 298 2572
rect 206 2548 210 2552
rect 270 2548 274 2552
rect 142 2538 146 2542
rect 110 2528 114 2532
rect 102 2518 106 2522
rect 150 2518 154 2522
rect 134 2508 138 2512
rect 150 2498 154 2502
rect 22 2488 26 2492
rect 142 2488 146 2492
rect 14 2468 18 2472
rect 182 2468 186 2472
rect 110 2459 114 2463
rect 134 2458 138 2462
rect 30 2448 34 2452
rect 6 2378 10 2382
rect 14 2288 18 2292
rect 350 2718 354 2722
rect 374 2688 378 2692
rect 462 2858 466 2862
rect 446 2698 450 2702
rect 470 2688 474 2692
rect 334 2668 338 2672
rect 350 2668 354 2672
rect 366 2668 370 2672
rect 406 2668 410 2672
rect 318 2538 322 2542
rect 246 2508 250 2512
rect 246 2488 250 2492
rect 438 2618 442 2622
rect 342 2598 346 2602
rect 390 2578 394 2582
rect 430 2578 434 2582
rect 382 2558 386 2562
rect 510 2948 514 2952
rect 526 2928 530 2932
rect 566 2938 570 2942
rect 654 3068 658 3072
rect 686 3148 690 3152
rect 686 3118 690 3122
rect 838 3388 842 3392
rect 910 3518 914 3522
rect 878 3378 882 3382
rect 870 3368 874 3372
rect 878 3358 882 3362
rect 894 3348 898 3352
rect 862 3328 866 3332
rect 902 3288 906 3292
rect 870 3278 874 3282
rect 734 3268 738 3272
rect 774 3268 778 3272
rect 854 3268 858 3272
rect 878 3268 882 3272
rect 742 3258 746 3262
rect 854 3258 858 3262
rect 734 3238 738 3242
rect 798 3188 802 3192
rect 774 3158 778 3162
rect 934 3548 938 3552
rect 926 3478 930 3482
rect 942 3518 946 3522
rect 982 3538 986 3542
rect 990 3538 994 3542
rect 974 3518 978 3522
rect 950 3498 954 3502
rect 990 3508 994 3512
rect 942 3488 946 3492
rect 982 3488 986 3492
rect 958 3458 962 3462
rect 998 3458 1002 3462
rect 966 3398 970 3402
rect 982 3398 986 3402
rect 958 3378 962 3382
rect 982 3368 986 3372
rect 926 3348 930 3352
rect 918 3328 922 3332
rect 934 3298 938 3302
rect 950 3288 954 3292
rect 998 3358 1002 3362
rect 982 3328 986 3332
rect 982 3318 986 3322
rect 974 3298 978 3302
rect 926 3268 930 3272
rect 958 3268 962 3272
rect 966 3268 970 3272
rect 982 3268 986 3272
rect 886 3258 890 3262
rect 886 3248 890 3252
rect 862 3168 866 3172
rect 814 3158 818 3162
rect 838 3158 842 3162
rect 854 3158 858 3162
rect 702 3138 706 3142
rect 742 3138 746 3142
rect 766 3138 770 3142
rect 806 3138 810 3142
rect 710 3118 714 3122
rect 702 3088 706 3092
rect 678 3078 682 3082
rect 838 3128 842 3132
rect 782 3118 786 3122
rect 726 3088 730 3092
rect 734 3078 738 3082
rect 694 3048 698 3052
rect 622 3038 626 3042
rect 614 3018 618 3022
rect 662 2958 666 2962
rect 670 2958 674 2962
rect 686 2958 690 2962
rect 582 2908 586 2912
rect 574 2898 578 2902
rect 654 2938 658 2942
rect 678 2938 682 2942
rect 734 2938 738 2942
rect 638 2898 642 2902
rect 646 2888 650 2892
rect 526 2868 530 2872
rect 598 2868 602 2872
rect 494 2858 498 2862
rect 494 2848 498 2852
rect 494 2758 498 2762
rect 510 2748 514 2752
rect 502 2718 506 2722
rect 478 2658 482 2662
rect 494 2648 498 2652
rect 486 2568 490 2572
rect 494 2568 498 2572
rect 510 2668 514 2672
rect 542 2858 546 2862
rect 590 2858 594 2862
rect 558 2848 562 2852
rect 538 2803 542 2807
rect 545 2803 549 2807
rect 678 2928 682 2932
rect 670 2888 674 2892
rect 702 2888 706 2892
rect 702 2868 706 2872
rect 606 2798 610 2802
rect 646 2798 650 2802
rect 710 2848 714 2852
rect 694 2838 698 2842
rect 694 2828 698 2832
rect 662 2778 666 2782
rect 582 2768 586 2772
rect 550 2758 554 2762
rect 566 2748 570 2752
rect 638 2748 642 2752
rect 654 2748 658 2752
rect 574 2718 578 2722
rect 582 2708 586 2712
rect 574 2688 578 2692
rect 526 2648 530 2652
rect 558 2648 562 2652
rect 534 2628 538 2632
rect 538 2603 542 2607
rect 545 2603 549 2607
rect 534 2568 538 2572
rect 398 2538 402 2542
rect 478 2538 482 2542
rect 486 2538 490 2542
rect 510 2538 514 2542
rect 382 2518 386 2522
rect 414 2518 418 2522
rect 422 2508 426 2512
rect 270 2488 274 2492
rect 334 2488 338 2492
rect 374 2478 378 2482
rect 310 2468 314 2472
rect 262 2458 266 2462
rect 230 2448 234 2452
rect 302 2448 306 2452
rect 214 2428 218 2432
rect 126 2388 130 2392
rect 206 2388 210 2392
rect 94 2358 98 2362
rect 166 2368 170 2372
rect 158 2358 162 2362
rect 182 2358 186 2362
rect 214 2358 218 2362
rect 158 2348 162 2352
rect 70 2278 74 2282
rect 118 2278 122 2282
rect 110 2268 114 2272
rect 134 2308 138 2312
rect 134 2288 138 2292
rect 110 2258 114 2262
rect 126 2258 130 2262
rect 270 2368 274 2372
rect 342 2418 346 2422
rect 318 2368 322 2372
rect 326 2358 330 2362
rect 358 2368 362 2372
rect 382 2468 386 2472
rect 470 2528 474 2532
rect 494 2528 498 2532
rect 454 2508 458 2512
rect 446 2488 450 2492
rect 502 2488 506 2492
rect 574 2638 578 2642
rect 606 2618 610 2622
rect 622 2588 626 2592
rect 582 2568 586 2572
rect 574 2558 578 2562
rect 590 2548 594 2552
rect 718 2828 722 2832
rect 646 2738 650 2742
rect 702 2698 706 2702
rect 710 2688 714 2692
rect 686 2668 690 2672
rect 646 2648 650 2652
rect 646 2548 650 2552
rect 558 2538 562 2542
rect 566 2508 570 2512
rect 638 2528 642 2532
rect 614 2518 618 2522
rect 534 2478 538 2482
rect 542 2478 546 2482
rect 590 2478 594 2482
rect 398 2448 402 2452
rect 502 2438 506 2442
rect 478 2388 482 2392
rect 382 2368 386 2372
rect 430 2368 434 2372
rect 478 2368 482 2372
rect 494 2368 498 2372
rect 350 2348 354 2352
rect 366 2348 370 2352
rect 302 2318 306 2322
rect 294 2288 298 2292
rect 326 2288 330 2292
rect 294 2268 298 2272
rect 302 2268 306 2272
rect 150 2188 154 2192
rect 110 2158 114 2162
rect 6 2148 10 2152
rect 14 2088 18 2092
rect 86 2147 90 2151
rect 118 2118 122 2122
rect 166 2258 170 2262
rect 270 2258 274 2262
rect 230 2248 234 2252
rect 198 2228 202 2232
rect 158 2178 162 2182
rect 166 2148 170 2152
rect 182 2138 186 2142
rect 166 2098 170 2102
rect 158 2088 162 2092
rect 70 2078 74 2082
rect 118 2068 122 2072
rect 134 2068 138 2072
rect 190 2078 194 2082
rect 174 2068 178 2072
rect 102 2048 106 2052
rect 182 2048 186 2052
rect 158 2038 162 2042
rect 222 2168 226 2172
rect 246 2168 250 2172
rect 230 2158 234 2162
rect 246 2148 250 2152
rect 214 2108 218 2112
rect 230 2108 234 2112
rect 246 2108 250 2112
rect 222 2088 226 2092
rect 238 2088 242 2092
rect 230 2078 234 2082
rect 206 2048 210 2052
rect 86 2008 90 2012
rect 134 2008 138 2012
rect 182 1978 186 1982
rect 118 1948 122 1952
rect 14 1938 18 1942
rect 70 1938 74 1942
rect 6 1878 10 1882
rect 6 1828 10 1832
rect 198 1938 202 1942
rect 158 1898 162 1902
rect 134 1878 138 1882
rect 102 1858 106 1862
rect 70 1848 74 1852
rect 110 1848 114 1852
rect 174 1888 178 1892
rect 166 1868 170 1872
rect 158 1858 162 1862
rect 142 1848 146 1852
rect 126 1838 130 1842
rect 166 1798 170 1802
rect 86 1748 90 1752
rect 62 1738 66 1742
rect 190 1858 194 1862
rect 238 1958 242 1962
rect 302 2238 306 2242
rect 294 2208 298 2212
rect 278 2178 282 2182
rect 358 2298 362 2302
rect 350 2278 354 2282
rect 342 2268 346 2272
rect 486 2338 490 2342
rect 502 2338 506 2342
rect 406 2318 410 2322
rect 382 2298 386 2302
rect 390 2298 394 2302
rect 534 2458 538 2462
rect 538 2403 542 2407
rect 545 2403 549 2407
rect 590 2458 594 2462
rect 606 2458 610 2462
rect 574 2448 578 2452
rect 606 2448 610 2452
rect 598 2398 602 2402
rect 542 2378 546 2382
rect 558 2378 562 2382
rect 566 2378 570 2382
rect 526 2368 530 2372
rect 526 2338 530 2342
rect 510 2308 514 2312
rect 446 2298 450 2302
rect 470 2298 474 2302
rect 502 2298 506 2302
rect 454 2288 458 2292
rect 478 2288 482 2292
rect 470 2268 474 2272
rect 510 2268 514 2272
rect 350 2258 354 2262
rect 366 2258 370 2262
rect 366 2188 370 2192
rect 574 2368 578 2372
rect 550 2298 554 2302
rect 486 2228 490 2232
rect 542 2228 546 2232
rect 538 2203 542 2207
rect 545 2203 549 2207
rect 422 2188 426 2192
rect 406 2148 410 2152
rect 310 2138 314 2142
rect 334 2138 338 2142
rect 270 2038 274 2042
rect 262 2008 266 2012
rect 254 1988 258 1992
rect 294 2128 298 2132
rect 366 2128 370 2132
rect 294 2118 298 2122
rect 278 1978 282 1982
rect 278 1958 282 1962
rect 326 2078 330 2082
rect 462 2178 466 2182
rect 478 2168 482 2172
rect 510 2158 514 2162
rect 502 2148 506 2152
rect 494 2138 498 2142
rect 478 2108 482 2112
rect 486 2108 490 2112
rect 486 2078 490 2082
rect 438 2068 442 2072
rect 422 2058 426 2062
rect 366 2048 370 2052
rect 342 2008 346 2012
rect 302 1978 306 1982
rect 246 1948 250 1952
rect 254 1938 258 1942
rect 246 1928 250 1932
rect 222 1918 226 1922
rect 422 1948 426 1952
rect 294 1918 298 1922
rect 342 1928 346 1932
rect 310 1918 314 1922
rect 302 1898 306 1902
rect 222 1868 226 1872
rect 238 1868 242 1872
rect 206 1808 210 1812
rect 270 1848 274 1852
rect 262 1818 266 1822
rect 262 1758 266 1762
rect 214 1748 218 1752
rect 158 1738 162 1742
rect 182 1738 186 1742
rect 222 1738 226 1742
rect 126 1718 130 1722
rect 78 1698 82 1702
rect 182 1728 186 1732
rect 166 1708 170 1712
rect 158 1678 162 1682
rect 94 1668 98 1672
rect 110 1668 114 1672
rect 214 1728 218 1732
rect 190 1688 194 1692
rect 102 1568 106 1572
rect 46 1548 50 1552
rect 278 1818 282 1822
rect 270 1698 274 1702
rect 262 1678 266 1682
rect 270 1658 274 1662
rect 254 1628 258 1632
rect 150 1568 154 1572
rect 126 1548 130 1552
rect 102 1538 106 1542
rect 62 1528 66 1532
rect 94 1478 98 1482
rect 166 1528 170 1532
rect 110 1508 114 1512
rect 134 1508 138 1512
rect 134 1488 138 1492
rect 46 1458 50 1462
rect 126 1458 130 1462
rect 174 1508 178 1512
rect 166 1478 170 1482
rect 190 1488 194 1492
rect 182 1468 186 1472
rect 110 1438 114 1442
rect 102 1378 106 1382
rect 102 1368 106 1372
rect 54 1348 58 1352
rect 102 1338 106 1342
rect 62 1318 66 1322
rect 102 1288 106 1292
rect 126 1388 130 1392
rect 134 1378 138 1382
rect 134 1358 138 1362
rect 150 1358 154 1362
rect 118 1338 122 1342
rect 134 1288 138 1292
rect 102 1258 106 1262
rect 38 1248 42 1252
rect 110 1238 114 1242
rect 110 1158 114 1162
rect 14 1138 18 1142
rect 62 1128 66 1132
rect 86 1128 90 1132
rect 38 1078 42 1082
rect 46 1058 50 1062
rect 102 1068 106 1072
rect 110 1068 114 1072
rect 94 1048 98 1052
rect 174 1458 178 1462
rect 246 1618 250 1622
rect 382 1898 386 1902
rect 374 1888 378 1892
rect 390 1878 394 1882
rect 414 1908 418 1912
rect 406 1888 410 1892
rect 422 1888 426 1892
rect 374 1868 378 1872
rect 398 1868 402 1872
rect 406 1858 410 1862
rect 422 1838 426 1842
rect 326 1818 330 1822
rect 318 1788 322 1792
rect 358 1778 362 1782
rect 342 1758 346 1762
rect 382 1748 386 1752
rect 374 1738 378 1742
rect 358 1718 362 1722
rect 326 1698 330 1702
rect 374 1678 378 1682
rect 446 2058 450 2062
rect 438 2048 442 2052
rect 462 2048 466 2052
rect 470 2038 474 2042
rect 454 2028 458 2032
rect 470 1958 474 1962
rect 446 1948 450 1952
rect 438 1928 442 1932
rect 446 1918 450 1922
rect 446 1868 450 1872
rect 590 2288 594 2292
rect 582 2278 586 2282
rect 606 2358 610 2362
rect 622 2498 626 2502
rect 630 2488 634 2492
rect 646 2508 650 2512
rect 718 2678 722 2682
rect 774 3098 778 3102
rect 758 3088 762 3092
rect 750 2978 754 2982
rect 798 3088 802 3092
rect 838 3108 842 3112
rect 846 3088 850 3092
rect 878 3148 882 3152
rect 902 3188 906 3192
rect 902 3178 906 3182
rect 1006 3258 1010 3262
rect 966 3248 970 3252
rect 1038 3618 1042 3622
rect 1022 3578 1026 3582
rect 1134 3598 1138 3602
rect 1142 3568 1146 3572
rect 1182 3568 1186 3572
rect 1070 3558 1074 3562
rect 1134 3558 1138 3562
rect 1054 3548 1058 3552
rect 1038 3538 1042 3542
rect 1050 3503 1054 3507
rect 1057 3503 1061 3507
rect 1046 3488 1050 3492
rect 1166 3548 1170 3552
rect 1126 3528 1130 3532
rect 1126 3518 1130 3522
rect 1094 3508 1098 3512
rect 1118 3508 1122 3512
rect 1046 3458 1050 3462
rect 1062 3458 1066 3462
rect 1030 3438 1034 3442
rect 1022 3378 1026 3382
rect 1022 3358 1026 3362
rect 1110 3438 1114 3442
rect 1086 3368 1090 3372
rect 1102 3358 1106 3362
rect 1070 3348 1074 3352
rect 1102 3348 1106 3352
rect 1070 3338 1074 3342
rect 1110 3338 1114 3342
rect 1050 3303 1054 3307
rect 1057 3303 1061 3307
rect 1070 3298 1074 3302
rect 1190 3498 1194 3502
rect 1134 3438 1138 3442
rect 1126 3358 1130 3362
rect 1142 3408 1146 3412
rect 1174 3398 1178 3402
rect 1150 3358 1154 3362
rect 1158 3358 1162 3362
rect 1126 3338 1130 3342
rect 1166 3338 1170 3342
rect 1118 3288 1122 3292
rect 1134 3288 1138 3292
rect 1174 3288 1178 3292
rect 1078 3268 1082 3272
rect 990 3228 994 3232
rect 1014 3228 1018 3232
rect 990 3208 994 3212
rect 1094 3248 1098 3252
rect 1126 3248 1130 3252
rect 1142 3248 1146 3252
rect 1054 3178 1058 3182
rect 918 3158 922 3162
rect 950 3138 954 3142
rect 894 3128 898 3132
rect 878 3118 882 3122
rect 958 3118 962 3122
rect 862 3078 866 3082
rect 870 3068 874 3072
rect 886 3098 890 3102
rect 886 3088 890 3092
rect 894 3078 898 3082
rect 838 3058 842 3062
rect 822 3048 826 3052
rect 830 3038 834 3042
rect 942 3078 946 3082
rect 934 3068 938 3072
rect 894 3028 898 3032
rect 942 3038 946 3042
rect 934 3028 938 3032
rect 958 3028 962 3032
rect 806 2978 810 2982
rect 918 2978 922 2982
rect 910 2968 914 2972
rect 782 2958 786 2962
rect 782 2948 786 2952
rect 822 2948 826 2952
rect 838 2948 842 2952
rect 878 2948 882 2952
rect 950 2948 954 2952
rect 798 2938 802 2942
rect 806 2938 810 2942
rect 782 2928 786 2932
rect 774 2908 778 2912
rect 758 2868 762 2872
rect 926 2938 930 2942
rect 1046 3158 1050 3162
rect 1110 3198 1114 3202
rect 1102 3188 1106 3192
rect 998 3148 1002 3152
rect 1078 3138 1082 3142
rect 1014 3128 1018 3132
rect 982 3118 986 3122
rect 982 3088 986 3092
rect 1030 3108 1034 3112
rect 1050 3103 1054 3107
rect 1057 3103 1061 3107
rect 1118 3178 1122 3182
rect 1134 3178 1138 3182
rect 1182 3278 1186 3282
rect 1294 3718 1298 3722
rect 1278 3708 1282 3712
rect 1326 3708 1330 3712
rect 1262 3668 1266 3672
rect 1206 3658 1210 3662
rect 1222 3658 1226 3662
rect 1254 3628 1258 3632
rect 1214 3618 1218 3622
rect 1302 3688 1306 3692
rect 1278 3608 1282 3612
rect 1246 3598 1250 3602
rect 1286 3598 1290 3602
rect 1238 3588 1242 3592
rect 1278 3588 1282 3592
rect 1230 3428 1234 3432
rect 1206 3328 1210 3332
rect 1230 3328 1234 3332
rect 1246 3548 1250 3552
rect 1318 3648 1322 3652
rect 1350 3798 1354 3802
rect 1358 3768 1362 3772
rect 1342 3738 1346 3742
rect 1366 3738 1370 3742
rect 1350 3698 1354 3702
rect 1366 3678 1370 3682
rect 1406 3848 1410 3852
rect 1422 3988 1426 3992
rect 1470 4028 1474 4032
rect 1454 3978 1458 3982
rect 1446 3968 1450 3972
rect 1494 3948 1498 3952
rect 1494 3938 1498 3942
rect 1494 3918 1498 3922
rect 1430 3898 1434 3902
rect 1470 3898 1474 3902
rect 1462 3888 1466 3892
rect 1446 3878 1450 3882
rect 1438 3868 1442 3872
rect 1478 3868 1482 3872
rect 1486 3858 1490 3862
rect 1750 4808 1754 4812
rect 1726 4768 1730 4772
rect 1822 4868 1826 4872
rect 1886 4818 1890 4822
rect 1814 4788 1818 4792
rect 1734 4738 1738 4742
rect 1710 4678 1714 4682
rect 1710 4658 1714 4662
rect 1694 4608 1698 4612
rect 1670 4588 1674 4592
rect 1710 4538 1714 4542
rect 1806 4738 1810 4742
rect 1790 4728 1794 4732
rect 1726 4718 1730 4722
rect 1774 4668 1778 4672
rect 1950 4778 1954 4782
rect 1950 4768 1954 4772
rect 1846 4748 1850 4752
rect 1886 4748 1890 4752
rect 1870 4738 1874 4742
rect 1878 4738 1882 4742
rect 1854 4718 1858 4722
rect 1862 4708 1866 4712
rect 1814 4698 1818 4702
rect 1782 4658 1786 4662
rect 1806 4658 1810 4662
rect 1798 4648 1802 4652
rect 1814 4638 1818 4642
rect 1774 4628 1778 4632
rect 1766 4618 1770 4622
rect 1798 4618 1802 4622
rect 1790 4588 1794 4592
rect 1798 4558 1802 4562
rect 1782 4538 1786 4542
rect 1718 4528 1722 4532
rect 1750 4518 1754 4522
rect 1766 4508 1770 4512
rect 1758 4488 1762 4492
rect 1678 4468 1682 4472
rect 1694 4448 1698 4452
rect 1686 4418 1690 4422
rect 1710 4418 1714 4422
rect 1670 4348 1674 4352
rect 1638 4238 1642 4242
rect 1614 4208 1618 4212
rect 1630 4198 1634 4202
rect 1630 4148 1634 4152
rect 1550 4058 1554 4062
rect 1606 4138 1610 4142
rect 1566 4118 1570 4122
rect 1606 4108 1610 4112
rect 1662 4228 1666 4232
rect 1654 4148 1658 4152
rect 1734 4418 1738 4422
rect 1750 4358 1754 4362
rect 1694 4328 1698 4332
rect 1686 4308 1690 4312
rect 1694 4298 1698 4302
rect 1686 4288 1690 4292
rect 1702 4268 1706 4272
rect 1838 4638 1842 4642
rect 1822 4608 1826 4612
rect 1814 4548 1818 4552
rect 1830 4548 1834 4552
rect 1774 4458 1778 4462
rect 1790 4458 1794 4462
rect 1782 4448 1786 4452
rect 1902 4718 1906 4722
rect 1886 4708 1890 4712
rect 1942 4688 1946 4692
rect 1910 4678 1914 4682
rect 2094 4868 2098 4872
rect 2134 4868 2138 4872
rect 2006 4858 2010 4862
rect 2062 4838 2066 4842
rect 2054 4818 2058 4822
rect 2038 4758 2042 4762
rect 2118 4858 2122 4862
rect 2118 4838 2122 4842
rect 2086 4818 2090 4822
rect 2078 4808 2082 4812
rect 2086 4778 2090 4782
rect 2118 4778 2122 4782
rect 1998 4748 2002 4752
rect 2046 4748 2050 4752
rect 2102 4758 2106 4762
rect 2054 4738 2058 4742
rect 2014 4728 2018 4732
rect 2022 4728 2026 4732
rect 2030 4718 2034 4722
rect 1998 4708 2002 4712
rect 2022 4708 2026 4712
rect 1974 4698 1978 4702
rect 1894 4668 1898 4672
rect 1958 4668 1962 4672
rect 1950 4658 1954 4662
rect 1926 4648 1930 4652
rect 1950 4648 1954 4652
rect 1942 4638 1946 4642
rect 1974 4638 1978 4642
rect 1918 4628 1922 4632
rect 1982 4628 1986 4632
rect 1886 4558 1890 4562
rect 1950 4578 1954 4582
rect 1926 4568 1930 4572
rect 1974 4568 1978 4572
rect 2038 4668 2042 4672
rect 1998 4658 2002 4662
rect 2014 4628 2018 4632
rect 2038 4598 2042 4602
rect 1918 4528 1922 4532
rect 1926 4528 1930 4532
rect 1902 4508 1906 4512
rect 1878 4478 1882 4482
rect 2254 4868 2258 4872
rect 2302 4868 2306 4872
rect 2190 4858 2194 4862
rect 2246 4858 2250 4862
rect 2174 4768 2178 4772
rect 2182 4768 2186 4772
rect 2150 4748 2154 4752
rect 2254 4828 2258 4832
rect 2230 4788 2234 4792
rect 2206 4768 2210 4772
rect 2198 4758 2202 4762
rect 2230 4758 2234 4762
rect 2246 4748 2250 4752
rect 2166 4728 2170 4732
rect 2102 4718 2106 4722
rect 2134 4718 2138 4722
rect 2074 4703 2078 4707
rect 2081 4703 2085 4707
rect 2270 4838 2274 4842
rect 2270 4778 2274 4782
rect 2262 4738 2266 4742
rect 2230 4728 2234 4732
rect 2174 4708 2178 4712
rect 2214 4698 2218 4702
rect 2062 4688 2066 4692
rect 2134 4678 2138 4682
rect 2158 4678 2162 4682
rect 2054 4668 2058 4672
rect 2078 4658 2082 4662
rect 2118 4648 2122 4652
rect 2238 4688 2242 4692
rect 2238 4668 2242 4672
rect 2214 4638 2218 4642
rect 2102 4608 2106 4612
rect 2158 4588 2162 4592
rect 2086 4558 2090 4562
rect 2142 4558 2146 4562
rect 2046 4548 2050 4552
rect 2126 4548 2130 4552
rect 1982 4538 1986 4542
rect 2030 4538 2034 4542
rect 2094 4538 2098 4542
rect 1966 4528 1970 4532
rect 2118 4528 2122 4532
rect 1846 4468 1850 4472
rect 1926 4468 1930 4472
rect 1830 4448 1834 4452
rect 1846 4448 1850 4452
rect 1886 4448 1890 4452
rect 1910 4448 1914 4452
rect 1854 4438 1858 4442
rect 1934 4438 1938 4442
rect 1822 4428 1826 4432
rect 1878 4428 1882 4432
rect 1870 4418 1874 4422
rect 1798 4398 1802 4402
rect 1814 4378 1818 4382
rect 1822 4378 1826 4382
rect 1790 4368 1794 4372
rect 1814 4368 1818 4372
rect 1846 4358 1850 4362
rect 1838 4348 1842 4352
rect 1766 4298 1770 4302
rect 1798 4288 1802 4292
rect 1694 4258 1698 4262
rect 1694 4248 1698 4252
rect 1758 4248 1762 4252
rect 1678 4238 1682 4242
rect 1694 4228 1698 4232
rect 1734 4208 1738 4212
rect 1726 4198 1730 4202
rect 1710 4168 1714 4172
rect 1686 4158 1690 4162
rect 1702 4148 1706 4152
rect 1718 4148 1722 4152
rect 1670 4138 1674 4142
rect 1638 4098 1642 4102
rect 1694 4128 1698 4132
rect 1750 4128 1754 4132
rect 1758 4128 1762 4132
rect 1670 4108 1674 4112
rect 1678 4098 1682 4102
rect 1742 4098 1746 4102
rect 1646 4088 1650 4092
rect 1630 4078 1634 4082
rect 1542 4048 1546 4052
rect 1558 4048 1562 4052
rect 1614 4048 1618 4052
rect 1566 4028 1570 4032
rect 1562 4003 1566 4007
rect 1569 4003 1573 4007
rect 1534 3988 1538 3992
rect 1598 3988 1602 3992
rect 1542 3978 1546 3982
rect 1606 3978 1610 3982
rect 1662 3978 1666 3982
rect 1542 3968 1546 3972
rect 1582 3948 1586 3952
rect 1566 3938 1570 3942
rect 1622 3938 1626 3942
rect 1550 3918 1554 3922
rect 1590 3918 1594 3922
rect 1646 3928 1650 3932
rect 1654 3928 1658 3932
rect 1590 3908 1594 3912
rect 1598 3908 1602 3912
rect 1638 3908 1642 3912
rect 1502 3898 1506 3902
rect 1534 3888 1538 3892
rect 1558 3868 1562 3872
rect 1438 3848 1442 3852
rect 1502 3848 1506 3852
rect 1414 3838 1418 3842
rect 1510 3838 1514 3842
rect 1582 3838 1586 3842
rect 1518 3818 1522 3822
rect 1562 3803 1566 3807
rect 1569 3803 1573 3807
rect 1462 3788 1466 3792
rect 1446 3778 1450 3782
rect 1414 3748 1418 3752
rect 1414 3738 1418 3742
rect 1390 3678 1394 3682
rect 1614 3878 1618 3882
rect 1646 3878 1650 3882
rect 1654 3878 1658 3882
rect 1622 3868 1626 3872
rect 1638 3858 1642 3862
rect 1638 3838 1642 3842
rect 1606 3828 1610 3832
rect 1670 3968 1674 3972
rect 1846 4298 1850 4302
rect 1822 4268 1826 4272
rect 1814 4258 1818 4262
rect 1798 4118 1802 4122
rect 1758 4068 1762 4072
rect 1782 4068 1786 4072
rect 1718 4058 1722 4062
rect 1742 4058 1746 4062
rect 1774 4038 1778 4042
rect 1686 3978 1690 3982
rect 1734 3968 1738 3972
rect 1726 3958 1730 3962
rect 1678 3948 1682 3952
rect 1726 3928 1730 3932
rect 1686 3918 1690 3922
rect 1694 3878 1698 3882
rect 1710 3878 1714 3882
rect 1774 3978 1778 3982
rect 1750 3938 1754 3942
rect 1766 3928 1770 3932
rect 1750 3878 1754 3882
rect 1822 4198 1826 4202
rect 1822 4168 1826 4172
rect 1838 4128 1842 4132
rect 1854 4118 1858 4122
rect 1846 4098 1850 4102
rect 1822 4088 1826 4092
rect 1838 4058 1842 4062
rect 1814 4028 1818 4032
rect 1950 4428 1954 4432
rect 1942 4418 1946 4422
rect 1942 4408 1946 4412
rect 1910 4368 1914 4372
rect 1902 4358 1906 4362
rect 1886 4338 1890 4342
rect 1910 4308 1914 4312
rect 1886 4258 1890 4262
rect 1886 4168 1890 4172
rect 1870 4138 1874 4142
rect 1862 4028 1866 4032
rect 1862 4008 1866 4012
rect 1854 3978 1858 3982
rect 1918 4288 1922 4292
rect 1918 4238 1922 4242
rect 2022 4508 2026 4512
rect 2014 4488 2018 4492
rect 2074 4503 2078 4507
rect 2081 4503 2085 4507
rect 2190 4568 2194 4572
rect 2150 4548 2154 4552
rect 2166 4548 2170 4552
rect 2190 4538 2194 4542
rect 2150 4528 2154 4532
rect 2206 4528 2210 4532
rect 2222 4568 2226 4572
rect 2286 4768 2290 4772
rect 2278 4758 2282 4762
rect 2342 4858 2346 4862
rect 2358 4859 2362 4863
rect 2462 4878 2466 4882
rect 2598 4878 2602 4882
rect 2894 4878 2898 4882
rect 3070 4878 3074 4882
rect 2430 4868 2434 4872
rect 2478 4868 2482 4872
rect 2686 4868 2690 4872
rect 2734 4868 2738 4872
rect 2438 4858 2442 4862
rect 2502 4858 2506 4862
rect 2654 4858 2658 4862
rect 2710 4858 2714 4862
rect 2782 4858 2786 4862
rect 2814 4858 2818 4862
rect 2838 4858 2842 4862
rect 2302 4808 2306 4812
rect 2318 4768 2322 4772
rect 2366 4768 2370 4772
rect 2350 4758 2354 4762
rect 2326 4738 2330 4742
rect 2294 4678 2298 4682
rect 2374 4738 2378 4742
rect 2366 4708 2370 4712
rect 2262 4668 2266 4672
rect 2318 4668 2322 4672
rect 2342 4668 2346 4672
rect 2374 4668 2378 4672
rect 2294 4658 2298 4662
rect 2326 4658 2330 4662
rect 2246 4608 2250 4612
rect 2414 4698 2418 4702
rect 2446 4838 2450 4842
rect 2502 4838 2506 4842
rect 2478 4768 2482 4772
rect 2502 4758 2506 4762
rect 2550 4848 2554 4852
rect 2686 4838 2690 4842
rect 2670 4828 2674 4832
rect 2518 4818 2522 4822
rect 2534 4818 2538 4822
rect 2586 4803 2590 4807
rect 2593 4803 2597 4807
rect 2566 4758 2570 4762
rect 2702 4838 2706 4842
rect 2694 4768 2698 4772
rect 2702 4768 2706 4772
rect 2718 4758 2722 4762
rect 2446 4748 2450 4752
rect 2510 4748 2514 4752
rect 2550 4748 2554 4752
rect 2430 4738 2434 4742
rect 2494 4718 2498 4722
rect 2390 4688 2394 4692
rect 2422 4678 2426 4682
rect 2542 4738 2546 4742
rect 2558 4738 2562 4742
rect 2526 4728 2530 4732
rect 2534 4668 2538 4672
rect 2398 4658 2402 4662
rect 2478 4658 2482 4662
rect 2398 4638 2402 4642
rect 2422 4638 2426 4642
rect 2382 4628 2386 4632
rect 2270 4608 2274 4612
rect 2254 4568 2258 4572
rect 2278 4558 2282 4562
rect 2270 4548 2274 4552
rect 2238 4528 2242 4532
rect 2190 4508 2194 4512
rect 2254 4498 2258 4502
rect 2174 4488 2178 4492
rect 2038 4478 2042 4482
rect 2134 4478 2138 4482
rect 1998 4468 2002 4472
rect 2006 4468 2010 4472
rect 2022 4468 2026 4472
rect 2030 4468 2034 4472
rect 2246 4468 2250 4472
rect 1982 4458 1986 4462
rect 1966 4438 1970 4442
rect 1958 4408 1962 4412
rect 1950 4388 1954 4392
rect 2062 4458 2066 4462
rect 2022 4428 2026 4432
rect 2150 4448 2154 4452
rect 2246 4448 2250 4452
rect 2182 4438 2186 4442
rect 2086 4418 2090 4422
rect 2166 4418 2170 4422
rect 2062 4378 2066 4382
rect 2078 4368 2082 4372
rect 2094 4388 2098 4392
rect 2054 4348 2058 4352
rect 1982 4338 1986 4342
rect 2062 4338 2066 4342
rect 1966 4308 1970 4312
rect 1958 4298 1962 4302
rect 1958 4268 1962 4272
rect 2038 4328 2042 4332
rect 1998 4308 2002 4312
rect 1966 4258 1970 4262
rect 1990 4258 1994 4262
rect 2038 4258 2042 4262
rect 1926 4228 1930 4232
rect 1958 4218 1962 4222
rect 1918 4178 1922 4182
rect 1942 4168 1946 4172
rect 1886 4138 1890 4142
rect 1878 4118 1882 4122
rect 1886 4068 1890 4072
rect 1894 4068 1898 4072
rect 1966 4158 1970 4162
rect 1934 4138 1938 4142
rect 1934 4118 1938 4122
rect 1918 4078 1922 4082
rect 1918 4028 1922 4032
rect 1910 3998 1914 4002
rect 1902 3978 1906 3982
rect 1902 3968 1906 3972
rect 1822 3958 1826 3962
rect 1846 3958 1850 3962
rect 1782 3948 1786 3952
rect 1790 3928 1794 3932
rect 1814 3948 1818 3952
rect 1886 3948 1890 3952
rect 1806 3918 1810 3922
rect 1798 3868 1802 3872
rect 1758 3858 1762 3862
rect 1702 3838 1706 3842
rect 1590 3758 1594 3762
rect 1494 3748 1498 3752
rect 1518 3738 1522 3742
rect 1478 3718 1482 3722
rect 1510 3698 1514 3702
rect 1470 3678 1474 3682
rect 1462 3668 1466 3672
rect 1622 3748 1626 3752
rect 1646 3748 1650 3752
rect 1606 3698 1610 3702
rect 1590 3678 1594 3682
rect 1598 3678 1602 3682
rect 1526 3668 1530 3672
rect 1558 3668 1562 3672
rect 1470 3658 1474 3662
rect 1406 3648 1410 3652
rect 1494 3648 1498 3652
rect 1382 3598 1386 3602
rect 1310 3578 1314 3582
rect 1358 3568 1362 3572
rect 1310 3558 1314 3562
rect 1318 3548 1322 3552
rect 1302 3518 1306 3522
rect 1350 3518 1354 3522
rect 1270 3498 1274 3502
rect 1294 3498 1298 3502
rect 1254 3488 1258 3492
rect 1286 3488 1290 3492
rect 1246 3458 1250 3462
rect 1262 3458 1266 3462
rect 1310 3458 1314 3462
rect 1318 3448 1322 3452
rect 1286 3408 1290 3412
rect 1318 3398 1322 3402
rect 1294 3368 1298 3372
rect 1278 3358 1282 3362
rect 1238 3318 1242 3322
rect 1318 3358 1322 3362
rect 1254 3308 1258 3312
rect 1270 3288 1274 3292
rect 1254 3278 1258 3282
rect 1190 3258 1194 3262
rect 1174 3248 1178 3252
rect 1302 3328 1306 3332
rect 1310 3268 1314 3272
rect 1222 3258 1226 3262
rect 1286 3258 1290 3262
rect 1198 3238 1202 3242
rect 1238 3238 1242 3242
rect 1166 3158 1170 3162
rect 1182 3158 1186 3162
rect 1126 3148 1130 3152
rect 1134 3148 1138 3152
rect 1150 3148 1154 3152
rect 1110 3138 1114 3142
rect 1142 3138 1146 3142
rect 1198 3198 1202 3202
rect 1190 3148 1194 3152
rect 1198 3138 1202 3142
rect 1118 3118 1122 3122
rect 1038 3068 1042 3072
rect 990 3048 994 3052
rect 998 3018 1002 3022
rect 974 3008 978 3012
rect 998 3008 1002 3012
rect 974 2988 978 2992
rect 966 2948 970 2952
rect 862 2928 866 2932
rect 958 2928 962 2932
rect 950 2908 954 2912
rect 862 2898 866 2902
rect 942 2888 946 2892
rect 910 2878 914 2882
rect 902 2868 906 2872
rect 934 2868 938 2872
rect 958 2898 962 2902
rect 1070 3038 1074 3042
rect 1038 3008 1042 3012
rect 1038 2998 1042 3002
rect 1014 2978 1018 2982
rect 1014 2968 1018 2972
rect 1022 2958 1026 2962
rect 1038 2948 1042 2952
rect 1014 2928 1018 2932
rect 1070 2928 1074 2932
rect 1006 2918 1010 2922
rect 998 2878 1002 2882
rect 982 2868 986 2872
rect 782 2858 786 2862
rect 814 2858 818 2862
rect 870 2858 874 2862
rect 758 2848 762 2852
rect 870 2838 874 2842
rect 758 2808 762 2812
rect 790 2798 794 2802
rect 870 2778 874 2782
rect 806 2758 810 2762
rect 854 2758 858 2762
rect 814 2748 818 2752
rect 822 2738 826 2742
rect 814 2728 818 2732
rect 742 2718 746 2722
rect 734 2668 738 2672
rect 726 2628 730 2632
rect 750 2608 754 2612
rect 726 2598 730 2602
rect 718 2588 722 2592
rect 766 2618 770 2622
rect 782 2618 786 2622
rect 758 2598 762 2602
rect 742 2548 746 2552
rect 774 2598 778 2602
rect 774 2538 778 2542
rect 758 2508 762 2512
rect 662 2498 666 2502
rect 702 2498 706 2502
rect 710 2498 714 2502
rect 702 2468 706 2472
rect 758 2468 762 2472
rect 766 2468 770 2472
rect 646 2458 650 2462
rect 662 2458 666 2462
rect 638 2448 642 2452
rect 662 2448 666 2452
rect 654 2418 658 2422
rect 798 2648 802 2652
rect 806 2628 810 2632
rect 790 2598 794 2602
rect 806 2598 810 2602
rect 790 2578 794 2582
rect 782 2448 786 2452
rect 782 2428 786 2432
rect 646 2358 650 2362
rect 766 2358 770 2362
rect 798 2568 802 2572
rect 878 2748 882 2752
rect 870 2738 874 2742
rect 878 2738 882 2742
rect 838 2728 842 2732
rect 862 2728 866 2732
rect 846 2718 850 2722
rect 934 2848 938 2852
rect 982 2848 986 2852
rect 934 2838 938 2842
rect 974 2788 978 2792
rect 958 2778 962 2782
rect 1070 2918 1074 2922
rect 1050 2903 1054 2907
rect 1057 2903 1061 2907
rect 1030 2878 1034 2882
rect 1054 2878 1058 2882
rect 990 2758 994 2762
rect 958 2748 962 2752
rect 974 2738 978 2742
rect 950 2718 954 2722
rect 902 2688 906 2692
rect 838 2678 842 2682
rect 878 2678 882 2682
rect 982 2678 986 2682
rect 838 2658 842 2662
rect 870 2648 874 2652
rect 950 2648 954 2652
rect 846 2638 850 2642
rect 902 2628 906 2632
rect 830 2608 834 2612
rect 822 2578 826 2582
rect 862 2578 866 2582
rect 814 2558 818 2562
rect 846 2558 850 2562
rect 854 2548 858 2552
rect 934 2598 938 2602
rect 902 2578 906 2582
rect 910 2578 914 2582
rect 918 2548 922 2552
rect 830 2538 834 2542
rect 870 2538 874 2542
rect 886 2538 890 2542
rect 798 2528 802 2532
rect 870 2528 874 2532
rect 878 2528 882 2532
rect 798 2488 802 2492
rect 814 2488 818 2492
rect 806 2468 810 2472
rect 870 2478 874 2482
rect 886 2478 890 2482
rect 830 2468 834 2472
rect 830 2458 834 2462
rect 838 2448 842 2452
rect 926 2528 930 2532
rect 982 2658 986 2662
rect 990 2638 994 2642
rect 1046 2788 1050 2792
rect 1094 3048 1098 3052
rect 1102 3038 1106 3042
rect 1094 3028 1098 3032
rect 1118 2958 1122 2962
rect 1118 2948 1122 2952
rect 1110 2938 1114 2942
rect 1094 2898 1098 2902
rect 1086 2888 1090 2892
rect 1094 2878 1098 2882
rect 1110 2868 1114 2872
rect 1102 2858 1106 2862
rect 1126 2858 1130 2862
rect 1078 2838 1082 2842
rect 1182 3128 1186 3132
rect 1174 3098 1178 3102
rect 1166 3088 1170 3092
rect 1142 3078 1146 3082
rect 1222 3178 1226 3182
rect 1238 3158 1242 3162
rect 1238 3138 1242 3142
rect 1262 3158 1266 3162
rect 1286 3248 1290 3252
rect 1302 3208 1306 3212
rect 1286 3178 1290 3182
rect 1318 3178 1322 3182
rect 1302 3168 1306 3172
rect 1286 3148 1290 3152
rect 1270 3118 1274 3122
rect 1238 3108 1242 3112
rect 1246 3108 1250 3112
rect 1206 3088 1210 3092
rect 1286 3128 1290 3132
rect 1334 3498 1338 3502
rect 1438 3628 1442 3632
rect 1478 3598 1482 3602
rect 1462 3568 1466 3572
rect 1486 3568 1490 3572
rect 1374 3548 1378 3552
rect 1486 3548 1490 3552
rect 1358 3488 1362 3492
rect 1390 3498 1394 3502
rect 1406 3488 1410 3492
rect 1358 3478 1362 3482
rect 1374 3478 1378 3482
rect 1470 3528 1474 3532
rect 1478 3528 1482 3532
rect 1430 3518 1434 3522
rect 1454 3518 1458 3522
rect 1462 3508 1466 3512
rect 1422 3498 1426 3502
rect 1358 3468 1362 3472
rect 1342 3448 1346 3452
rect 1414 3468 1418 3472
rect 1382 3448 1386 3452
rect 1398 3448 1402 3452
rect 1366 3438 1370 3442
rect 1382 3438 1386 3442
rect 1350 3428 1354 3432
rect 1414 3418 1418 3422
rect 1414 3378 1418 3382
rect 1406 3368 1410 3372
rect 1358 3358 1362 3362
rect 1438 3458 1442 3462
rect 1430 3448 1434 3452
rect 1454 3428 1458 3432
rect 1430 3398 1434 3402
rect 1462 3378 1466 3382
rect 1430 3348 1434 3352
rect 1334 3278 1338 3282
rect 1310 3108 1314 3112
rect 1326 3108 1330 3112
rect 1326 3088 1330 3092
rect 1278 3078 1282 3082
rect 1214 3068 1218 3072
rect 1222 3068 1226 3072
rect 1198 3058 1202 3062
rect 1286 3058 1290 3062
rect 1294 3058 1298 3062
rect 1182 3048 1186 3052
rect 1198 3018 1202 3022
rect 1142 2998 1146 3002
rect 1158 2978 1162 2982
rect 1150 2948 1154 2952
rect 1158 2948 1162 2952
rect 1190 2948 1194 2952
rect 1150 2938 1154 2942
rect 1150 2928 1154 2932
rect 1182 2928 1186 2932
rect 1270 3038 1274 3042
rect 1286 3038 1290 3042
rect 1230 3028 1234 3032
rect 1254 3028 1258 3032
rect 1238 2998 1242 3002
rect 1222 2918 1226 2922
rect 1166 2858 1170 2862
rect 1142 2848 1146 2852
rect 1222 2888 1226 2892
rect 1182 2868 1186 2872
rect 1230 2868 1234 2872
rect 1190 2858 1194 2862
rect 1134 2788 1138 2792
rect 1062 2748 1066 2752
rect 1078 2748 1082 2752
rect 1046 2738 1050 2742
rect 1102 2738 1106 2742
rect 1046 2718 1050 2722
rect 1050 2703 1054 2707
rect 1057 2703 1061 2707
rect 1070 2698 1074 2702
rect 1046 2678 1050 2682
rect 1014 2658 1018 2662
rect 1030 2658 1034 2662
rect 1062 2658 1066 2662
rect 1006 2608 1010 2612
rect 998 2558 1002 2562
rect 1038 2568 1042 2572
rect 1014 2548 1018 2552
rect 1030 2548 1034 2552
rect 1014 2538 1018 2542
rect 918 2498 922 2502
rect 902 2468 906 2472
rect 894 2458 898 2462
rect 910 2458 914 2462
rect 862 2448 866 2452
rect 886 2448 890 2452
rect 886 2408 890 2412
rect 854 2388 858 2392
rect 814 2368 818 2372
rect 846 2368 850 2372
rect 822 2358 826 2362
rect 846 2358 850 2362
rect 878 2358 882 2362
rect 622 2348 626 2352
rect 638 2338 642 2342
rect 630 2298 634 2302
rect 630 2288 634 2292
rect 614 2278 618 2282
rect 566 2258 570 2262
rect 614 2258 618 2262
rect 606 2248 610 2252
rect 574 2238 578 2242
rect 622 2228 626 2232
rect 598 2198 602 2202
rect 662 2318 666 2322
rect 790 2338 794 2342
rect 766 2328 770 2332
rect 710 2298 714 2302
rect 678 2268 682 2272
rect 646 2258 650 2262
rect 686 2248 690 2252
rect 782 2308 786 2312
rect 726 2258 730 2262
rect 742 2258 746 2262
rect 718 2248 722 2252
rect 702 2238 706 2242
rect 678 2228 682 2232
rect 582 2188 586 2192
rect 678 2188 682 2192
rect 702 2178 706 2182
rect 614 2168 618 2172
rect 646 2168 650 2172
rect 702 2158 706 2162
rect 566 2138 570 2142
rect 606 2148 610 2152
rect 630 2148 634 2152
rect 646 2148 650 2152
rect 686 2148 690 2152
rect 750 2148 754 2152
rect 662 2138 666 2142
rect 590 2128 594 2132
rect 646 2128 650 2132
rect 526 2118 530 2122
rect 558 2118 562 2122
rect 502 2108 506 2112
rect 518 2078 522 2082
rect 534 2078 538 2082
rect 510 2048 514 2052
rect 494 2028 498 2032
rect 518 2008 522 2012
rect 486 1948 490 1952
rect 502 1948 506 1952
rect 538 2003 542 2007
rect 545 2003 549 2007
rect 542 1958 546 1962
rect 486 1928 490 1932
rect 462 1898 466 1902
rect 462 1858 466 1862
rect 454 1838 458 1842
rect 502 1828 506 1832
rect 470 1808 474 1812
rect 446 1798 450 1802
rect 538 1803 542 1807
rect 545 1803 549 1807
rect 470 1788 474 1792
rect 486 1768 490 1772
rect 542 1768 546 1772
rect 430 1758 434 1762
rect 422 1698 426 1702
rect 398 1678 402 1682
rect 334 1668 338 1672
rect 382 1668 386 1672
rect 286 1658 290 1662
rect 334 1658 338 1662
rect 382 1658 386 1662
rect 374 1648 378 1652
rect 366 1608 370 1612
rect 510 1748 514 1752
rect 486 1738 490 1742
rect 494 1738 498 1742
rect 518 1738 522 1742
rect 518 1718 522 1722
rect 494 1698 498 1702
rect 494 1688 498 1692
rect 446 1678 450 1682
rect 470 1678 474 1682
rect 494 1678 498 1682
rect 486 1668 490 1672
rect 510 1668 514 1672
rect 582 2078 586 2082
rect 574 2058 578 2062
rect 646 2098 650 2102
rect 622 2078 626 2082
rect 574 2048 578 2052
rect 598 2048 602 2052
rect 566 1988 570 1992
rect 606 1968 610 1972
rect 622 1958 626 1962
rect 638 1958 642 1962
rect 622 1948 626 1952
rect 566 1938 570 1942
rect 606 1908 610 1912
rect 598 1868 602 1872
rect 654 2018 658 2022
rect 694 2108 698 2112
rect 686 2068 690 2072
rect 678 2048 682 2052
rect 718 2098 722 2102
rect 702 2078 706 2082
rect 774 2278 778 2282
rect 798 2318 802 2322
rect 790 2268 794 2272
rect 806 2268 810 2272
rect 790 2258 794 2262
rect 766 2118 770 2122
rect 774 2088 778 2092
rect 758 2068 762 2072
rect 670 2038 674 2042
rect 686 2038 690 2042
rect 662 2008 666 2012
rect 718 2048 722 2052
rect 742 2048 746 2052
rect 734 2018 738 2022
rect 798 2158 802 2162
rect 830 2298 834 2302
rect 878 2338 882 2342
rect 846 2328 850 2332
rect 854 2298 858 2302
rect 814 2258 818 2262
rect 870 2278 874 2282
rect 934 2508 938 2512
rect 1030 2528 1034 2532
rect 1038 2528 1042 2532
rect 1054 2548 1058 2552
rect 1118 2678 1122 2682
rect 1078 2668 1082 2672
rect 1070 2618 1074 2622
rect 1102 2658 1106 2662
rect 1086 2648 1090 2652
rect 1094 2648 1098 2652
rect 1134 2648 1138 2652
rect 1230 2828 1234 2832
rect 1190 2798 1194 2802
rect 1166 2788 1170 2792
rect 1174 2748 1178 2752
rect 1158 2708 1162 2712
rect 1206 2748 1210 2752
rect 1190 2738 1194 2742
rect 1214 2738 1218 2742
rect 1182 2728 1186 2732
rect 1198 2708 1202 2712
rect 1166 2698 1170 2702
rect 1198 2658 1202 2662
rect 1198 2608 1202 2612
rect 1142 2598 1146 2602
rect 1182 2598 1186 2602
rect 1166 2578 1170 2582
rect 1078 2568 1082 2572
rect 1094 2568 1098 2572
rect 1078 2538 1082 2542
rect 1014 2488 1018 2492
rect 950 2468 954 2472
rect 1050 2503 1054 2507
rect 1057 2503 1061 2507
rect 1054 2488 1058 2492
rect 1038 2458 1042 2462
rect 982 2448 986 2452
rect 1142 2558 1146 2562
rect 1110 2538 1114 2542
rect 1190 2558 1194 2562
rect 1206 2568 1210 2572
rect 1166 2548 1170 2552
rect 1182 2548 1186 2552
rect 1214 2548 1218 2552
rect 1158 2538 1162 2542
rect 1134 2528 1138 2532
rect 1126 2498 1130 2502
rect 1158 2498 1162 2502
rect 1078 2438 1082 2442
rect 1094 2438 1098 2442
rect 942 2388 946 2392
rect 1014 2348 1018 2352
rect 918 2338 922 2342
rect 910 2308 914 2312
rect 894 2268 898 2272
rect 918 2268 922 2272
rect 902 2248 906 2252
rect 846 2238 850 2242
rect 910 2228 914 2232
rect 934 2338 938 2342
rect 958 2298 962 2302
rect 950 2258 954 2262
rect 1050 2303 1054 2307
rect 1057 2303 1061 2307
rect 1046 2278 1050 2282
rect 982 2248 986 2252
rect 846 2218 850 2222
rect 886 2218 890 2222
rect 830 2198 834 2202
rect 814 2178 818 2182
rect 822 2138 826 2142
rect 822 2128 826 2132
rect 814 2118 818 2122
rect 806 2058 810 2062
rect 766 2048 770 2052
rect 790 2048 794 2052
rect 758 2008 762 2012
rect 702 1968 706 1972
rect 710 1958 714 1962
rect 758 1958 762 1962
rect 790 1958 794 1962
rect 798 1958 802 1962
rect 694 1948 698 1952
rect 654 1928 658 1932
rect 678 1928 682 1932
rect 662 1878 666 1882
rect 654 1868 658 1872
rect 702 1868 706 1872
rect 566 1858 570 1862
rect 646 1858 650 1862
rect 574 1748 578 1752
rect 430 1658 434 1662
rect 470 1658 474 1662
rect 454 1648 458 1652
rect 486 1638 490 1642
rect 538 1603 542 1607
rect 545 1603 549 1607
rect 422 1578 426 1582
rect 366 1558 370 1562
rect 278 1538 282 1542
rect 326 1538 330 1542
rect 334 1528 338 1532
rect 278 1518 282 1522
rect 270 1508 274 1512
rect 342 1498 346 1502
rect 550 1558 554 1562
rect 406 1548 410 1552
rect 438 1548 442 1552
rect 446 1538 450 1542
rect 422 1518 426 1522
rect 422 1508 426 1512
rect 390 1498 394 1502
rect 262 1488 266 1492
rect 294 1478 298 1482
rect 166 1408 170 1412
rect 270 1468 274 1472
rect 214 1448 218 1452
rect 222 1428 226 1432
rect 246 1458 250 1462
rect 278 1458 282 1462
rect 238 1428 242 1432
rect 198 1398 202 1402
rect 230 1398 234 1402
rect 222 1368 226 1372
rect 190 1318 194 1322
rect 254 1428 258 1432
rect 366 1448 370 1452
rect 366 1428 370 1432
rect 310 1418 314 1422
rect 302 1398 306 1402
rect 334 1398 338 1402
rect 278 1388 282 1392
rect 294 1368 298 1372
rect 294 1348 298 1352
rect 254 1338 258 1342
rect 254 1318 258 1322
rect 278 1318 282 1322
rect 166 1288 170 1292
rect 198 1288 202 1292
rect 182 1278 186 1282
rect 278 1308 282 1312
rect 230 1268 234 1272
rect 150 1148 154 1152
rect 134 1068 138 1072
rect 230 1248 234 1252
rect 214 1238 218 1242
rect 238 1238 242 1242
rect 166 1228 170 1232
rect 166 1208 170 1212
rect 198 1178 202 1182
rect 190 1168 194 1172
rect 182 1148 186 1152
rect 126 1058 130 1062
rect 102 988 106 992
rect 110 948 114 952
rect 62 938 66 942
rect 102 888 106 892
rect 110 868 114 872
rect 46 858 50 862
rect 118 848 122 852
rect 134 1018 138 1022
rect 134 988 138 992
rect 182 1068 186 1072
rect 206 1168 210 1172
rect 214 1158 218 1162
rect 246 1148 250 1152
rect 214 1088 218 1092
rect 166 1048 170 1052
rect 182 1048 186 1052
rect 198 1048 202 1052
rect 214 1038 218 1042
rect 198 1028 202 1032
rect 214 1008 218 1012
rect 198 988 202 992
rect 158 978 162 982
rect 134 958 138 962
rect 134 888 138 892
rect 198 968 202 972
rect 206 968 210 972
rect 174 938 178 942
rect 150 868 154 872
rect 134 828 138 832
rect 54 798 58 802
rect 110 798 114 802
rect 126 798 130 802
rect 38 728 42 732
rect 14 668 18 672
rect 38 558 42 562
rect 14 488 18 492
rect 30 468 34 472
rect 38 458 42 462
rect 110 748 114 752
rect 134 748 138 752
rect 94 738 98 742
rect 70 708 74 712
rect 150 738 154 742
rect 118 718 122 722
rect 102 698 106 702
rect 126 698 130 702
rect 86 678 90 682
rect 118 658 122 662
rect 102 568 106 572
rect 118 558 122 562
rect 94 538 98 542
rect 94 528 98 532
rect 62 518 66 522
rect 86 478 90 482
rect 46 288 50 292
rect 102 508 106 512
rect 102 468 106 472
rect 78 458 82 462
rect 150 568 154 572
rect 134 558 138 562
rect 214 878 218 882
rect 174 848 178 852
rect 198 848 202 852
rect 166 728 170 732
rect 182 818 186 822
rect 198 778 202 782
rect 270 1128 274 1132
rect 246 1118 250 1122
rect 230 1068 234 1072
rect 294 1138 298 1142
rect 238 1058 242 1062
rect 230 988 234 992
rect 222 808 226 812
rect 206 768 210 772
rect 182 748 186 752
rect 222 748 226 752
rect 174 718 178 722
rect 174 698 178 702
rect 262 998 266 1002
rect 278 1038 282 1042
rect 270 968 274 972
rect 262 938 266 942
rect 254 928 258 932
rect 246 918 250 922
rect 246 858 250 862
rect 238 788 242 792
rect 238 758 242 762
rect 262 758 266 762
rect 286 878 290 882
rect 310 1388 314 1392
rect 326 1358 330 1362
rect 382 1388 386 1392
rect 350 1358 354 1362
rect 350 1348 354 1352
rect 350 1338 354 1342
rect 350 1328 354 1332
rect 334 1298 338 1302
rect 366 1318 370 1322
rect 358 1308 362 1312
rect 510 1547 514 1551
rect 454 1518 458 1522
rect 470 1518 474 1522
rect 462 1498 466 1502
rect 398 1478 402 1482
rect 422 1478 426 1482
rect 406 1418 410 1422
rect 398 1398 402 1402
rect 374 1298 378 1302
rect 358 1288 362 1292
rect 366 1288 370 1292
rect 446 1468 450 1472
rect 430 1448 434 1452
rect 422 1388 426 1392
rect 430 1368 434 1372
rect 406 1348 410 1352
rect 422 1348 426 1352
rect 414 1338 418 1342
rect 350 1258 354 1262
rect 382 1258 386 1262
rect 334 1248 338 1252
rect 390 1238 394 1242
rect 406 1228 410 1232
rect 398 1218 402 1222
rect 374 1188 378 1192
rect 390 1188 394 1192
rect 382 1178 386 1182
rect 366 1128 370 1132
rect 326 1078 330 1082
rect 342 1078 346 1082
rect 318 988 322 992
rect 342 1068 346 1072
rect 350 1068 354 1072
rect 406 1088 410 1092
rect 518 1498 522 1502
rect 486 1488 490 1492
rect 494 1488 498 1492
rect 462 1448 466 1452
rect 454 1398 458 1402
rect 526 1418 530 1422
rect 538 1403 542 1407
rect 545 1403 549 1407
rect 478 1388 482 1392
rect 518 1388 522 1392
rect 462 1358 466 1362
rect 470 1347 474 1351
rect 526 1328 530 1332
rect 462 1318 466 1322
rect 462 1308 466 1312
rect 446 1278 450 1282
rect 454 1268 458 1272
rect 446 1248 450 1252
rect 510 1298 514 1302
rect 486 1288 490 1292
rect 470 1258 474 1262
rect 486 1258 490 1262
rect 502 1228 506 1232
rect 430 1188 434 1192
rect 438 1188 442 1192
rect 470 1158 474 1162
rect 550 1278 554 1282
rect 534 1248 538 1252
rect 574 1708 578 1712
rect 574 1668 578 1672
rect 606 1668 610 1672
rect 638 1738 642 1742
rect 662 1859 666 1863
rect 790 1948 794 1952
rect 774 1938 778 1942
rect 798 1938 802 1942
rect 734 1908 738 1912
rect 758 1908 762 1912
rect 750 1888 754 1892
rect 758 1868 762 1872
rect 718 1858 722 1862
rect 710 1848 714 1852
rect 734 1848 738 1852
rect 782 1908 786 1912
rect 870 2188 874 2192
rect 846 2158 850 2162
rect 854 2158 858 2162
rect 838 2078 842 2082
rect 926 2218 930 2222
rect 918 2198 922 2202
rect 918 2188 922 2192
rect 934 2188 938 2192
rect 982 2178 986 2182
rect 942 2158 946 2162
rect 958 2158 962 2162
rect 910 2148 914 2152
rect 894 2138 898 2142
rect 902 2138 906 2142
rect 862 2128 866 2132
rect 886 2108 890 2112
rect 886 2098 890 2102
rect 854 2078 858 2082
rect 830 2018 834 2022
rect 846 2018 850 2022
rect 822 1948 826 1952
rect 814 1928 818 1932
rect 798 1918 802 1922
rect 806 1918 810 1922
rect 790 1888 794 1892
rect 790 1868 794 1872
rect 798 1868 802 1872
rect 774 1858 778 1862
rect 766 1848 770 1852
rect 782 1838 786 1842
rect 838 2008 842 2012
rect 854 1908 858 1912
rect 902 2028 906 2032
rect 910 2028 914 2032
rect 894 1968 898 1972
rect 878 1958 882 1962
rect 886 1958 890 1962
rect 942 2138 946 2142
rect 974 2138 978 2142
rect 1022 2138 1026 2142
rect 974 2128 978 2132
rect 990 2128 994 2132
rect 982 2108 986 2112
rect 1050 2103 1054 2107
rect 1057 2103 1061 2107
rect 1006 2098 1010 2102
rect 1030 2068 1034 2072
rect 990 2058 994 2062
rect 974 2048 978 2052
rect 974 2038 978 2042
rect 982 2018 986 2022
rect 926 1958 930 1962
rect 838 1878 842 1882
rect 886 1858 890 1862
rect 814 1848 818 1852
rect 798 1828 802 1832
rect 750 1818 754 1822
rect 702 1758 706 1762
rect 710 1758 714 1762
rect 734 1758 738 1762
rect 686 1738 690 1742
rect 814 1798 818 1802
rect 838 1798 842 1802
rect 870 1778 874 1782
rect 774 1758 778 1762
rect 718 1748 722 1752
rect 758 1748 762 1752
rect 878 1768 882 1772
rect 734 1738 738 1742
rect 742 1738 746 1742
rect 694 1728 698 1732
rect 718 1728 722 1732
rect 678 1718 682 1722
rect 686 1718 690 1722
rect 702 1718 706 1722
rect 686 1668 690 1672
rect 614 1658 618 1662
rect 670 1658 674 1662
rect 582 1648 586 1652
rect 598 1648 602 1652
rect 590 1608 594 1612
rect 614 1638 618 1642
rect 654 1648 658 1652
rect 662 1648 666 1652
rect 710 1648 714 1652
rect 606 1628 610 1632
rect 622 1628 626 1632
rect 646 1598 650 1602
rect 614 1568 618 1572
rect 662 1638 666 1642
rect 670 1638 674 1642
rect 710 1638 714 1642
rect 686 1608 690 1612
rect 670 1588 674 1592
rect 662 1558 666 1562
rect 598 1548 602 1552
rect 566 1538 570 1542
rect 582 1538 586 1542
rect 638 1538 642 1542
rect 566 1528 570 1532
rect 574 1488 578 1492
rect 566 1398 570 1402
rect 654 1518 658 1522
rect 622 1498 626 1502
rect 630 1488 634 1492
rect 606 1468 610 1472
rect 598 1458 602 1462
rect 646 1448 650 1452
rect 606 1438 610 1442
rect 614 1438 618 1442
rect 598 1368 602 1372
rect 574 1348 578 1352
rect 606 1348 610 1352
rect 606 1338 610 1342
rect 574 1328 578 1332
rect 598 1318 602 1322
rect 574 1288 578 1292
rect 590 1278 594 1282
rect 558 1208 562 1212
rect 538 1203 542 1207
rect 545 1203 549 1207
rect 590 1168 594 1172
rect 582 1158 586 1162
rect 630 1388 634 1392
rect 622 1348 626 1352
rect 686 1558 690 1562
rect 670 1518 674 1522
rect 670 1468 674 1472
rect 702 1468 706 1472
rect 654 1408 658 1412
rect 662 1368 666 1372
rect 646 1358 650 1362
rect 694 1458 698 1462
rect 702 1428 706 1432
rect 678 1408 682 1412
rect 678 1368 682 1372
rect 662 1298 666 1302
rect 694 1338 698 1342
rect 766 1708 770 1712
rect 758 1688 762 1692
rect 734 1638 738 1642
rect 726 1598 730 1602
rect 734 1508 738 1512
rect 758 1618 762 1622
rect 950 1958 954 1962
rect 1006 2048 1010 2052
rect 1022 2048 1026 2052
rect 998 1998 1002 2002
rect 1014 1998 1018 2002
rect 1014 1958 1018 1962
rect 966 1948 970 1952
rect 982 1948 986 1952
rect 926 1938 930 1942
rect 918 1838 922 1842
rect 902 1738 906 1742
rect 894 1728 898 1732
rect 886 1708 890 1712
rect 782 1678 786 1682
rect 822 1678 826 1682
rect 806 1658 810 1662
rect 790 1628 794 1632
rect 814 1628 818 1632
rect 782 1618 786 1622
rect 774 1608 778 1612
rect 782 1598 786 1602
rect 774 1578 778 1582
rect 774 1558 778 1562
rect 782 1548 786 1552
rect 766 1508 770 1512
rect 1038 2038 1042 2042
rect 1054 2038 1058 2042
rect 1166 2428 1170 2432
rect 1182 2498 1186 2502
rect 1182 2468 1186 2472
rect 1270 2948 1274 2952
rect 1246 2938 1250 2942
rect 1310 3058 1314 3062
rect 1478 3428 1482 3432
rect 1358 3338 1362 3342
rect 1454 3338 1458 3342
rect 1358 3318 1362 3322
rect 1446 3318 1450 3322
rect 1414 3258 1418 3262
rect 1366 3228 1370 3232
rect 1374 3188 1378 3192
rect 1358 3078 1362 3082
rect 1342 3068 1346 3072
rect 1382 3158 1386 3162
rect 1478 3288 1482 3292
rect 1574 3658 1578 3662
rect 1526 3648 1530 3652
rect 1614 3658 1618 3662
rect 1526 3628 1530 3632
rect 1582 3628 1586 3632
rect 1590 3628 1594 3632
rect 1526 3618 1530 3622
rect 1510 3508 1514 3512
rect 1502 3498 1506 3502
rect 1502 3478 1506 3482
rect 1562 3603 1566 3607
rect 1569 3603 1573 3607
rect 1598 3618 1602 3622
rect 1606 3568 1610 3572
rect 1590 3548 1594 3552
rect 1550 3518 1554 3522
rect 1582 3488 1586 3492
rect 1502 3458 1506 3462
rect 1550 3458 1554 3462
rect 1534 3398 1538 3402
rect 1526 3378 1530 3382
rect 1494 3358 1498 3362
rect 1502 3358 1506 3362
rect 1562 3403 1566 3407
rect 1569 3403 1573 3407
rect 1542 3388 1546 3392
rect 1550 3378 1554 3382
rect 1574 3378 1578 3382
rect 1494 3338 1498 3342
rect 1638 3738 1642 3742
rect 1742 3848 1746 3852
rect 1710 3828 1714 3832
rect 1694 3768 1698 3772
rect 1670 3748 1674 3752
rect 1686 3748 1690 3752
rect 1662 3658 1666 3662
rect 1654 3608 1658 3612
rect 1622 3568 1626 3572
rect 1630 3548 1634 3552
rect 1606 3478 1610 3482
rect 1606 3458 1610 3462
rect 1614 3448 1618 3452
rect 1662 3598 1666 3602
rect 1726 3768 1730 3772
rect 1718 3738 1722 3742
rect 1718 3718 1722 3722
rect 1726 3708 1730 3712
rect 1726 3688 1730 3692
rect 1702 3678 1706 3682
rect 1798 3838 1802 3842
rect 1822 3878 1826 3882
rect 1814 3868 1818 3872
rect 1806 3828 1810 3832
rect 1830 3818 1834 3822
rect 1750 3778 1754 3782
rect 1766 3778 1770 3782
rect 1766 3768 1770 3772
rect 1750 3758 1754 3762
rect 1766 3718 1770 3722
rect 1742 3698 1746 3702
rect 1758 3688 1762 3692
rect 1678 3648 1682 3652
rect 1694 3558 1698 3562
rect 1686 3548 1690 3552
rect 1686 3528 1690 3532
rect 1710 3528 1714 3532
rect 1718 3528 1722 3532
rect 1678 3478 1682 3482
rect 1678 3438 1682 3442
rect 1694 3488 1698 3492
rect 1694 3448 1698 3452
rect 1654 3428 1658 3432
rect 1686 3428 1690 3432
rect 1638 3408 1642 3412
rect 1598 3398 1602 3402
rect 1630 3398 1634 3402
rect 1526 3338 1530 3342
rect 1606 3338 1610 3342
rect 1510 3328 1514 3332
rect 1478 3268 1482 3272
rect 1486 3268 1490 3272
rect 1494 3258 1498 3262
rect 1470 3228 1474 3232
rect 1518 3248 1522 3252
rect 1502 3228 1506 3232
rect 1486 3198 1490 3202
rect 1478 3188 1482 3192
rect 1470 3158 1474 3162
rect 1382 3128 1386 3132
rect 1422 3128 1426 3132
rect 1446 3128 1450 3132
rect 1350 3058 1354 3062
rect 1374 3058 1378 3062
rect 1398 3118 1402 3122
rect 1406 3118 1410 3122
rect 1422 3088 1426 3092
rect 1542 3318 1546 3322
rect 1598 3288 1602 3292
rect 1534 3178 1538 3182
rect 1494 3158 1498 3162
rect 1502 3148 1506 3152
rect 1526 3148 1530 3152
rect 1510 3138 1514 3142
rect 1526 3128 1530 3132
rect 1398 3078 1402 3082
rect 1430 3078 1434 3082
rect 1478 3078 1482 3082
rect 1390 3068 1394 3072
rect 1534 3118 1538 3122
rect 1534 3088 1538 3092
rect 1446 3068 1450 3072
rect 1510 3068 1514 3072
rect 1366 2988 1370 2992
rect 1562 3203 1566 3207
rect 1569 3203 1573 3207
rect 1550 3158 1554 3162
rect 1582 3158 1586 3162
rect 1590 3158 1594 3162
rect 1582 3138 1586 3142
rect 1542 3078 1546 3082
rect 1454 3058 1458 3062
rect 1486 3048 1490 3052
rect 1462 2998 1466 3002
rect 1438 2978 1442 2982
rect 1358 2968 1362 2972
rect 1350 2958 1354 2962
rect 1366 2958 1370 2962
rect 1334 2948 1338 2952
rect 1374 2948 1378 2952
rect 1310 2938 1314 2942
rect 1342 2938 1346 2942
rect 1302 2928 1306 2932
rect 1294 2918 1298 2922
rect 1350 2918 1354 2922
rect 1302 2888 1306 2892
rect 1342 2888 1346 2892
rect 1318 2868 1322 2872
rect 1270 2848 1274 2852
rect 1278 2838 1282 2842
rect 1406 2938 1410 2942
rect 1414 2938 1418 2942
rect 1430 2928 1434 2932
rect 1414 2918 1418 2922
rect 1358 2888 1362 2892
rect 1342 2848 1346 2852
rect 1334 2838 1338 2842
rect 1302 2828 1306 2832
rect 1294 2768 1298 2772
rect 1270 2758 1274 2762
rect 1382 2848 1386 2852
rect 1390 2848 1394 2852
rect 1350 2838 1354 2842
rect 1390 2798 1394 2802
rect 1350 2758 1354 2762
rect 1238 2748 1242 2752
rect 1254 2748 1258 2752
rect 1342 2748 1346 2752
rect 1262 2728 1266 2732
rect 1254 2708 1258 2712
rect 1278 2708 1282 2712
rect 1358 2708 1362 2712
rect 1238 2668 1242 2672
rect 1254 2658 1258 2662
rect 1270 2648 1274 2652
rect 1230 2608 1234 2612
rect 1230 2528 1234 2532
rect 1262 2508 1266 2512
rect 1246 2458 1250 2462
rect 1230 2448 1234 2452
rect 1238 2448 1242 2452
rect 1206 2418 1210 2422
rect 1222 2418 1226 2422
rect 1174 2408 1178 2412
rect 1182 2388 1186 2392
rect 1198 2368 1202 2372
rect 1214 2368 1218 2372
rect 1102 2358 1106 2362
rect 1206 2358 1210 2362
rect 1110 2348 1114 2352
rect 1126 2348 1130 2352
rect 1214 2348 1218 2352
rect 1102 2338 1106 2342
rect 1118 2338 1122 2342
rect 1150 2338 1154 2342
rect 1110 2278 1114 2282
rect 1102 2268 1106 2272
rect 1110 2258 1114 2262
rect 1078 2228 1082 2232
rect 1086 2158 1090 2162
rect 1118 2238 1122 2242
rect 1118 2178 1122 2182
rect 1118 2158 1122 2162
rect 1150 2328 1154 2332
rect 1158 2328 1162 2332
rect 1238 2338 1242 2342
rect 1174 2308 1178 2312
rect 1198 2278 1202 2282
rect 1174 2268 1178 2272
rect 1230 2298 1234 2302
rect 1254 2378 1258 2382
rect 1246 2268 1250 2272
rect 1198 2258 1202 2262
rect 1150 2248 1154 2252
rect 1214 2258 1218 2262
rect 1230 2258 1234 2262
rect 1166 2228 1170 2232
rect 1238 2228 1242 2232
rect 1206 2218 1210 2222
rect 1214 2218 1218 2222
rect 1174 2188 1178 2192
rect 1134 2178 1138 2182
rect 1150 2178 1154 2182
rect 1134 2158 1138 2162
rect 1182 2158 1186 2162
rect 1126 2148 1130 2152
rect 1134 2138 1138 2142
rect 1126 2128 1130 2132
rect 1094 2108 1098 2112
rect 1094 2078 1098 2082
rect 1110 2058 1114 2062
rect 1126 2058 1130 2062
rect 1102 2038 1106 2042
rect 1110 2038 1114 2042
rect 1038 2028 1042 2032
rect 1070 2028 1074 2032
rect 1030 2018 1034 2022
rect 1054 2008 1058 2012
rect 1110 2008 1114 2012
rect 1118 1998 1122 2002
rect 1166 2088 1170 2092
rect 1150 2078 1154 2082
rect 1166 2078 1170 2082
rect 1190 2078 1194 2082
rect 1246 2188 1250 2192
rect 1294 2648 1298 2652
rect 1286 2598 1290 2602
rect 1350 2568 1354 2572
rect 1278 2558 1282 2562
rect 1342 2548 1346 2552
rect 1302 2538 1306 2542
rect 1350 2508 1354 2512
rect 1302 2488 1306 2492
rect 1278 2468 1282 2472
rect 1294 2468 1298 2472
rect 1286 2448 1290 2452
rect 1342 2448 1346 2452
rect 1302 2428 1306 2432
rect 1286 2408 1290 2412
rect 1310 2408 1314 2412
rect 1318 2408 1322 2412
rect 1278 2388 1282 2392
rect 1286 2388 1290 2392
rect 1310 2378 1314 2382
rect 1278 2368 1282 2372
rect 1286 2368 1290 2372
rect 1374 2668 1378 2672
rect 1406 2708 1410 2712
rect 1462 2908 1466 2912
rect 1446 2878 1450 2882
rect 1446 2868 1450 2872
rect 1502 3018 1506 3022
rect 1606 3259 1610 3263
rect 1614 3248 1618 3252
rect 1606 3238 1610 3242
rect 1614 3198 1618 3202
rect 1702 3428 1706 3432
rect 1662 3378 1666 3382
rect 1638 3368 1642 3372
rect 1678 3358 1682 3362
rect 1670 3278 1674 3282
rect 1654 3258 1658 3262
rect 1662 3248 1666 3252
rect 1646 3238 1650 3242
rect 1670 3228 1674 3232
rect 1686 3328 1690 3332
rect 1694 3288 1698 3292
rect 1686 3198 1690 3202
rect 1662 3188 1666 3192
rect 1678 3188 1682 3192
rect 1710 3418 1714 3422
rect 1710 3288 1714 3292
rect 1734 3658 1738 3662
rect 1742 3598 1746 3602
rect 1734 3458 1738 3462
rect 1726 3428 1730 3432
rect 1782 3678 1786 3682
rect 1822 3778 1826 3782
rect 1814 3748 1818 3752
rect 1846 3878 1850 3882
rect 1854 3868 1858 3872
rect 1846 3808 1850 3812
rect 1854 3798 1858 3802
rect 1854 3788 1858 3792
rect 1878 3928 1882 3932
rect 1878 3878 1882 3882
rect 1886 3878 1890 3882
rect 1886 3868 1890 3872
rect 1998 4168 2002 4172
rect 1998 4158 2002 4162
rect 1998 4148 2002 4152
rect 2022 4128 2026 4132
rect 2074 4303 2078 4307
rect 2081 4303 2085 4307
rect 2062 4278 2066 4282
rect 2086 4238 2090 4242
rect 2046 4218 2050 4222
rect 2062 4158 2066 4162
rect 2142 4378 2146 4382
rect 2118 4368 2122 4372
rect 2134 4368 2138 4372
rect 2118 4348 2122 4352
rect 2158 4348 2162 4352
rect 2142 4328 2146 4332
rect 2190 4368 2194 4372
rect 2214 4368 2218 4372
rect 2174 4328 2178 4332
rect 2174 4318 2178 4322
rect 2134 4278 2138 4282
rect 2150 4278 2154 4282
rect 2166 4278 2170 4282
rect 2150 4258 2154 4262
rect 2190 4298 2194 4302
rect 2214 4288 2218 4292
rect 2262 4438 2266 4442
rect 2278 4508 2282 4512
rect 2390 4558 2394 4562
rect 2358 4538 2362 4542
rect 2374 4538 2378 4542
rect 2342 4528 2346 4532
rect 2358 4528 2362 4532
rect 2278 4468 2282 4472
rect 2294 4458 2298 4462
rect 2350 4498 2354 4502
rect 2302 4438 2306 4442
rect 2326 4438 2330 4442
rect 2334 4438 2338 4442
rect 2278 4318 2282 4322
rect 2302 4318 2306 4322
rect 2246 4298 2250 4302
rect 2270 4298 2274 4302
rect 2222 4278 2226 4282
rect 2238 4268 2242 4272
rect 2182 4258 2186 4262
rect 2198 4258 2202 4262
rect 2414 4618 2418 4622
rect 2526 4618 2530 4622
rect 2630 4747 2634 4751
rect 2686 4728 2690 4732
rect 2694 4718 2698 4722
rect 2694 4688 2698 4692
rect 2558 4668 2562 4672
rect 2630 4668 2634 4672
rect 2654 4668 2658 4672
rect 2550 4658 2554 4662
rect 2574 4638 2578 4642
rect 2694 4658 2698 4662
rect 2582 4628 2586 4632
rect 2718 4738 2722 4742
rect 2742 4828 2746 4832
rect 2726 4698 2730 4702
rect 2726 4658 2730 4662
rect 2718 4628 2722 4632
rect 2586 4603 2590 4607
rect 2593 4603 2597 4607
rect 2542 4598 2546 4602
rect 2534 4578 2538 4582
rect 2694 4578 2698 4582
rect 2726 4588 2730 4592
rect 2710 4578 2714 4582
rect 2590 4568 2594 4572
rect 2702 4568 2706 4572
rect 2422 4558 2426 4562
rect 2470 4558 2474 4562
rect 2462 4548 2466 4552
rect 2486 4548 2490 4552
rect 2518 4548 2522 4552
rect 2534 4548 2538 4552
rect 2454 4538 2458 4542
rect 2454 4518 2458 4522
rect 2430 4508 2434 4512
rect 2446 4508 2450 4512
rect 2414 4468 2418 4472
rect 2502 4528 2506 4532
rect 2462 4498 2466 4502
rect 2486 4468 2490 4472
rect 2358 4458 2362 4462
rect 2422 4458 2426 4462
rect 2390 4438 2394 4442
rect 2342 4318 2346 4322
rect 2270 4288 2274 4292
rect 2446 4378 2450 4382
rect 2390 4368 2394 4372
rect 2414 4368 2418 4372
rect 2446 4348 2450 4352
rect 2478 4428 2482 4432
rect 2574 4548 2578 4552
rect 2718 4568 2722 4572
rect 2614 4547 2618 4551
rect 2694 4548 2698 4552
rect 2670 4538 2674 4542
rect 2574 4518 2578 4522
rect 2518 4488 2522 4492
rect 2534 4488 2538 4492
rect 2534 4468 2538 4472
rect 2550 4468 2554 4472
rect 2518 4458 2522 4462
rect 2510 4448 2514 4452
rect 2686 4528 2690 4532
rect 2662 4518 2666 4522
rect 2670 4488 2674 4492
rect 2694 4468 2698 4472
rect 2614 4438 2618 4442
rect 2542 4418 2546 4422
rect 2494 4398 2498 4402
rect 2510 4378 2514 4382
rect 2462 4358 2466 4362
rect 2486 4358 2490 4362
rect 2526 4358 2530 4362
rect 2542 4358 2546 4362
rect 2694 4428 2698 4432
rect 2718 4508 2722 4512
rect 2854 4818 2858 4822
rect 2750 4768 2754 4772
rect 2750 4758 2754 4762
rect 2814 4758 2818 4762
rect 2758 4738 2762 4742
rect 2838 4738 2842 4742
rect 2958 4858 2962 4862
rect 2982 4858 2986 4862
rect 3014 4858 3018 4862
rect 3086 4858 3090 4862
rect 3054 4838 3058 4842
rect 2894 4798 2898 4802
rect 3062 4758 3066 4762
rect 2742 4698 2746 4702
rect 2862 4688 2866 4692
rect 2742 4658 2746 4662
rect 2974 4728 2978 4732
rect 3038 4728 3042 4732
rect 2998 4718 3002 4722
rect 2902 4708 2906 4712
rect 2782 4658 2786 4662
rect 2878 4658 2882 4662
rect 2798 4648 2802 4652
rect 2742 4638 2746 4642
rect 2766 4638 2770 4642
rect 2854 4638 2858 4642
rect 2902 4638 2906 4642
rect 2790 4548 2794 4552
rect 3030 4708 3034 4712
rect 3014 4688 3018 4692
rect 2982 4658 2986 4662
rect 2982 4648 2986 4652
rect 2998 4648 3002 4652
rect 2958 4598 2962 4602
rect 2870 4568 2874 4572
rect 2862 4558 2866 4562
rect 2798 4538 2802 4542
rect 2862 4538 2866 4542
rect 2742 4488 2746 4492
rect 2790 4488 2794 4492
rect 2734 4478 2738 4482
rect 2822 4508 2826 4512
rect 2814 4498 2818 4502
rect 2742 4468 2746 4472
rect 2774 4468 2778 4472
rect 2806 4468 2810 4472
rect 2726 4458 2730 4462
rect 2710 4418 2714 4422
rect 2586 4403 2590 4407
rect 2593 4403 2597 4407
rect 2662 4388 2666 4392
rect 2694 4368 2698 4372
rect 2710 4368 2714 4372
rect 2718 4368 2722 4372
rect 2470 4348 2474 4352
rect 2502 4348 2506 4352
rect 2454 4328 2458 4332
rect 2462 4328 2466 4332
rect 2486 4328 2490 4332
rect 2422 4308 2426 4312
rect 2398 4298 2402 4302
rect 2406 4298 2410 4302
rect 2382 4288 2386 4292
rect 2350 4278 2354 4282
rect 2366 4278 2370 4282
rect 2302 4268 2306 4272
rect 2374 4268 2378 4272
rect 2278 4258 2282 4262
rect 2310 4258 2314 4262
rect 2382 4258 2386 4262
rect 2110 4248 2114 4252
rect 2182 4238 2186 4242
rect 2126 4138 2130 4142
rect 2038 4118 2042 4122
rect 1982 4108 1986 4112
rect 1990 4108 1994 4112
rect 2074 4103 2078 4107
rect 2081 4103 2085 4107
rect 1990 4088 1994 4092
rect 1998 4088 2002 4092
rect 1958 4048 1962 4052
rect 1942 4028 1946 4032
rect 1950 4028 1954 4032
rect 1934 3988 1938 3992
rect 1958 4008 1962 4012
rect 2158 4148 2162 4152
rect 2174 4148 2178 4152
rect 2134 4128 2138 4132
rect 2142 4118 2146 4122
rect 2158 4098 2162 4102
rect 2006 4048 2010 4052
rect 2022 4048 2026 4052
rect 2078 4048 2082 4052
rect 1982 4018 1986 4022
rect 2022 4008 2026 4012
rect 1966 3988 1970 3992
rect 1974 3978 1978 3982
rect 2086 3978 2090 3982
rect 1958 3958 1962 3962
rect 1942 3948 1946 3952
rect 1998 3958 2002 3962
rect 2022 3958 2026 3962
rect 1990 3948 1994 3952
rect 2014 3948 2018 3952
rect 2046 3948 2050 3952
rect 2006 3938 2010 3942
rect 2022 3938 2026 3942
rect 2054 3938 2058 3942
rect 1934 3888 1938 3892
rect 2078 3918 2082 3922
rect 2110 3918 2114 3922
rect 2074 3903 2078 3907
rect 2081 3903 2085 3907
rect 2102 3898 2106 3902
rect 2022 3888 2026 3892
rect 1990 3868 1994 3872
rect 2062 3868 2066 3872
rect 1870 3858 1874 3862
rect 2038 3858 2042 3862
rect 2086 3858 2090 3862
rect 1878 3848 1882 3852
rect 2070 3828 2074 3832
rect 2110 3828 2114 3832
rect 1926 3818 1930 3822
rect 1878 3758 1882 3762
rect 1894 3758 1898 3762
rect 1838 3738 1842 3742
rect 1862 3738 1866 3742
rect 1870 3718 1874 3722
rect 1806 3698 1810 3702
rect 1798 3688 1802 3692
rect 1782 3648 1786 3652
rect 1774 3598 1778 3602
rect 1774 3558 1778 3562
rect 1790 3548 1794 3552
rect 1846 3688 1850 3692
rect 1886 3688 1890 3692
rect 1814 3678 1818 3682
rect 1854 3678 1858 3682
rect 1846 3668 1850 3672
rect 1910 3758 1914 3762
rect 1902 3678 1906 3682
rect 1902 3668 1906 3672
rect 1822 3658 1826 3662
rect 1894 3658 1898 3662
rect 1838 3648 1842 3652
rect 1822 3618 1826 3622
rect 1814 3568 1818 3572
rect 1814 3518 1818 3522
rect 1750 3378 1754 3382
rect 1774 3398 1778 3402
rect 1838 3598 1842 3602
rect 1846 3588 1850 3592
rect 2014 3768 2018 3772
rect 1958 3758 1962 3762
rect 2038 3758 2042 3762
rect 2054 3758 2058 3762
rect 2134 4038 2138 4042
rect 2206 4198 2210 4202
rect 2230 4158 2234 4162
rect 2214 4098 2218 4102
rect 2174 4088 2178 4092
rect 2190 4088 2194 4092
rect 2158 4058 2162 4062
rect 2150 4028 2154 4032
rect 2126 3928 2130 3932
rect 2126 3868 2130 3872
rect 2142 3868 2146 3872
rect 2158 3848 2162 3852
rect 2222 4088 2226 4092
rect 2190 4058 2194 4062
rect 2198 4008 2202 4012
rect 2230 4018 2234 4022
rect 2222 3978 2226 3982
rect 2198 3938 2202 3942
rect 2286 4248 2290 4252
rect 2342 4248 2346 4252
rect 2302 4238 2306 4242
rect 2358 4208 2362 4212
rect 2414 4208 2418 4212
rect 2358 4198 2362 4202
rect 2270 4188 2274 4192
rect 2398 4178 2402 4182
rect 2262 4168 2266 4172
rect 2310 4168 2314 4172
rect 2286 4158 2290 4162
rect 2318 4158 2322 4162
rect 2270 4148 2274 4152
rect 2278 4148 2282 4152
rect 2246 4078 2250 4082
rect 2262 4118 2266 4122
rect 2270 4108 2274 4112
rect 2302 4148 2306 4152
rect 2438 4288 2442 4292
rect 2438 4158 2442 4162
rect 2334 4148 2338 4152
rect 2366 4148 2370 4152
rect 2414 4148 2418 4152
rect 2438 4148 2442 4152
rect 2326 4138 2330 4142
rect 2294 4128 2298 4132
rect 2390 4138 2394 4142
rect 2454 4168 2458 4172
rect 2366 4128 2370 4132
rect 2446 4128 2450 4132
rect 2438 4118 2442 4122
rect 2342 4108 2346 4112
rect 2294 4098 2298 4102
rect 2302 4098 2306 4102
rect 2310 4088 2314 4092
rect 2278 4058 2282 4062
rect 2302 4058 2306 4062
rect 2270 4028 2274 4032
rect 2302 3988 2306 3992
rect 2254 3978 2258 3982
rect 2270 3958 2274 3962
rect 2302 3958 2306 3962
rect 2286 3938 2290 3942
rect 2254 3928 2258 3932
rect 2262 3898 2266 3902
rect 2286 3898 2290 3902
rect 2238 3878 2242 3882
rect 2198 3868 2202 3872
rect 2246 3868 2250 3872
rect 2166 3798 2170 3802
rect 2190 3798 2194 3802
rect 2254 3808 2258 3812
rect 2246 3768 2250 3772
rect 2174 3758 2178 3762
rect 2206 3758 2210 3762
rect 2270 3768 2274 3772
rect 1982 3748 1986 3752
rect 2118 3748 2122 3752
rect 2134 3748 2138 3752
rect 2214 3748 2218 3752
rect 2230 3748 2234 3752
rect 2262 3748 2266 3752
rect 2030 3728 2034 3732
rect 2054 3728 2058 3732
rect 1926 3668 1930 3672
rect 1934 3658 1938 3662
rect 1918 3618 1922 3622
rect 1950 3648 1954 3652
rect 1942 3608 1946 3612
rect 1894 3598 1898 3602
rect 2262 3728 2266 3732
rect 2030 3718 2034 3722
rect 2206 3718 2210 3722
rect 2230 3718 2234 3722
rect 2278 3718 2282 3722
rect 2030 3678 2034 3682
rect 1982 3668 1986 3672
rect 2006 3668 2010 3672
rect 1974 3648 1978 3652
rect 1998 3648 2002 3652
rect 1974 3628 1978 3632
rect 1926 3588 1930 3592
rect 1958 3588 1962 3592
rect 1966 3588 1970 3592
rect 1870 3568 1874 3572
rect 1838 3528 1842 3532
rect 1902 3558 1906 3562
rect 1966 3568 1970 3572
rect 1982 3558 1986 3562
rect 1998 3558 2002 3562
rect 1926 3548 1930 3552
rect 1958 3548 1962 3552
rect 1862 3528 1866 3532
rect 1854 3508 1858 3512
rect 1886 3488 1890 3492
rect 1958 3528 1962 3532
rect 1966 3528 1970 3532
rect 1974 3518 1978 3522
rect 1998 3518 2002 3522
rect 1950 3488 1954 3492
rect 1990 3468 1994 3472
rect 1934 3458 1938 3462
rect 1982 3458 1986 3462
rect 1998 3458 2002 3462
rect 1838 3448 1842 3452
rect 1878 3448 1882 3452
rect 1886 3448 1890 3452
rect 1838 3418 1842 3422
rect 1782 3378 1786 3382
rect 1782 3358 1786 3362
rect 1742 3338 1746 3342
rect 1750 3338 1754 3342
rect 1766 3328 1770 3332
rect 1726 3308 1730 3312
rect 1726 3258 1730 3262
rect 1766 3308 1770 3312
rect 1758 3268 1762 3272
rect 1742 3248 1746 3252
rect 1702 3198 1706 3202
rect 1670 3158 1674 3162
rect 1734 3158 1738 3162
rect 1622 3148 1626 3152
rect 1670 3148 1674 3152
rect 1694 3148 1698 3152
rect 1726 3148 1730 3152
rect 1686 3138 1690 3142
rect 1638 3088 1642 3092
rect 1654 3088 1658 3092
rect 1622 3078 1626 3082
rect 1630 3078 1634 3082
rect 1654 3078 1658 3082
rect 1590 3048 1594 3052
rect 1562 3003 1566 3007
rect 1569 3003 1573 3007
rect 1662 3068 1666 3072
rect 1670 3058 1674 3062
rect 1646 3048 1650 3052
rect 1726 3108 1730 3112
rect 1710 3078 1714 3082
rect 1694 3068 1698 3072
rect 1622 3028 1626 3032
rect 1662 3028 1666 3032
rect 1606 3018 1610 3022
rect 1598 2998 1602 3002
rect 1550 2978 1554 2982
rect 1590 2968 1594 2972
rect 1478 2948 1482 2952
rect 1542 2948 1546 2952
rect 1718 3048 1722 3052
rect 1734 3048 1738 3052
rect 1710 3028 1714 3032
rect 1702 3008 1706 3012
rect 1662 2968 1666 2972
rect 1686 2958 1690 2962
rect 1622 2948 1626 2952
rect 1638 2948 1642 2952
rect 1702 2948 1706 2952
rect 1734 2948 1738 2952
rect 1750 3128 1754 3132
rect 1750 3078 1754 3082
rect 1470 2888 1474 2892
rect 1486 2878 1490 2882
rect 1694 2938 1698 2942
rect 1710 2938 1714 2942
rect 1726 2938 1730 2942
rect 1678 2918 1682 2922
rect 1598 2908 1602 2912
rect 1630 2908 1634 2912
rect 1542 2888 1546 2892
rect 1550 2888 1554 2892
rect 1534 2878 1538 2882
rect 1502 2868 1506 2872
rect 1518 2868 1522 2872
rect 1582 2868 1586 2872
rect 1670 2888 1674 2892
rect 1622 2878 1626 2882
rect 1638 2868 1642 2872
rect 1646 2868 1650 2872
rect 1582 2858 1586 2862
rect 1470 2848 1474 2852
rect 1494 2848 1498 2852
rect 1510 2848 1514 2852
rect 1534 2848 1538 2852
rect 1502 2838 1506 2842
rect 1518 2828 1522 2832
rect 1502 2798 1506 2802
rect 1470 2758 1474 2762
rect 1494 2758 1498 2762
rect 1454 2738 1458 2742
rect 1470 2738 1474 2742
rect 1486 2738 1490 2742
rect 1438 2708 1442 2712
rect 1430 2698 1434 2702
rect 1406 2668 1410 2672
rect 1414 2668 1418 2672
rect 1406 2658 1410 2662
rect 1374 2648 1378 2652
rect 1390 2648 1394 2652
rect 1390 2608 1394 2612
rect 1374 2558 1378 2562
rect 1382 2558 1386 2562
rect 1366 2528 1370 2532
rect 1358 2498 1362 2502
rect 1430 2648 1434 2652
rect 1422 2598 1426 2602
rect 1414 2538 1418 2542
rect 1390 2528 1394 2532
rect 1358 2488 1362 2492
rect 1406 2488 1410 2492
rect 1494 2698 1498 2702
rect 1446 2668 1450 2672
rect 1502 2668 1506 2672
rect 1470 2658 1474 2662
rect 1478 2648 1482 2652
rect 1470 2628 1474 2632
rect 1438 2618 1442 2622
rect 1446 2598 1450 2602
rect 1430 2548 1434 2552
rect 1454 2538 1458 2542
rect 1462 2538 1466 2542
rect 1558 2848 1562 2852
rect 1550 2808 1554 2812
rect 1562 2803 1566 2807
rect 1569 2803 1573 2807
rect 1574 2748 1578 2752
rect 1534 2718 1538 2722
rect 1550 2678 1554 2682
rect 1526 2648 1530 2652
rect 1494 2558 1498 2562
rect 1510 2558 1514 2562
rect 1478 2548 1482 2552
rect 1494 2548 1498 2552
rect 1478 2538 1482 2542
rect 1502 2538 1506 2542
rect 1470 2528 1474 2532
rect 1430 2498 1434 2502
rect 1494 2528 1498 2532
rect 1470 2488 1474 2492
rect 1478 2488 1482 2492
rect 1510 2498 1514 2502
rect 1526 2488 1530 2492
rect 1502 2458 1506 2462
rect 1470 2448 1474 2452
rect 1542 2498 1546 2502
rect 1598 2848 1602 2852
rect 1742 2888 1746 2892
rect 1750 2868 1754 2872
rect 1686 2848 1690 2852
rect 1710 2848 1714 2852
rect 1734 2848 1738 2852
rect 1678 2838 1682 2842
rect 1686 2828 1690 2832
rect 1718 2828 1722 2832
rect 1614 2798 1618 2802
rect 1726 2798 1730 2802
rect 1590 2758 1594 2762
rect 1662 2758 1666 2762
rect 1638 2748 1642 2752
rect 1670 2748 1674 2752
rect 1710 2738 1714 2742
rect 1630 2728 1634 2732
rect 1710 2728 1714 2732
rect 1718 2688 1722 2692
rect 1678 2668 1682 2672
rect 1694 2668 1698 2672
rect 1710 2668 1714 2672
rect 1566 2618 1570 2622
rect 1582 2618 1586 2622
rect 1662 2608 1666 2612
rect 1562 2603 1566 2607
rect 1569 2603 1573 2607
rect 1598 2598 1602 2602
rect 1734 2788 1738 2792
rect 1750 2828 1754 2832
rect 1742 2768 1746 2772
rect 1750 2758 1754 2762
rect 1734 2738 1738 2742
rect 1774 3238 1778 3242
rect 1766 3188 1770 3192
rect 1766 3148 1770 3152
rect 1830 3378 1834 3382
rect 1830 3368 1834 3372
rect 1806 3348 1810 3352
rect 1814 3308 1818 3312
rect 1822 3308 1826 3312
rect 1798 3268 1802 3272
rect 1798 3258 1802 3262
rect 1806 3248 1810 3252
rect 1782 3098 1786 3102
rect 1806 3078 1810 3082
rect 1766 3048 1770 3052
rect 1766 3038 1770 3042
rect 1838 3248 1842 3252
rect 1918 3408 1922 3412
rect 1942 3438 1946 3442
rect 1870 3348 1874 3352
rect 1902 3348 1906 3352
rect 1934 3338 1938 3342
rect 1910 3268 1914 3272
rect 1862 3158 1866 3162
rect 1886 3148 1890 3152
rect 1846 3128 1850 3132
rect 1830 3118 1834 3122
rect 1902 3138 1906 3142
rect 1910 3118 1914 3122
rect 1862 3098 1866 3102
rect 1830 3078 1834 3082
rect 1846 3078 1850 3082
rect 1870 3068 1874 3072
rect 1878 3068 1882 3072
rect 1998 3418 2002 3422
rect 1974 3398 1978 3402
rect 1950 3368 1954 3372
rect 2038 3648 2042 3652
rect 2198 3708 2202 3712
rect 2074 3703 2078 3707
rect 2081 3703 2085 3707
rect 2134 3698 2138 3702
rect 2150 3678 2154 3682
rect 2166 3668 2170 3672
rect 2110 3659 2114 3663
rect 2158 3648 2162 3652
rect 2190 3648 2194 3652
rect 2166 3618 2170 3622
rect 2126 3608 2130 3612
rect 2110 3568 2114 3572
rect 2030 3548 2034 3552
rect 2046 3548 2050 3552
rect 2062 3548 2066 3552
rect 2030 3518 2034 3522
rect 2014 3508 2018 3512
rect 2094 3518 2098 3522
rect 2074 3503 2078 3507
rect 2081 3503 2085 3507
rect 2038 3488 2042 3492
rect 2062 3488 2066 3492
rect 2142 3558 2146 3562
rect 2174 3568 2178 3572
rect 2190 3558 2194 3562
rect 2158 3548 2162 3552
rect 2014 3468 2018 3472
rect 2022 3468 2026 3472
rect 2062 3468 2066 3472
rect 2086 3468 2090 3472
rect 2014 3438 2018 3442
rect 2006 3358 2010 3362
rect 2046 3458 2050 3462
rect 2038 3448 2042 3452
rect 2030 3438 2034 3442
rect 2038 3378 2042 3382
rect 2006 3348 2010 3352
rect 2054 3448 2058 3452
rect 2078 3448 2082 3452
rect 2062 3438 2066 3442
rect 2110 3448 2114 3452
rect 2142 3448 2146 3452
rect 2134 3438 2138 3442
rect 2094 3428 2098 3432
rect 2062 3358 2066 3362
rect 1958 3278 1962 3282
rect 1958 3258 1962 3262
rect 1950 3248 1954 3252
rect 1958 3248 1962 3252
rect 2014 3338 2018 3342
rect 2030 3338 2034 3342
rect 2038 3298 2042 3302
rect 2038 3278 2042 3282
rect 2070 3338 2074 3342
rect 2102 3338 2106 3342
rect 2062 3308 2066 3312
rect 2014 3268 2018 3272
rect 2074 3303 2078 3307
rect 2081 3303 2085 3307
rect 2078 3268 2082 3272
rect 2070 3258 2074 3262
rect 1982 3218 1986 3222
rect 1974 3208 1978 3212
rect 1966 3158 1970 3162
rect 1958 3148 1962 3152
rect 1934 3138 1938 3142
rect 1942 3118 1946 3122
rect 1974 3118 1978 3122
rect 1966 3108 1970 3112
rect 1958 3088 1962 3092
rect 1910 3068 1914 3072
rect 1838 3048 1842 3052
rect 1790 3028 1794 3032
rect 1822 3028 1826 3032
rect 1774 2998 1778 3002
rect 1782 2998 1786 3002
rect 1766 2978 1770 2982
rect 1774 2968 1778 2972
rect 1870 3028 1874 3032
rect 1854 3018 1858 3022
rect 1798 2988 1802 2992
rect 1822 2988 1826 2992
rect 1878 2978 1882 2982
rect 1822 2958 1826 2962
rect 1838 2958 1842 2962
rect 1846 2958 1850 2962
rect 1806 2948 1810 2952
rect 1822 2948 1826 2952
rect 1782 2938 1786 2942
rect 1782 2888 1786 2892
rect 1766 2738 1770 2742
rect 1750 2728 1754 2732
rect 1758 2728 1762 2732
rect 1742 2678 1746 2682
rect 1726 2668 1730 2672
rect 1750 2668 1754 2672
rect 1822 2928 1826 2932
rect 1830 2928 1834 2932
rect 1838 2888 1842 2892
rect 1790 2868 1794 2872
rect 1854 2868 1858 2872
rect 1846 2848 1850 2852
rect 1878 2848 1882 2852
rect 1870 2828 1874 2832
rect 1798 2788 1802 2792
rect 1790 2778 1794 2782
rect 1790 2768 1794 2772
rect 1918 3058 1922 3062
rect 1926 3058 1930 3062
rect 1942 3058 1946 3062
rect 1942 3038 1946 3042
rect 1934 3008 1938 3012
rect 1918 2988 1922 2992
rect 1910 2928 1914 2932
rect 1926 2898 1930 2902
rect 1894 2868 1898 2872
rect 1942 2958 1946 2962
rect 1934 2888 1938 2892
rect 2014 3148 2018 3152
rect 2014 3128 2018 3132
rect 1998 3048 2002 3052
rect 2094 3238 2098 3242
rect 2078 3158 2082 3162
rect 2094 3138 2098 3142
rect 2062 3118 2066 3122
rect 2074 3103 2078 3107
rect 2081 3103 2085 3107
rect 2070 3078 2074 3082
rect 2038 3058 2042 3062
rect 2078 3058 2082 3062
rect 2014 3048 2018 3052
rect 2046 3038 2050 3042
rect 2054 3038 2058 3042
rect 2006 3028 2010 3032
rect 2118 3308 2122 3312
rect 2134 3308 2138 3312
rect 2262 3698 2266 3702
rect 2230 3598 2234 3602
rect 2230 3548 2234 3552
rect 2278 3668 2282 3672
rect 2318 4058 2322 4062
rect 2334 4028 2338 4032
rect 2446 4068 2450 4072
rect 2398 4058 2402 4062
rect 2430 4058 2434 4062
rect 2358 4048 2362 4052
rect 2510 4338 2514 4342
rect 2542 4338 2546 4342
rect 2630 4338 2634 4342
rect 2566 4328 2570 4332
rect 2558 4318 2562 4322
rect 2494 4278 2498 4282
rect 2494 4238 2498 4242
rect 2518 4238 2522 4242
rect 2542 4238 2546 4242
rect 2526 4198 2530 4202
rect 2486 4178 2490 4182
rect 2478 4168 2482 4172
rect 2470 4158 2474 4162
rect 2478 4148 2482 4152
rect 2470 4108 2474 4112
rect 2350 4038 2354 4042
rect 2462 4038 2466 4042
rect 2342 4018 2346 4022
rect 2374 3998 2378 4002
rect 2342 3968 2346 3972
rect 2350 3968 2354 3972
rect 2390 3968 2394 3972
rect 2414 3968 2418 3972
rect 2374 3938 2378 3942
rect 2366 3928 2370 3932
rect 2318 3918 2322 3922
rect 2342 3878 2346 3882
rect 2334 3868 2338 3872
rect 2302 3858 2306 3862
rect 2374 3858 2378 3862
rect 2310 3818 2314 3822
rect 2326 3848 2330 3852
rect 2358 3848 2362 3852
rect 2342 3838 2346 3842
rect 2318 3808 2322 3812
rect 2318 3698 2322 3702
rect 2310 3668 2314 3672
rect 2334 3668 2338 3672
rect 2326 3658 2330 3662
rect 2334 3638 2338 3642
rect 2294 3598 2298 3602
rect 2406 3918 2410 3922
rect 2462 3978 2466 3982
rect 2430 3928 2434 3932
rect 2502 4118 2506 4122
rect 2518 4088 2522 4092
rect 2534 4158 2538 4162
rect 2678 4318 2682 4322
rect 2686 4318 2690 4322
rect 2662 4288 2666 4292
rect 2662 4258 2666 4262
rect 2702 4298 2706 4302
rect 2686 4288 2690 4292
rect 2718 4308 2722 4312
rect 2734 4308 2738 4312
rect 2718 4288 2722 4292
rect 2702 4268 2706 4272
rect 2750 4428 2754 4432
rect 2782 4438 2786 4442
rect 2766 4428 2770 4432
rect 2758 4418 2762 4422
rect 2750 4408 2754 4412
rect 2798 4438 2802 4442
rect 2790 4418 2794 4422
rect 2942 4558 2946 4562
rect 2990 4628 2994 4632
rect 3014 4618 3018 4622
rect 3022 4568 3026 4572
rect 2982 4558 2986 4562
rect 3022 4558 3026 4562
rect 3030 4558 3034 4562
rect 2990 4548 2994 4552
rect 3022 4548 3026 4552
rect 2982 4538 2986 4542
rect 2966 4528 2970 4532
rect 2910 4518 2914 4522
rect 2838 4488 2842 4492
rect 2806 4388 2810 4392
rect 2790 4368 2794 4372
rect 2782 4348 2786 4352
rect 2790 4348 2794 4352
rect 2710 4258 2714 4262
rect 2726 4258 2730 4262
rect 2742 4258 2746 4262
rect 2598 4228 2602 4232
rect 2586 4203 2590 4207
rect 2593 4203 2597 4207
rect 2574 4158 2578 4162
rect 2622 4158 2626 4162
rect 2670 4158 2674 4162
rect 2678 4158 2682 4162
rect 2614 4138 2618 4142
rect 2566 4098 2570 4102
rect 2542 4068 2546 4072
rect 2438 3918 2442 3922
rect 2422 3908 2426 3912
rect 2422 3878 2426 3882
rect 2470 3918 2474 3922
rect 2414 3858 2418 3862
rect 2438 3858 2442 3862
rect 2406 3848 2410 3852
rect 2446 3828 2450 3832
rect 2398 3818 2402 3822
rect 2382 3808 2386 3812
rect 2382 3788 2386 3792
rect 2350 3768 2354 3772
rect 2390 3778 2394 3782
rect 2382 3748 2386 3752
rect 2414 3748 2418 3752
rect 2422 3738 2426 3742
rect 2366 3728 2370 3732
rect 2526 4018 2530 4022
rect 2542 4018 2546 4022
rect 2486 3958 2490 3962
rect 2558 4008 2562 4012
rect 2542 3988 2546 3992
rect 2510 3928 2514 3932
rect 2518 3898 2522 3902
rect 2486 3878 2490 3882
rect 2510 3878 2514 3882
rect 2534 3878 2538 3882
rect 2606 4128 2610 4132
rect 2670 4128 2674 4132
rect 2654 4108 2658 4112
rect 2614 4098 2618 4102
rect 2582 4068 2586 4072
rect 2654 4068 2658 4072
rect 2590 4038 2594 4042
rect 2586 4003 2590 4007
rect 2593 4003 2597 4007
rect 2598 3978 2602 3982
rect 2574 3938 2578 3942
rect 2598 3938 2602 3942
rect 2702 4208 2706 4212
rect 2726 4238 2730 4242
rect 2726 4228 2730 4232
rect 2750 4228 2754 4232
rect 2750 4168 2754 4172
rect 2710 4148 2714 4152
rect 2718 4148 2722 4152
rect 2750 4148 2754 4152
rect 2694 4128 2698 4132
rect 2822 4398 2826 4402
rect 2846 4388 2850 4392
rect 2814 4368 2818 4372
rect 2814 4348 2818 4352
rect 2830 4338 2834 4342
rect 2854 4288 2858 4292
rect 2838 4268 2842 4272
rect 2782 4248 2786 4252
rect 2806 4228 2810 4232
rect 2782 4208 2786 4212
rect 2790 4148 2794 4152
rect 2710 4128 2714 4132
rect 2766 4128 2770 4132
rect 2774 4128 2778 4132
rect 2686 4118 2690 4122
rect 2702 4118 2706 4122
rect 2774 4098 2778 4102
rect 2758 4088 2762 4092
rect 2678 4058 2682 4062
rect 2638 4048 2642 4052
rect 2622 4038 2626 4042
rect 2614 4018 2618 4022
rect 2606 3928 2610 3932
rect 2558 3898 2562 3902
rect 2566 3848 2570 3852
rect 2542 3818 2546 3822
rect 2534 3798 2538 3802
rect 2518 3758 2522 3762
rect 2446 3748 2450 3752
rect 2462 3748 2466 3752
rect 2478 3748 2482 3752
rect 2486 3748 2490 3752
rect 2382 3718 2386 3722
rect 2398 3718 2402 3722
rect 2438 3718 2442 3722
rect 2374 3698 2378 3702
rect 2398 3678 2402 3682
rect 2358 3668 2362 3672
rect 2366 3648 2370 3652
rect 2326 3588 2330 3592
rect 2342 3588 2346 3592
rect 2310 3568 2314 3572
rect 2286 3548 2290 3552
rect 2190 3538 2194 3542
rect 2214 3538 2218 3542
rect 2230 3538 2234 3542
rect 2174 3528 2178 3532
rect 2166 3518 2170 3522
rect 2158 3498 2162 3502
rect 2166 3488 2170 3492
rect 2158 3458 2162 3462
rect 2174 3448 2178 3452
rect 2158 3398 2162 3402
rect 2158 3368 2162 3372
rect 2222 3458 2226 3462
rect 2206 3368 2210 3372
rect 2190 3358 2194 3362
rect 2214 3358 2218 3362
rect 2174 3348 2178 3352
rect 2198 3338 2202 3342
rect 2214 3338 2218 3342
rect 2214 3308 2218 3312
rect 2166 3298 2170 3302
rect 2134 3268 2138 3272
rect 2182 3258 2186 3262
rect 2134 3248 2138 3252
rect 2150 3238 2154 3242
rect 2158 3188 2162 3192
rect 2126 3168 2130 3172
rect 2150 3168 2154 3172
rect 2110 3158 2114 3162
rect 2134 3148 2138 3152
rect 2278 3498 2282 3502
rect 2478 3718 2482 3722
rect 2462 3668 2466 3672
rect 2446 3658 2450 3662
rect 2454 3638 2458 3642
rect 2398 3608 2402 3612
rect 2382 3588 2386 3592
rect 2398 3568 2402 3572
rect 2422 3568 2426 3572
rect 2462 3568 2466 3572
rect 2334 3548 2338 3552
rect 2374 3548 2378 3552
rect 2390 3548 2394 3552
rect 2366 3538 2370 3542
rect 2414 3538 2418 3542
rect 2374 3518 2378 3522
rect 2350 3488 2354 3492
rect 2446 3548 2450 3552
rect 2470 3538 2474 3542
rect 2518 3738 2522 3742
rect 2502 3728 2506 3732
rect 2518 3668 2522 3672
rect 2550 3778 2554 3782
rect 2590 3858 2594 3862
rect 2638 4008 2642 4012
rect 2638 3988 2642 3992
rect 2630 3958 2634 3962
rect 2758 4058 2762 4062
rect 2678 4048 2682 4052
rect 2742 4048 2746 4052
rect 2686 4018 2690 4022
rect 2702 4018 2706 4022
rect 2718 4018 2722 4022
rect 2654 3988 2658 3992
rect 2694 3988 2698 3992
rect 2662 3968 2666 3972
rect 2670 3948 2674 3952
rect 2646 3938 2650 3942
rect 2630 3918 2634 3922
rect 2654 3918 2658 3922
rect 2614 3878 2618 3882
rect 2622 3878 2626 3882
rect 2630 3868 2634 3872
rect 2646 3868 2650 3872
rect 2606 3838 2610 3842
rect 2586 3803 2590 3807
rect 2593 3803 2597 3807
rect 2630 3808 2634 3812
rect 2630 3798 2634 3802
rect 2606 3788 2610 3792
rect 2574 3758 2578 3762
rect 2598 3758 2602 3762
rect 2574 3738 2578 3742
rect 2614 3738 2618 3742
rect 2566 3698 2570 3702
rect 2550 3688 2554 3692
rect 2542 3668 2546 3672
rect 2574 3678 2578 3682
rect 2526 3658 2530 3662
rect 2494 3618 2498 3622
rect 2486 3528 2490 3532
rect 2430 3518 2434 3522
rect 2478 3508 2482 3512
rect 2446 3498 2450 3502
rect 2334 3468 2338 3472
rect 2302 3458 2306 3462
rect 2398 3459 2402 3463
rect 2270 3448 2274 3452
rect 2318 3448 2322 3452
rect 2286 3438 2290 3442
rect 2230 3348 2234 3352
rect 2230 3308 2234 3312
rect 2238 3298 2242 3302
rect 2238 3278 2242 3282
rect 2222 3178 2226 3182
rect 2214 3158 2218 3162
rect 2270 3358 2274 3362
rect 2302 3358 2306 3362
rect 2262 3338 2266 3342
rect 2286 3338 2290 3342
rect 2278 3328 2282 3332
rect 2278 3288 2282 3292
rect 2470 3488 2474 3492
rect 2454 3468 2458 3472
rect 2446 3448 2450 3452
rect 2438 3438 2442 3442
rect 2446 3418 2450 3422
rect 2422 3368 2426 3372
rect 2334 3358 2338 3362
rect 2366 3358 2370 3362
rect 2334 3348 2338 3352
rect 2350 3348 2354 3352
rect 2326 3288 2330 3292
rect 2310 3278 2314 3282
rect 2318 3278 2322 3282
rect 2286 3268 2290 3272
rect 2310 3258 2314 3262
rect 2326 3248 2330 3252
rect 2294 3238 2298 3242
rect 2278 3208 2282 3212
rect 2270 3198 2274 3202
rect 2174 3148 2178 3152
rect 2206 3148 2210 3152
rect 2246 3148 2250 3152
rect 2190 3138 2194 3142
rect 2254 3138 2258 3142
rect 2126 3118 2130 3122
rect 2182 3118 2186 3122
rect 2102 3078 2106 3082
rect 2134 3068 2138 3072
rect 2158 3068 2162 3072
rect 2270 3068 2274 3072
rect 2062 3018 2066 3022
rect 1990 3008 1994 3012
rect 2022 2988 2026 2992
rect 2014 2978 2018 2982
rect 2038 2978 2042 2982
rect 2006 2968 2010 2972
rect 2102 2958 2106 2962
rect 2030 2948 2034 2952
rect 2070 2948 2074 2952
rect 1998 2938 2002 2942
rect 1958 2898 1962 2902
rect 1998 2928 2002 2932
rect 2014 2928 2018 2932
rect 2074 2903 2078 2907
rect 2081 2903 2085 2907
rect 2022 2898 2026 2902
rect 1958 2888 1962 2892
rect 1966 2888 1970 2892
rect 1942 2868 1946 2872
rect 1902 2848 1906 2852
rect 1910 2848 1914 2852
rect 1966 2798 1970 2802
rect 1886 2788 1890 2792
rect 1950 2778 1954 2782
rect 1854 2758 1858 2762
rect 1862 2758 1866 2762
rect 1870 2758 1874 2762
rect 1838 2748 1842 2752
rect 1790 2738 1794 2742
rect 1774 2658 1778 2662
rect 1726 2648 1730 2652
rect 1734 2648 1738 2652
rect 1766 2628 1770 2632
rect 1734 2608 1738 2612
rect 1702 2598 1706 2602
rect 1686 2578 1690 2582
rect 1686 2568 1690 2572
rect 1670 2558 1674 2562
rect 1702 2558 1706 2562
rect 1574 2548 1578 2552
rect 1662 2548 1666 2552
rect 1742 2538 1746 2542
rect 1574 2508 1578 2512
rect 1654 2508 1658 2512
rect 1598 2488 1602 2492
rect 1550 2478 1554 2482
rect 1582 2478 1586 2482
rect 1654 2478 1658 2482
rect 1550 2458 1554 2462
rect 1422 2428 1426 2432
rect 1406 2388 1410 2392
rect 1366 2378 1370 2382
rect 1382 2378 1386 2382
rect 1358 2368 1362 2372
rect 1326 2348 1330 2352
rect 1350 2348 1354 2352
rect 1262 2338 1266 2342
rect 1294 2338 1298 2342
rect 1302 2338 1306 2342
rect 1262 2278 1266 2282
rect 1350 2338 1354 2342
rect 1342 2278 1346 2282
rect 1398 2368 1402 2372
rect 1454 2368 1458 2372
rect 1446 2348 1450 2352
rect 1390 2338 1394 2342
rect 1430 2328 1434 2332
rect 1374 2308 1378 2312
rect 1430 2308 1434 2312
rect 1286 2268 1290 2272
rect 1310 2258 1314 2262
rect 1278 2248 1282 2252
rect 1294 2238 1298 2242
rect 1302 2238 1306 2242
rect 1294 2228 1298 2232
rect 1286 2178 1290 2182
rect 1278 2158 1282 2162
rect 1318 2218 1322 2222
rect 1318 2148 1322 2152
rect 1294 2138 1298 2142
rect 1270 2128 1274 2132
rect 1374 2258 1378 2262
rect 1334 2238 1338 2242
rect 1350 2188 1354 2192
rect 1366 2178 1370 2182
rect 1350 2168 1354 2172
rect 1358 2168 1362 2172
rect 1366 2158 1370 2162
rect 1302 2118 1306 2122
rect 1326 2118 1330 2122
rect 1230 2088 1234 2092
rect 1238 2088 1242 2092
rect 1246 2088 1250 2092
rect 1214 2078 1218 2082
rect 1150 2058 1154 2062
rect 1206 2038 1210 2042
rect 1190 2028 1194 2032
rect 1182 2008 1186 2012
rect 1158 1958 1162 1962
rect 1070 1948 1074 1952
rect 1094 1948 1098 1952
rect 1206 1948 1210 1952
rect 1062 1938 1066 1942
rect 1030 1898 1034 1902
rect 1022 1878 1026 1882
rect 982 1868 986 1872
rect 1014 1858 1018 1862
rect 1050 1903 1054 1907
rect 1057 1903 1061 1907
rect 1062 1888 1066 1892
rect 998 1848 1002 1852
rect 1038 1848 1042 1852
rect 958 1818 962 1822
rect 958 1738 962 1742
rect 958 1718 962 1722
rect 950 1708 954 1712
rect 982 1728 986 1732
rect 982 1698 986 1702
rect 942 1688 946 1692
rect 926 1678 930 1682
rect 926 1668 930 1672
rect 966 1678 970 1682
rect 918 1658 922 1662
rect 1142 1938 1146 1942
rect 1094 1918 1098 1922
rect 1150 1878 1154 1882
rect 1166 1938 1170 1942
rect 1174 1938 1178 1942
rect 1190 1938 1194 1942
rect 1086 1858 1090 1862
rect 1078 1848 1082 1852
rect 1086 1818 1090 1822
rect 1022 1738 1026 1742
rect 1126 1848 1130 1852
rect 1134 1828 1138 1832
rect 1102 1818 1106 1822
rect 1118 1808 1122 1812
rect 1118 1788 1122 1792
rect 1102 1738 1106 1742
rect 1118 1738 1122 1742
rect 1030 1728 1034 1732
rect 1086 1728 1090 1732
rect 1094 1728 1098 1732
rect 1050 1703 1054 1707
rect 1057 1703 1061 1707
rect 1054 1688 1058 1692
rect 1118 1728 1122 1732
rect 1110 1708 1114 1712
rect 1022 1668 1026 1672
rect 1046 1668 1050 1672
rect 1102 1668 1106 1672
rect 982 1658 986 1662
rect 1006 1658 1010 1662
rect 1038 1658 1042 1662
rect 862 1648 866 1652
rect 934 1648 938 1652
rect 950 1648 954 1652
rect 870 1568 874 1572
rect 926 1558 930 1562
rect 878 1548 882 1552
rect 894 1548 898 1552
rect 918 1548 922 1552
rect 838 1538 842 1542
rect 886 1538 890 1542
rect 790 1528 794 1532
rect 878 1478 882 1482
rect 718 1468 722 1472
rect 750 1468 754 1472
rect 774 1468 778 1472
rect 790 1458 794 1462
rect 806 1458 810 1462
rect 854 1459 858 1463
rect 742 1418 746 1422
rect 734 1388 738 1392
rect 758 1388 762 1392
rect 726 1348 730 1352
rect 774 1348 778 1352
rect 878 1448 882 1452
rect 798 1428 802 1432
rect 830 1418 834 1422
rect 902 1418 906 1422
rect 854 1398 858 1402
rect 846 1368 850 1372
rect 806 1358 810 1362
rect 830 1358 834 1362
rect 870 1358 874 1362
rect 902 1358 906 1362
rect 998 1648 1002 1652
rect 1006 1648 1010 1652
rect 1006 1558 1010 1562
rect 1022 1578 1026 1582
rect 1046 1648 1050 1652
rect 1110 1648 1114 1652
rect 1110 1628 1114 1632
rect 1070 1578 1074 1582
rect 1038 1568 1042 1572
rect 1022 1558 1026 1562
rect 950 1548 954 1552
rect 998 1548 1002 1552
rect 1046 1548 1050 1552
rect 958 1538 962 1542
rect 974 1538 978 1542
rect 1030 1538 1034 1542
rect 1014 1518 1018 1522
rect 966 1508 970 1512
rect 934 1498 938 1502
rect 1050 1503 1054 1507
rect 1057 1503 1061 1507
rect 942 1458 946 1462
rect 958 1458 962 1462
rect 1014 1458 1018 1462
rect 1078 1548 1082 1552
rect 1134 1678 1138 1682
rect 1182 1888 1186 1892
rect 1230 2068 1234 2072
rect 1238 2048 1242 2052
rect 1230 2028 1234 2032
rect 1230 1908 1234 1912
rect 1206 1868 1210 1872
rect 1214 1868 1218 1872
rect 1222 1868 1226 1872
rect 1198 1858 1202 1862
rect 1270 2088 1274 2092
rect 1294 2068 1298 2072
rect 1310 2078 1314 2082
rect 1270 2058 1274 2062
rect 1286 2058 1290 2062
rect 1270 2048 1274 2052
rect 1310 2038 1314 2042
rect 1318 2038 1322 2042
rect 1286 1958 1290 1962
rect 1294 1958 1298 1962
rect 1310 1958 1314 1962
rect 1302 1948 1306 1952
rect 1278 1938 1282 1942
rect 1294 1938 1298 1942
rect 1278 1908 1282 1912
rect 1230 1858 1234 1862
rect 1230 1848 1234 1852
rect 1254 1848 1258 1852
rect 1238 1838 1242 1842
rect 1214 1808 1218 1812
rect 1246 1808 1250 1812
rect 1238 1798 1242 1802
rect 1214 1788 1218 1792
rect 1158 1758 1162 1762
rect 1278 1818 1282 1822
rect 1262 1778 1266 1782
rect 1174 1748 1178 1752
rect 1254 1748 1258 1752
rect 1206 1738 1210 1742
rect 1214 1738 1218 1742
rect 1198 1698 1202 1702
rect 1190 1688 1194 1692
rect 1206 1688 1210 1692
rect 1166 1678 1170 1682
rect 1182 1658 1186 1662
rect 1174 1638 1178 1642
rect 1126 1558 1130 1562
rect 1174 1628 1178 1632
rect 1262 1738 1266 1742
rect 1286 1748 1290 1752
rect 1286 1738 1290 1742
rect 1246 1688 1250 1692
rect 1238 1668 1242 1672
rect 1278 1728 1282 1732
rect 1286 1728 1290 1732
rect 1270 1718 1274 1722
rect 1262 1708 1266 1712
rect 1406 2248 1410 2252
rect 1422 2198 1426 2202
rect 1398 2168 1402 2172
rect 1414 2168 1418 2172
rect 1398 2158 1402 2162
rect 1382 2138 1386 2142
rect 1350 2098 1354 2102
rect 1374 2098 1378 2102
rect 1342 2078 1346 2082
rect 1390 2059 1394 2063
rect 1366 2038 1370 2042
rect 1334 2018 1338 2022
rect 1350 2018 1354 2022
rect 1334 1978 1338 1982
rect 1382 1978 1386 1982
rect 1358 1958 1362 1962
rect 1382 1948 1386 1952
rect 1358 1938 1362 1942
rect 1406 2138 1410 2142
rect 1462 2238 1466 2242
rect 1438 2198 1442 2202
rect 1454 2168 1458 2172
rect 1454 2148 1458 2152
rect 1446 2138 1450 2142
rect 1446 2048 1450 2052
rect 1414 1998 1418 2002
rect 1398 1938 1402 1942
rect 1462 2078 1466 2082
rect 1430 1958 1434 1962
rect 1454 1958 1458 1962
rect 1454 1948 1458 1952
rect 1526 2418 1530 2422
rect 1518 2338 1522 2342
rect 1494 2308 1498 2312
rect 1494 2288 1498 2292
rect 1502 2288 1506 2292
rect 1502 2278 1506 2282
rect 1478 2268 1482 2272
rect 1486 2258 1490 2262
rect 1510 2268 1514 2272
rect 1562 2403 1566 2407
rect 1569 2403 1573 2407
rect 1542 2378 1546 2382
rect 1702 2528 1706 2532
rect 1678 2508 1682 2512
rect 1670 2488 1674 2492
rect 1686 2498 1690 2502
rect 1726 2508 1730 2512
rect 1742 2508 1746 2512
rect 1710 2498 1714 2502
rect 1694 2488 1698 2492
rect 1662 2468 1666 2472
rect 1678 2468 1682 2472
rect 1702 2478 1706 2482
rect 1726 2478 1730 2482
rect 1758 2488 1762 2492
rect 1758 2478 1762 2482
rect 1878 2748 1882 2752
rect 1926 2747 1930 2751
rect 1822 2738 1826 2742
rect 1886 2738 1890 2742
rect 1822 2728 1826 2732
rect 1814 2718 1818 2722
rect 1806 2678 1810 2682
rect 1854 2708 1858 2712
rect 1894 2718 1898 2722
rect 1918 2718 1922 2722
rect 1942 2708 1946 2712
rect 1894 2678 1898 2682
rect 1950 2678 1954 2682
rect 1862 2668 1866 2672
rect 1822 2648 1826 2652
rect 1830 2618 1834 2622
rect 1798 2578 1802 2582
rect 1822 2558 1826 2562
rect 1862 2588 1866 2592
rect 1838 2578 1842 2582
rect 1998 2848 2002 2852
rect 1990 2808 1994 2812
rect 1990 2758 1994 2762
rect 1990 2738 1994 2742
rect 1982 2728 1986 2732
rect 2006 2728 2010 2732
rect 2038 2888 2042 2892
rect 2070 2888 2074 2892
rect 2094 2888 2098 2892
rect 2102 2858 2106 2862
rect 2046 2848 2050 2852
rect 2046 2808 2050 2812
rect 2030 2798 2034 2802
rect 2054 2798 2058 2802
rect 2030 2768 2034 2772
rect 2030 2748 2034 2752
rect 2038 2738 2042 2742
rect 2022 2678 2026 2682
rect 2134 3048 2138 3052
rect 2126 3028 2130 3032
rect 2230 3048 2234 3052
rect 2230 3038 2234 3042
rect 2142 3008 2146 3012
rect 2182 2988 2186 2992
rect 2134 2968 2138 2972
rect 2222 2978 2226 2982
rect 2262 3058 2266 3062
rect 2270 3038 2274 3042
rect 2270 3008 2274 3012
rect 2262 2978 2266 2982
rect 2246 2968 2250 2972
rect 2166 2948 2170 2952
rect 2158 2938 2162 2942
rect 2174 2938 2178 2942
rect 2206 2938 2210 2942
rect 2238 2938 2242 2942
rect 2318 3178 2322 3182
rect 2326 3178 2330 3182
rect 2318 3168 2322 3172
rect 2366 3308 2370 3312
rect 2398 3298 2402 3302
rect 2438 3298 2442 3302
rect 2358 3268 2362 3272
rect 2374 3258 2378 3262
rect 2438 3278 2442 3282
rect 2462 3358 2466 3362
rect 2454 3328 2458 3332
rect 2518 3608 2522 3612
rect 2510 3538 2514 3542
rect 2510 3528 2514 3532
rect 2494 3448 2498 3452
rect 2502 3448 2506 3452
rect 2494 3438 2498 3442
rect 2502 3418 2506 3422
rect 2478 3288 2482 3292
rect 2494 3288 2498 3292
rect 2502 3268 2506 3272
rect 2494 3258 2498 3262
rect 2350 3228 2354 3232
rect 2430 3198 2434 3202
rect 2502 3238 2506 3242
rect 2486 3198 2490 3202
rect 2454 3188 2458 3192
rect 2366 3168 2370 3172
rect 2446 3168 2450 3172
rect 2334 3158 2338 3162
rect 2350 3158 2354 3162
rect 2446 3158 2450 3162
rect 2454 3158 2458 3162
rect 2430 3148 2434 3152
rect 2502 3148 2506 3152
rect 2342 3138 2346 3142
rect 2374 3128 2378 3132
rect 2294 3118 2298 3122
rect 2302 3118 2306 3122
rect 2286 3058 2290 3062
rect 2454 3098 2458 3102
rect 2486 3098 2490 3102
rect 2310 3078 2314 3082
rect 2350 3078 2354 3082
rect 2422 3068 2426 3072
rect 2310 3048 2314 3052
rect 2334 3008 2338 3012
rect 2278 2988 2282 2992
rect 2254 2918 2258 2922
rect 2158 2898 2162 2902
rect 2150 2888 2154 2892
rect 2126 2868 2130 2872
rect 2134 2858 2138 2862
rect 2118 2828 2122 2832
rect 2174 2838 2178 2842
rect 2150 2818 2154 2822
rect 2134 2768 2138 2772
rect 2094 2758 2098 2762
rect 2126 2758 2130 2762
rect 2086 2738 2090 2742
rect 2110 2738 2114 2742
rect 2074 2703 2078 2707
rect 2081 2703 2085 2707
rect 2078 2678 2082 2682
rect 2110 2678 2114 2682
rect 2022 2668 2026 2672
rect 2046 2668 2050 2672
rect 1934 2658 1938 2662
rect 1950 2658 1954 2662
rect 2006 2658 2010 2662
rect 2038 2658 2042 2662
rect 2102 2658 2106 2662
rect 1998 2648 2002 2652
rect 2030 2638 2034 2642
rect 1958 2628 1962 2632
rect 1934 2598 1938 2602
rect 1918 2588 1922 2592
rect 1894 2548 1898 2552
rect 1782 2538 1786 2542
rect 2022 2558 2026 2562
rect 1926 2548 1930 2552
rect 1950 2548 1954 2552
rect 1990 2548 1994 2552
rect 1998 2548 2002 2552
rect 2006 2548 2010 2552
rect 1886 2538 1890 2542
rect 1918 2538 1922 2542
rect 1942 2538 1946 2542
rect 1862 2518 1866 2522
rect 1830 2508 1834 2512
rect 1798 2488 1802 2492
rect 1814 2488 1818 2492
rect 1822 2488 1826 2492
rect 1830 2478 1834 2482
rect 1854 2478 1858 2482
rect 1758 2468 1762 2472
rect 1766 2468 1770 2472
rect 1622 2458 1626 2462
rect 1710 2458 1714 2462
rect 1734 2458 1738 2462
rect 1750 2458 1754 2462
rect 1798 2458 1802 2462
rect 1590 2438 1594 2442
rect 1702 2438 1706 2442
rect 1622 2408 1626 2412
rect 1558 2368 1562 2372
rect 1582 2368 1586 2372
rect 1606 2368 1610 2372
rect 1646 2368 1650 2372
rect 1622 2348 1626 2352
rect 1646 2348 1650 2352
rect 1574 2328 1578 2332
rect 1598 2338 1602 2342
rect 1630 2338 1634 2342
rect 1590 2308 1594 2312
rect 1622 2308 1626 2312
rect 1582 2278 1586 2282
rect 1542 2268 1546 2272
rect 1622 2268 1626 2272
rect 1502 2148 1506 2152
rect 1486 2118 1490 2122
rect 1494 2098 1498 2102
rect 1550 2248 1554 2252
rect 1598 2248 1602 2252
rect 1526 2198 1530 2202
rect 1526 2148 1530 2152
rect 1518 2138 1522 2142
rect 1562 2203 1566 2207
rect 1569 2203 1573 2207
rect 1542 2158 1546 2162
rect 1550 2118 1554 2122
rect 1574 2098 1578 2102
rect 1518 2088 1522 2092
rect 1502 2078 1506 2082
rect 1550 2078 1554 2082
rect 1598 2168 1602 2172
rect 1598 2088 1602 2092
rect 1638 2328 1642 2332
rect 1702 2388 1706 2392
rect 1702 2378 1706 2382
rect 1718 2378 1722 2382
rect 1670 2368 1674 2372
rect 1670 2348 1674 2352
rect 1686 2328 1690 2332
rect 1694 2318 1698 2322
rect 1654 2308 1658 2312
rect 1670 2298 1674 2302
rect 1710 2358 1714 2362
rect 1726 2348 1730 2352
rect 1814 2438 1818 2442
rect 1790 2348 1794 2352
rect 1694 2278 1698 2282
rect 1662 2268 1666 2272
rect 1678 2268 1682 2272
rect 1670 2248 1674 2252
rect 1662 2228 1666 2232
rect 1638 2218 1642 2222
rect 1686 2208 1690 2212
rect 1734 2298 1738 2302
rect 1718 2268 1722 2272
rect 1726 2258 1730 2262
rect 1742 2288 1746 2292
rect 1758 2298 1762 2302
rect 1750 2278 1754 2282
rect 1782 2268 1786 2272
rect 1750 2258 1754 2262
rect 1710 2248 1714 2252
rect 1702 2238 1706 2242
rect 1742 2238 1746 2242
rect 1710 2228 1714 2232
rect 1630 2168 1634 2172
rect 1662 2168 1666 2172
rect 1694 2168 1698 2172
rect 1622 2138 1626 2142
rect 1662 2108 1666 2112
rect 1670 2108 1674 2112
rect 1638 2078 1642 2082
rect 1590 2068 1594 2072
rect 1614 2068 1618 2072
rect 1742 2208 1746 2212
rect 1726 2168 1730 2172
rect 1734 2168 1738 2172
rect 1710 2138 1714 2142
rect 1702 2118 1706 2122
rect 1678 2088 1682 2092
rect 1718 2088 1722 2092
rect 1742 2138 1746 2142
rect 1726 2078 1730 2082
rect 1798 2338 1802 2342
rect 1798 2308 1802 2312
rect 1806 2298 1810 2302
rect 1862 2458 1866 2462
rect 1878 2478 1882 2482
rect 1902 2498 1906 2502
rect 1894 2488 1898 2492
rect 1942 2518 1946 2522
rect 1910 2488 1914 2492
rect 1934 2498 1938 2502
rect 1926 2478 1930 2482
rect 1910 2458 1914 2462
rect 1870 2448 1874 2452
rect 1878 2448 1882 2452
rect 1942 2448 1946 2452
rect 1846 2438 1850 2442
rect 1854 2438 1858 2442
rect 1854 2418 1858 2422
rect 1830 2388 1834 2392
rect 1822 2368 1826 2372
rect 1862 2368 1866 2372
rect 1902 2388 1906 2392
rect 1886 2348 1890 2352
rect 1870 2328 1874 2332
rect 1870 2318 1874 2322
rect 1854 2308 1858 2312
rect 1846 2298 1850 2302
rect 1838 2278 1842 2282
rect 1862 2278 1866 2282
rect 1894 2318 1898 2322
rect 1886 2308 1890 2312
rect 1878 2298 1882 2302
rect 1886 2298 1890 2302
rect 1782 2248 1786 2252
rect 1774 2158 1778 2162
rect 1806 2218 1810 2222
rect 1782 2128 1786 2132
rect 1758 2098 1762 2102
rect 1766 2098 1770 2102
rect 1486 2058 1490 2062
rect 1694 2058 1698 2062
rect 1734 2058 1738 2062
rect 1526 2048 1530 2052
rect 1606 2048 1610 2052
rect 1542 2038 1546 2042
rect 1562 2003 1566 2007
rect 1569 2003 1573 2007
rect 1510 1998 1514 2002
rect 1502 1978 1506 1982
rect 1542 1968 1546 1972
rect 1550 1968 1554 1972
rect 1486 1938 1490 1942
rect 1414 1918 1418 1922
rect 1366 1898 1370 1902
rect 1430 1888 1434 1892
rect 1422 1868 1426 1872
rect 1446 1868 1450 1872
rect 1486 1918 1490 1922
rect 1526 1898 1530 1902
rect 1494 1888 1498 1892
rect 1502 1878 1506 1882
rect 1478 1868 1482 1872
rect 1326 1858 1330 1862
rect 1342 1858 1346 1862
rect 1358 1848 1362 1852
rect 1534 1868 1538 1872
rect 1510 1858 1514 1862
rect 1414 1838 1418 1842
rect 1438 1838 1442 1842
rect 1478 1838 1482 1842
rect 1470 1818 1474 1822
rect 1366 1768 1370 1772
rect 1318 1738 1322 1742
rect 1302 1688 1306 1692
rect 1310 1688 1314 1692
rect 1358 1718 1362 1722
rect 1406 1748 1410 1752
rect 1422 1748 1426 1752
rect 1382 1738 1386 1742
rect 1398 1738 1402 1742
rect 1406 1738 1410 1742
rect 1430 1738 1434 1742
rect 1446 1738 1450 1742
rect 1302 1668 1306 1672
rect 1334 1668 1338 1672
rect 1374 1668 1378 1672
rect 1262 1658 1266 1662
rect 1278 1658 1282 1662
rect 1214 1638 1218 1642
rect 1206 1598 1210 1602
rect 1198 1588 1202 1592
rect 1190 1578 1194 1582
rect 1190 1558 1194 1562
rect 1174 1548 1178 1552
rect 1142 1538 1146 1542
rect 1150 1538 1154 1542
rect 1118 1528 1122 1532
rect 1230 1548 1234 1552
rect 1158 1518 1162 1522
rect 1166 1498 1170 1502
rect 1174 1498 1178 1502
rect 1150 1488 1154 1492
rect 982 1448 986 1452
rect 1014 1448 1018 1452
rect 1054 1448 1058 1452
rect 1070 1448 1074 1452
rect 934 1438 938 1442
rect 966 1438 970 1442
rect 966 1398 970 1402
rect 950 1358 954 1362
rect 974 1358 978 1362
rect 870 1348 874 1352
rect 910 1348 914 1352
rect 934 1348 938 1352
rect 750 1338 754 1342
rect 782 1338 786 1342
rect 886 1338 890 1342
rect 774 1328 778 1332
rect 798 1328 802 1332
rect 878 1328 882 1332
rect 910 1328 914 1332
rect 726 1298 730 1302
rect 678 1288 682 1292
rect 702 1288 706 1292
rect 638 1278 642 1282
rect 646 1268 650 1272
rect 646 1258 650 1262
rect 654 1258 658 1262
rect 702 1258 706 1262
rect 686 1248 690 1252
rect 678 1168 682 1172
rect 566 1148 570 1152
rect 598 1148 602 1152
rect 614 1148 618 1152
rect 502 1138 506 1142
rect 510 1138 514 1142
rect 558 1138 562 1142
rect 462 1128 466 1132
rect 414 1068 418 1072
rect 422 1068 426 1072
rect 334 1058 338 1062
rect 398 1058 402 1062
rect 374 1048 378 1052
rect 382 1048 386 1052
rect 366 1038 370 1042
rect 350 1028 354 1032
rect 390 998 394 1002
rect 374 988 378 992
rect 430 1058 434 1062
rect 414 1038 418 1042
rect 502 1118 506 1122
rect 486 1088 490 1092
rect 462 1068 466 1072
rect 446 1018 450 1022
rect 414 1008 418 1012
rect 438 1008 442 1012
rect 406 988 410 992
rect 414 978 418 982
rect 358 958 362 962
rect 374 948 378 952
rect 342 938 346 942
rect 342 908 346 912
rect 310 868 314 872
rect 326 868 330 872
rect 286 858 290 862
rect 318 858 322 862
rect 278 758 282 762
rect 254 748 258 752
rect 270 748 274 752
rect 190 738 194 742
rect 238 738 242 742
rect 206 728 210 732
rect 230 728 234 732
rect 222 688 226 692
rect 206 678 210 682
rect 214 678 218 682
rect 190 668 194 672
rect 214 668 218 672
rect 174 648 178 652
rect 206 648 210 652
rect 230 578 234 582
rect 238 578 242 582
rect 182 558 186 562
rect 206 558 210 562
rect 158 548 162 552
rect 166 538 170 542
rect 190 548 194 552
rect 214 538 218 542
rect 198 518 202 522
rect 150 478 154 482
rect 158 478 162 482
rect 150 468 154 472
rect 110 448 114 452
rect 70 388 74 392
rect 86 388 90 392
rect 102 348 106 352
rect 78 338 82 342
rect 62 278 66 282
rect 38 248 42 252
rect 38 158 42 162
rect 62 138 66 142
rect 102 278 106 282
rect 118 348 122 352
rect 294 848 298 852
rect 350 838 354 842
rect 302 738 306 742
rect 262 718 266 722
rect 254 678 258 682
rect 294 708 298 712
rect 294 698 298 702
rect 758 1248 762 1252
rect 718 1178 722 1182
rect 750 1168 754 1172
rect 758 1168 762 1172
rect 726 1158 730 1162
rect 766 1158 770 1162
rect 670 1148 674 1152
rect 734 1148 738 1152
rect 742 1148 746 1152
rect 662 1138 666 1142
rect 630 1128 634 1132
rect 582 1118 586 1122
rect 574 1098 578 1102
rect 614 1098 618 1102
rect 590 1078 594 1082
rect 534 1048 538 1052
rect 550 1048 554 1052
rect 538 1003 542 1007
rect 545 1003 549 1007
rect 518 998 522 1002
rect 454 988 458 992
rect 502 988 506 992
rect 534 988 538 992
rect 470 948 474 952
rect 494 948 498 952
rect 446 938 450 942
rect 470 938 474 942
rect 406 918 410 922
rect 422 898 426 902
rect 438 898 442 902
rect 430 868 434 872
rect 390 858 394 862
rect 406 858 410 862
rect 486 918 490 922
rect 526 928 530 932
rect 526 918 530 922
rect 510 898 514 902
rect 478 858 482 862
rect 518 858 522 862
rect 374 838 378 842
rect 454 838 458 842
rect 462 768 466 772
rect 518 768 522 772
rect 398 758 402 762
rect 478 758 482 762
rect 494 758 498 762
rect 630 998 634 1002
rect 646 998 650 1002
rect 750 1128 754 1132
rect 742 1098 746 1102
rect 686 1078 690 1082
rect 710 1078 714 1082
rect 734 1058 738 1062
rect 710 1028 714 1032
rect 678 988 682 992
rect 646 948 650 952
rect 614 938 618 942
rect 566 918 570 922
rect 614 918 618 922
rect 598 908 602 912
rect 574 888 578 892
rect 598 888 602 892
rect 590 868 594 872
rect 630 878 634 882
rect 574 858 578 862
rect 606 858 610 862
rect 670 948 674 952
rect 702 948 706 952
rect 694 938 698 942
rect 702 918 706 922
rect 670 908 674 912
rect 638 858 642 862
rect 654 848 658 852
rect 662 838 666 842
rect 590 808 594 812
rect 538 803 542 807
rect 545 803 549 807
rect 566 798 570 802
rect 598 788 602 792
rect 582 758 586 762
rect 462 748 466 752
rect 478 748 482 752
rect 382 678 386 682
rect 446 708 450 712
rect 334 668 338 672
rect 358 668 362 672
rect 326 658 330 662
rect 286 638 290 642
rect 270 628 274 632
rect 326 648 330 652
rect 302 638 306 642
rect 294 618 298 622
rect 254 578 258 582
rect 254 568 258 572
rect 350 638 354 642
rect 366 638 370 642
rect 358 588 362 592
rect 422 638 426 642
rect 694 848 698 852
rect 694 798 698 802
rect 718 968 722 972
rect 734 938 738 942
rect 718 868 722 872
rect 742 848 746 852
rect 614 768 618 772
rect 654 768 658 772
rect 630 758 634 762
rect 590 738 594 742
rect 486 698 490 702
rect 598 728 602 732
rect 574 698 578 702
rect 518 678 522 682
rect 582 678 586 682
rect 630 678 634 682
rect 494 668 498 672
rect 470 658 474 662
rect 518 658 522 662
rect 446 648 450 652
rect 478 648 482 652
rect 518 648 522 652
rect 550 648 554 652
rect 494 638 498 642
rect 382 568 386 572
rect 342 558 346 562
rect 262 548 266 552
rect 270 548 274 552
rect 390 547 394 551
rect 494 618 498 622
rect 538 603 542 607
rect 545 603 549 607
rect 534 588 538 592
rect 478 558 482 562
rect 310 538 314 542
rect 246 508 250 512
rect 302 508 306 512
rect 438 528 442 532
rect 270 468 274 472
rect 350 468 354 472
rect 414 468 418 472
rect 430 468 434 472
rect 142 448 146 452
rect 158 438 162 442
rect 158 418 162 422
rect 190 458 194 462
rect 174 428 178 432
rect 286 458 290 462
rect 318 458 322 462
rect 334 458 338 462
rect 406 458 410 462
rect 222 438 226 442
rect 206 418 210 422
rect 166 388 170 392
rect 150 348 154 352
rect 174 348 178 352
rect 126 338 130 342
rect 174 328 178 332
rect 166 318 170 322
rect 158 298 162 302
rect 94 258 98 262
rect 134 258 138 262
rect 142 258 146 262
rect 110 238 114 242
rect 102 188 106 192
rect 134 168 138 172
rect 110 148 114 152
rect 190 328 194 332
rect 182 298 186 302
rect 214 348 218 352
rect 286 428 290 432
rect 278 378 282 382
rect 222 338 226 342
rect 230 318 234 322
rect 198 308 202 312
rect 326 358 330 362
rect 502 518 506 522
rect 478 498 482 502
rect 566 628 570 632
rect 638 668 642 672
rect 686 758 690 762
rect 718 758 722 762
rect 718 748 722 752
rect 702 728 706 732
rect 702 718 706 722
rect 686 698 690 702
rect 694 698 698 702
rect 782 1298 786 1302
rect 790 1278 794 1282
rect 822 1268 826 1272
rect 838 1258 842 1262
rect 790 1248 794 1252
rect 830 1238 834 1242
rect 894 1288 898 1292
rect 854 1278 858 1282
rect 870 1258 874 1262
rect 838 1218 842 1222
rect 878 1208 882 1212
rect 878 1198 882 1202
rect 790 1168 794 1172
rect 870 1168 874 1172
rect 790 1158 794 1162
rect 838 1148 842 1152
rect 790 1108 794 1112
rect 790 1068 794 1072
rect 782 998 786 1002
rect 806 1138 810 1142
rect 806 1108 810 1112
rect 806 1088 810 1092
rect 806 1068 810 1072
rect 846 1108 850 1112
rect 838 1098 842 1102
rect 806 1038 810 1042
rect 902 1148 906 1152
rect 950 1318 954 1322
rect 934 1308 938 1312
rect 926 1298 930 1302
rect 1030 1358 1034 1362
rect 1070 1438 1074 1442
rect 1118 1458 1122 1462
rect 1142 1458 1146 1462
rect 1142 1448 1146 1452
rect 1110 1438 1114 1442
rect 1094 1418 1098 1422
rect 1158 1408 1162 1412
rect 1086 1378 1090 1382
rect 1094 1378 1098 1382
rect 1078 1368 1082 1372
rect 1110 1358 1114 1362
rect 1014 1348 1018 1352
rect 1038 1348 1042 1352
rect 1102 1348 1106 1352
rect 998 1328 1002 1332
rect 966 1278 970 1282
rect 990 1268 994 1272
rect 1006 1208 1010 1212
rect 974 1198 978 1202
rect 934 1158 938 1162
rect 942 1148 946 1152
rect 1014 1148 1018 1152
rect 942 1138 946 1142
rect 886 1128 890 1132
rect 910 1128 914 1132
rect 854 1078 858 1082
rect 870 1068 874 1072
rect 886 1068 890 1072
rect 958 1108 962 1112
rect 918 1058 922 1062
rect 934 1058 938 1062
rect 950 1058 954 1062
rect 830 1038 834 1042
rect 902 1038 906 1042
rect 870 1018 874 1022
rect 838 988 842 992
rect 822 968 826 972
rect 798 948 802 952
rect 814 948 818 952
rect 830 948 834 952
rect 822 938 826 942
rect 774 928 778 932
rect 758 878 762 882
rect 790 908 794 912
rect 798 878 802 882
rect 822 878 826 882
rect 854 938 858 942
rect 838 928 842 932
rect 958 988 962 992
rect 918 968 922 972
rect 902 938 906 942
rect 862 918 866 922
rect 838 888 842 892
rect 918 918 922 922
rect 878 898 882 902
rect 894 898 898 902
rect 990 1138 994 1142
rect 1046 1338 1050 1342
rect 1078 1338 1082 1342
rect 1142 1338 1146 1342
rect 1050 1303 1054 1307
rect 1057 1303 1061 1307
rect 1054 1288 1058 1292
rect 1118 1308 1122 1312
rect 1078 1268 1082 1272
rect 1086 1268 1090 1272
rect 1094 1268 1098 1272
rect 1110 1268 1114 1272
rect 1110 1238 1114 1242
rect 1094 1218 1098 1222
rect 1126 1288 1130 1292
rect 1142 1278 1146 1282
rect 1206 1448 1210 1452
rect 1198 1438 1202 1442
rect 1198 1368 1202 1372
rect 1262 1538 1266 1542
rect 1230 1488 1234 1492
rect 1254 1488 1258 1492
rect 1334 1648 1338 1652
rect 1318 1608 1322 1612
rect 1334 1588 1338 1592
rect 1318 1578 1322 1582
rect 1334 1578 1338 1582
rect 1366 1558 1370 1562
rect 1318 1548 1322 1552
rect 1374 1538 1378 1542
rect 1366 1528 1370 1532
rect 1262 1468 1266 1472
rect 1278 1458 1282 1462
rect 1302 1458 1306 1462
rect 1342 1458 1346 1462
rect 1238 1428 1242 1432
rect 1230 1388 1234 1392
rect 1270 1408 1274 1412
rect 1246 1378 1250 1382
rect 1214 1358 1218 1362
rect 1262 1358 1266 1362
rect 1230 1348 1234 1352
rect 1222 1338 1226 1342
rect 1270 1338 1274 1342
rect 1254 1328 1258 1332
rect 1174 1308 1178 1312
rect 1190 1308 1194 1312
rect 1206 1298 1210 1302
rect 1198 1278 1202 1282
rect 1126 1268 1130 1272
rect 1166 1268 1170 1272
rect 1214 1268 1218 1272
rect 1222 1268 1226 1272
rect 1142 1258 1146 1262
rect 1134 1238 1138 1242
rect 1078 1158 1082 1162
rect 1150 1158 1154 1162
rect 1182 1258 1186 1262
rect 1054 1148 1058 1152
rect 1126 1148 1130 1152
rect 1158 1148 1162 1152
rect 1054 1128 1058 1132
rect 1078 1128 1082 1132
rect 1050 1103 1054 1107
rect 1057 1103 1061 1107
rect 1006 1088 1010 1092
rect 1070 1078 1074 1082
rect 1030 1068 1034 1072
rect 1046 1058 1050 1062
rect 1062 1058 1066 1062
rect 998 1048 1002 1052
rect 1022 988 1026 992
rect 1030 968 1034 972
rect 1062 968 1066 972
rect 990 938 994 942
rect 990 918 994 922
rect 982 888 986 892
rect 782 858 786 862
rect 782 848 786 852
rect 806 848 810 852
rect 806 828 810 832
rect 782 808 786 812
rect 822 788 826 792
rect 806 758 810 762
rect 766 748 770 752
rect 734 708 738 712
rect 766 708 770 712
rect 758 698 762 702
rect 766 678 770 682
rect 726 668 730 672
rect 654 658 658 662
rect 718 658 722 662
rect 774 658 778 662
rect 606 638 610 642
rect 590 598 594 602
rect 566 578 570 582
rect 574 568 578 572
rect 606 568 610 572
rect 646 568 650 572
rect 622 558 626 562
rect 622 548 626 552
rect 630 548 634 552
rect 574 538 578 542
rect 614 538 618 542
rect 598 498 602 502
rect 558 488 562 492
rect 726 638 730 642
rect 750 598 754 602
rect 1050 903 1054 907
rect 1057 903 1061 907
rect 990 878 994 882
rect 1006 878 1010 882
rect 926 868 930 872
rect 870 858 874 862
rect 886 858 890 862
rect 910 848 914 852
rect 870 818 874 822
rect 910 828 914 832
rect 966 858 970 862
rect 934 838 938 842
rect 958 838 962 842
rect 926 828 930 832
rect 966 828 970 832
rect 942 818 946 822
rect 894 798 898 802
rect 950 798 954 802
rect 862 788 866 792
rect 926 788 930 792
rect 886 768 890 772
rect 838 758 842 762
rect 878 758 882 762
rect 830 728 834 732
rect 862 708 866 712
rect 822 698 826 702
rect 830 678 834 682
rect 902 758 906 762
rect 910 678 914 682
rect 846 668 850 672
rect 966 768 970 772
rect 974 758 978 762
rect 950 728 954 732
rect 966 718 970 722
rect 942 708 946 712
rect 1006 868 1010 872
rect 1070 868 1074 872
rect 1094 1098 1098 1102
rect 1102 1088 1106 1092
rect 1086 1068 1090 1072
rect 1118 1028 1122 1032
rect 1110 998 1114 1002
rect 1166 1138 1170 1142
rect 1150 1128 1154 1132
rect 1134 1078 1138 1082
rect 1134 1048 1138 1052
rect 1142 1048 1146 1052
rect 1158 1048 1162 1052
rect 1166 1038 1170 1042
rect 1166 1028 1170 1032
rect 1150 998 1154 1002
rect 1142 988 1146 992
rect 1134 968 1138 972
rect 1118 958 1122 962
rect 1262 1268 1266 1272
rect 1422 1688 1426 1692
rect 1438 1688 1442 1692
rect 1454 1688 1458 1692
rect 1526 1848 1530 1852
rect 1502 1808 1506 1812
rect 1558 1948 1562 1952
rect 1590 1948 1594 1952
rect 1702 2048 1706 2052
rect 1670 2038 1674 2042
rect 1670 2018 1674 2022
rect 1646 2008 1650 2012
rect 1678 1998 1682 2002
rect 1686 1958 1690 1962
rect 1662 1948 1666 1952
rect 1614 1928 1618 1932
rect 1598 1888 1602 1892
rect 1598 1868 1602 1872
rect 1614 1868 1618 1872
rect 1638 1868 1642 1872
rect 1566 1858 1570 1862
rect 1562 1803 1566 1807
rect 1569 1803 1573 1807
rect 1542 1788 1546 1792
rect 1526 1768 1530 1772
rect 1486 1728 1490 1732
rect 1494 1728 1498 1732
rect 1470 1708 1474 1712
rect 1478 1668 1482 1672
rect 1446 1658 1450 1662
rect 1446 1648 1450 1652
rect 1438 1578 1442 1582
rect 1462 1648 1466 1652
rect 1518 1688 1522 1692
rect 1678 1778 1682 1782
rect 1662 1768 1666 1772
rect 1550 1758 1554 1762
rect 1574 1748 1578 1752
rect 1662 1748 1666 1752
rect 1614 1738 1618 1742
rect 1614 1728 1618 1732
rect 1606 1698 1610 1702
rect 1502 1658 1506 1662
rect 1526 1658 1530 1662
rect 1598 1648 1602 1652
rect 1510 1638 1514 1642
rect 1562 1603 1566 1607
rect 1569 1603 1573 1607
rect 1478 1588 1482 1592
rect 1502 1588 1506 1592
rect 1486 1558 1490 1562
rect 1406 1548 1410 1552
rect 1390 1538 1394 1542
rect 1422 1508 1426 1512
rect 1414 1498 1418 1502
rect 1406 1488 1410 1492
rect 1430 1498 1434 1502
rect 1414 1458 1418 1462
rect 1286 1448 1290 1452
rect 1366 1448 1370 1452
rect 1390 1438 1394 1442
rect 1366 1418 1370 1422
rect 1406 1428 1410 1432
rect 1398 1408 1402 1412
rect 1366 1398 1370 1402
rect 1342 1358 1346 1362
rect 1366 1358 1370 1362
rect 1438 1458 1442 1462
rect 1446 1438 1450 1442
rect 1430 1398 1434 1402
rect 1438 1398 1442 1402
rect 1534 1578 1538 1582
rect 1590 1558 1594 1562
rect 1470 1548 1474 1552
rect 1550 1548 1554 1552
rect 1574 1548 1578 1552
rect 1494 1538 1498 1542
rect 1550 1538 1554 1542
rect 1598 1538 1602 1542
rect 1526 1528 1530 1532
rect 1518 1508 1522 1512
rect 1478 1488 1482 1492
rect 1502 1488 1506 1492
rect 1534 1488 1538 1492
rect 1470 1458 1474 1462
rect 1462 1448 1466 1452
rect 1510 1448 1514 1452
rect 1454 1388 1458 1392
rect 1422 1358 1426 1362
rect 1430 1348 1434 1352
rect 1286 1308 1290 1312
rect 1294 1298 1298 1302
rect 1334 1328 1338 1332
rect 1318 1318 1322 1322
rect 1406 1338 1410 1342
rect 1422 1338 1426 1342
rect 1470 1338 1474 1342
rect 1342 1308 1346 1312
rect 1334 1298 1338 1302
rect 1310 1288 1314 1292
rect 1342 1288 1346 1292
rect 1326 1278 1330 1282
rect 1342 1268 1346 1272
rect 1358 1268 1362 1272
rect 1214 1248 1218 1252
rect 1278 1248 1282 1252
rect 1206 1218 1210 1222
rect 1190 1188 1194 1192
rect 1182 1128 1186 1132
rect 1190 1068 1194 1072
rect 1190 1058 1194 1062
rect 1182 1028 1186 1032
rect 1174 1018 1178 1022
rect 1134 948 1138 952
rect 1142 948 1146 952
rect 1174 948 1178 952
rect 1126 878 1130 882
rect 1126 858 1130 862
rect 1022 768 1026 772
rect 1030 768 1034 772
rect 990 758 994 762
rect 990 738 994 742
rect 998 728 1002 732
rect 982 668 986 672
rect 822 648 826 652
rect 902 658 906 662
rect 918 658 922 662
rect 966 658 970 662
rect 686 558 690 562
rect 782 558 786 562
rect 790 558 794 562
rect 758 548 762 552
rect 646 538 650 542
rect 766 538 770 542
rect 790 538 794 542
rect 814 538 818 542
rect 630 498 634 502
rect 454 468 458 472
rect 494 468 498 472
rect 438 448 442 452
rect 406 438 410 442
rect 366 388 370 392
rect 350 378 354 382
rect 350 348 354 352
rect 358 348 362 352
rect 382 358 386 362
rect 390 358 394 362
rect 406 358 410 362
rect 414 358 418 362
rect 446 358 450 362
rect 334 328 338 332
rect 286 308 290 312
rect 310 298 314 302
rect 222 288 226 292
rect 374 298 378 302
rect 398 308 402 312
rect 318 288 322 292
rect 366 288 370 292
rect 206 248 210 252
rect 222 248 226 252
rect 166 188 170 192
rect 222 188 226 192
rect 198 178 202 182
rect 182 158 186 162
rect 190 158 194 162
rect 214 158 218 162
rect 206 148 210 152
rect 446 348 450 352
rect 542 448 546 452
rect 470 428 474 432
rect 598 418 602 422
rect 538 403 542 407
rect 545 403 549 407
rect 502 378 506 382
rect 590 378 594 382
rect 478 358 482 362
rect 438 338 442 342
rect 454 338 458 342
rect 422 318 426 322
rect 462 318 466 322
rect 422 308 426 312
rect 438 308 442 312
rect 430 298 434 302
rect 406 288 410 292
rect 542 347 546 351
rect 670 518 674 522
rect 686 518 690 522
rect 654 478 658 482
rect 622 458 626 462
rect 630 448 634 452
rect 614 438 618 442
rect 630 428 634 432
rect 614 398 618 402
rect 662 438 666 442
rect 678 378 682 382
rect 622 358 626 362
rect 654 358 658 362
rect 614 338 618 342
rect 470 298 474 302
rect 438 268 442 272
rect 454 268 458 272
rect 502 268 506 272
rect 422 248 426 252
rect 582 318 586 322
rect 566 298 570 302
rect 574 298 578 302
rect 542 258 546 262
rect 558 248 562 252
rect 358 228 362 232
rect 478 228 482 232
rect 326 218 330 222
rect 294 178 298 182
rect 278 168 282 172
rect 286 168 290 172
rect 230 158 234 162
rect 238 148 242 152
rect 254 148 258 152
rect 150 78 154 82
rect 310 168 314 172
rect 310 148 314 152
rect 318 138 322 142
rect 294 128 298 132
rect 230 78 234 82
rect 78 68 82 72
rect 158 68 162 72
rect 494 218 498 222
rect 430 188 434 192
rect 462 188 466 192
rect 406 168 410 172
rect 374 148 378 152
rect 310 118 314 122
rect 278 88 282 92
rect 302 88 306 92
rect 326 78 330 82
rect 538 203 542 207
rect 545 203 549 207
rect 566 198 570 202
rect 510 178 514 182
rect 494 168 498 172
rect 430 158 434 162
rect 454 148 458 152
rect 486 148 490 152
rect 510 148 514 152
rect 494 138 498 142
rect 526 138 530 142
rect 422 128 426 132
rect 438 128 442 132
rect 414 118 418 122
rect 206 58 210 62
rect 454 78 458 82
rect 478 78 482 82
rect 430 68 434 72
rect 366 58 370 62
rect 438 58 442 62
rect 598 298 602 302
rect 782 508 786 512
rect 758 488 762 492
rect 750 478 754 482
rect 870 648 874 652
rect 894 648 898 652
rect 846 638 850 642
rect 878 638 882 642
rect 886 638 890 642
rect 982 648 986 652
rect 1022 708 1026 712
rect 1022 698 1026 702
rect 1238 1238 1242 1242
rect 1246 1148 1250 1152
rect 1222 1038 1226 1042
rect 1342 1198 1346 1202
rect 1294 1138 1298 1142
rect 1254 1128 1258 1132
rect 1294 1128 1298 1132
rect 1246 1058 1250 1062
rect 1278 1058 1282 1062
rect 1390 1328 1394 1332
rect 1382 1278 1386 1282
rect 1382 1248 1386 1252
rect 1374 1208 1378 1212
rect 1398 1258 1402 1262
rect 1430 1298 1434 1302
rect 1494 1438 1498 1442
rect 1590 1438 1594 1442
rect 1510 1398 1514 1402
rect 1486 1288 1490 1292
rect 1454 1278 1458 1282
rect 1470 1278 1474 1282
rect 1470 1258 1474 1262
rect 1414 1248 1418 1252
rect 1422 1248 1426 1252
rect 1562 1403 1566 1407
rect 1569 1403 1573 1407
rect 1686 1758 1690 1762
rect 1726 2038 1730 2042
rect 1790 2118 1794 2122
rect 1798 2108 1802 2112
rect 1790 2078 1794 2082
rect 1838 2218 1842 2222
rect 1814 2178 1818 2182
rect 1926 2438 1930 2442
rect 1942 2428 1946 2432
rect 1926 2368 1930 2372
rect 1990 2528 1994 2532
rect 2006 2518 2010 2522
rect 1990 2508 1994 2512
rect 1966 2488 1970 2492
rect 2022 2518 2026 2522
rect 2014 2488 2018 2492
rect 2006 2478 2010 2482
rect 1966 2428 1970 2432
rect 1990 2388 1994 2392
rect 1926 2358 1930 2362
rect 1958 2358 1962 2362
rect 1934 2348 1938 2352
rect 1942 2348 1946 2352
rect 1950 2348 1954 2352
rect 1910 2318 1914 2322
rect 1918 2318 1922 2322
rect 1926 2308 1930 2312
rect 1942 2318 1946 2322
rect 1950 2298 1954 2302
rect 1950 2288 1954 2292
rect 2054 2628 2058 2632
rect 2062 2618 2066 2622
rect 2054 2578 2058 2582
rect 2046 2548 2050 2552
rect 2054 2528 2058 2532
rect 2038 2518 2042 2522
rect 2070 2598 2074 2602
rect 2158 2748 2162 2752
rect 2214 2868 2218 2872
rect 2262 2908 2266 2912
rect 2190 2778 2194 2782
rect 2238 2778 2242 2782
rect 2230 2768 2234 2772
rect 2206 2758 2210 2762
rect 2222 2758 2226 2762
rect 2230 2748 2234 2752
rect 2182 2738 2186 2742
rect 2190 2738 2194 2742
rect 2254 2738 2258 2742
rect 2158 2728 2162 2732
rect 2246 2728 2250 2732
rect 2206 2698 2210 2702
rect 2190 2678 2194 2682
rect 2238 2678 2242 2682
rect 2254 2678 2258 2682
rect 2294 2948 2298 2952
rect 2294 2938 2298 2942
rect 2318 2938 2322 2942
rect 2286 2928 2290 2932
rect 2278 2918 2282 2922
rect 2286 2808 2290 2812
rect 2318 2908 2322 2912
rect 2302 2888 2306 2892
rect 2310 2888 2314 2892
rect 2318 2868 2322 2872
rect 2302 2848 2306 2852
rect 2606 3718 2610 3722
rect 2630 3718 2634 3722
rect 2590 3708 2594 3712
rect 2742 3968 2746 3972
rect 2798 4048 2802 4052
rect 2790 3968 2794 3972
rect 2726 3958 2730 3962
rect 2734 3958 2738 3962
rect 2774 3958 2778 3962
rect 2822 4208 2826 4212
rect 2878 4488 2882 4492
rect 2886 4468 2890 4472
rect 2894 4458 2898 4462
rect 2886 4378 2890 4382
rect 2878 4328 2882 4332
rect 2846 4218 2850 4222
rect 2942 4508 2946 4512
rect 2950 4448 2954 4452
rect 2982 4468 2986 4472
rect 2998 4458 3002 4462
rect 2982 4448 2986 4452
rect 3022 4508 3026 4512
rect 4114 4903 4118 4907
rect 4121 4903 4125 4907
rect 3622 4888 3626 4892
rect 3830 4888 3834 4892
rect 3990 4888 3994 4892
rect 4078 4888 4082 4892
rect 5006 4888 5010 4892
rect 5166 4888 5170 4892
rect 3214 4878 3218 4882
rect 3342 4878 3346 4882
rect 3558 4878 3562 4882
rect 4238 4878 4242 4882
rect 3350 4868 3354 4872
rect 3190 4858 3194 4862
rect 3230 4858 3234 4862
rect 3286 4858 3290 4862
rect 3358 4858 3362 4862
rect 3190 4848 3194 4852
rect 3254 4848 3258 4852
rect 3126 4838 3130 4842
rect 3150 4838 3154 4842
rect 3222 4828 3226 4832
rect 3222 4818 3226 4822
rect 3094 4788 3098 4792
rect 3206 4778 3210 4782
rect 3238 4768 3242 4772
rect 3334 4798 3338 4802
rect 3238 4748 3242 4752
rect 3254 4748 3258 4752
rect 3334 4748 3338 4752
rect 3110 4728 3114 4732
rect 3118 4718 3122 4722
rect 3098 4703 3102 4707
rect 3105 4703 3109 4707
rect 3174 4738 3178 4742
rect 3206 4738 3210 4742
rect 3142 4698 3146 4702
rect 3078 4688 3082 4692
rect 3150 4688 3154 4692
rect 3190 4728 3194 4732
rect 3174 4718 3178 4722
rect 3070 4678 3074 4682
rect 3158 4678 3162 4682
rect 3062 4658 3066 4662
rect 3054 4648 3058 4652
rect 3062 4648 3066 4652
rect 3054 4598 3058 4602
rect 3062 4568 3066 4572
rect 2950 4438 2954 4442
rect 2958 4418 2962 4422
rect 2894 4368 2898 4372
rect 2910 4368 2914 4372
rect 2918 4328 2922 4332
rect 2910 4318 2914 4322
rect 2934 4318 2938 4322
rect 3022 4368 3026 4372
rect 3006 4348 3010 4352
rect 2982 4298 2986 4302
rect 2926 4258 2930 4262
rect 2966 4258 2970 4262
rect 2990 4248 2994 4252
rect 2918 4238 2922 4242
rect 2854 4198 2858 4202
rect 2846 4188 2850 4192
rect 2846 4148 2850 4152
rect 2862 4138 2866 4142
rect 2878 4198 2882 4202
rect 2918 4168 2922 4172
rect 2822 4098 2826 4102
rect 2870 4098 2874 4102
rect 2814 4088 2818 4092
rect 2838 4068 2842 4072
rect 2854 4068 2858 4072
rect 2814 4058 2818 4062
rect 2830 4048 2834 4052
rect 2830 4038 2834 4042
rect 2830 3988 2834 3992
rect 2814 3958 2818 3962
rect 2830 3958 2834 3962
rect 2782 3948 2786 3952
rect 2758 3938 2762 3942
rect 2726 3928 2730 3932
rect 2734 3928 2738 3932
rect 2766 3918 2770 3922
rect 2774 3908 2778 3912
rect 2758 3878 2762 3882
rect 2734 3868 2738 3872
rect 2774 3868 2778 3872
rect 2902 4118 2906 4122
rect 2902 4088 2906 4092
rect 2926 4128 2930 4132
rect 2950 4118 2954 4122
rect 2998 4188 3002 4192
rect 2998 4138 3002 4142
rect 3054 4438 3058 4442
rect 3062 4398 3066 4402
rect 3054 4388 3058 4392
rect 3046 4268 3050 4272
rect 3022 4248 3026 4252
rect 3030 4218 3034 4222
rect 3062 4268 3066 4272
rect 3038 4158 3042 4162
rect 3182 4708 3186 4712
rect 3198 4708 3202 4712
rect 3182 4698 3186 4702
rect 3238 4738 3242 4742
rect 3262 4738 3266 4742
rect 3222 4718 3226 4722
rect 3214 4698 3218 4702
rect 3230 4688 3234 4692
rect 3294 4728 3298 4732
rect 3150 4668 3154 4672
rect 3174 4668 3178 4672
rect 3214 4668 3218 4672
rect 3230 4668 3234 4672
rect 3238 4668 3242 4672
rect 3086 4638 3090 4642
rect 3078 4578 3082 4582
rect 3086 4568 3090 4572
rect 3086 4538 3090 4542
rect 3166 4658 3170 4662
rect 3110 4648 3114 4652
rect 3134 4558 3138 4562
rect 3102 4548 3106 4552
rect 3150 4548 3154 4552
rect 3190 4658 3194 4662
rect 3190 4638 3194 4642
rect 3142 4538 3146 4542
rect 3158 4538 3162 4542
rect 3126 4508 3130 4512
rect 3098 4503 3102 4507
rect 3105 4503 3109 4507
rect 3126 4488 3130 4492
rect 3086 4448 3090 4452
rect 3110 4448 3114 4452
rect 3134 4448 3138 4452
rect 3126 4408 3130 4412
rect 3086 4348 3090 4352
rect 3134 4368 3138 4372
rect 3150 4478 3154 4482
rect 3182 4508 3186 4512
rect 3198 4628 3202 4632
rect 3238 4588 3242 4592
rect 3230 4548 3234 4552
rect 3294 4638 3298 4642
rect 3334 4698 3338 4702
rect 3318 4658 3322 4662
rect 3318 4628 3322 4632
rect 3262 4478 3266 4482
rect 3206 4468 3210 4472
rect 3246 4468 3250 4472
rect 3278 4468 3282 4472
rect 3214 4458 3218 4462
rect 3230 4458 3234 4462
rect 3254 4458 3258 4462
rect 3174 4438 3178 4442
rect 3246 4448 3250 4452
rect 3214 4418 3218 4422
rect 3174 4398 3178 4402
rect 3190 4398 3194 4402
rect 3150 4368 3154 4372
rect 3142 4358 3146 4362
rect 3190 4368 3194 4372
rect 3134 4348 3138 4352
rect 3142 4348 3146 4352
rect 3166 4348 3170 4352
rect 3142 4338 3146 4342
rect 3158 4338 3162 4342
rect 3098 4303 3102 4307
rect 3105 4303 3109 4307
rect 3102 4268 3106 4272
rect 3070 4218 3074 4222
rect 3150 4278 3154 4282
rect 3158 4268 3162 4272
rect 3190 4338 3194 4342
rect 3198 4318 3202 4322
rect 3238 4278 3242 4282
rect 3150 4258 3154 4262
rect 3182 4258 3186 4262
rect 3198 4258 3202 4262
rect 3086 4188 3090 4192
rect 3078 4148 3082 4152
rect 3086 4138 3090 4142
rect 3294 4488 3298 4492
rect 3262 4378 3266 4382
rect 3302 4368 3306 4372
rect 3366 4828 3370 4832
rect 3398 4858 3402 4862
rect 3478 4858 3482 4862
rect 3790 4858 3794 4862
rect 3382 4838 3386 4842
rect 3406 4838 3410 4842
rect 3462 4828 3466 4832
rect 3582 4828 3586 4832
rect 3374 4818 3378 4822
rect 3446 4798 3450 4802
rect 3406 4788 3410 4792
rect 3430 4788 3434 4792
rect 3414 4778 3418 4782
rect 3430 4778 3434 4782
rect 3610 4803 3614 4807
rect 3617 4803 3621 4807
rect 3694 4828 3698 4832
rect 3734 4818 3738 4822
rect 3790 4838 3794 4842
rect 3782 4828 3786 4832
rect 3766 4808 3770 4812
rect 3670 4778 3674 4782
rect 3582 4768 3586 4772
rect 3382 4758 3386 4762
rect 3366 4728 3370 4732
rect 3406 4748 3410 4752
rect 3414 4738 3418 4742
rect 3438 4748 3442 4752
rect 3446 4738 3450 4742
rect 3382 4698 3386 4702
rect 3366 4678 3370 4682
rect 3414 4678 3418 4682
rect 3422 4678 3426 4682
rect 3374 4668 3378 4672
rect 3406 4668 3410 4672
rect 3366 4658 3370 4662
rect 3398 4658 3402 4662
rect 3350 4628 3354 4632
rect 3350 4568 3354 4572
rect 3334 4548 3338 4552
rect 3350 4548 3354 4552
rect 3318 4528 3322 4532
rect 3334 4478 3338 4482
rect 3406 4568 3410 4572
rect 3406 4558 3410 4562
rect 3374 4518 3378 4522
rect 3398 4508 3402 4512
rect 3438 4538 3442 4542
rect 3510 4758 3514 4762
rect 3470 4748 3474 4752
rect 3606 4748 3610 4752
rect 3470 4738 3474 4742
rect 3486 4728 3490 4732
rect 3574 4728 3578 4732
rect 3470 4688 3474 4692
rect 3550 4718 3554 4722
rect 3558 4718 3562 4722
rect 3574 4688 3578 4692
rect 3534 4678 3538 4682
rect 3582 4668 3586 4672
rect 3806 4788 3810 4792
rect 3862 4868 3866 4872
rect 3878 4868 3882 4872
rect 4206 4868 4210 4872
rect 3854 4858 3858 4862
rect 3870 4858 3874 4862
rect 3878 4848 3882 4852
rect 4046 4848 4050 4852
rect 3918 4838 3922 4842
rect 4182 4858 4186 4862
rect 4214 4858 4218 4862
rect 4142 4838 4146 4842
rect 3910 4828 3914 4832
rect 4062 4828 4066 4832
rect 4166 4828 4170 4832
rect 3830 4788 3834 4792
rect 3974 4798 3978 4802
rect 3822 4768 3826 4772
rect 3806 4758 3810 4762
rect 3846 4758 3850 4762
rect 3894 4758 3898 4762
rect 3774 4748 3778 4752
rect 3790 4748 3794 4752
rect 3622 4718 3626 4722
rect 3710 4738 3714 4742
rect 3766 4738 3770 4742
rect 3638 4708 3642 4712
rect 3654 4718 3658 4722
rect 3614 4678 3618 4682
rect 3646 4678 3650 4682
rect 3550 4658 3554 4662
rect 3470 4648 3474 4652
rect 3550 4648 3554 4652
rect 3582 4648 3586 4652
rect 3646 4648 3650 4652
rect 3494 4548 3498 4552
rect 3470 4538 3474 4542
rect 3462 4518 3466 4522
rect 3454 4498 3458 4502
rect 3486 4478 3490 4482
rect 3366 4468 3370 4472
rect 3454 4458 3458 4462
rect 3358 4448 3362 4452
rect 3374 4388 3378 4392
rect 3406 4388 3410 4392
rect 3270 4358 3274 4362
rect 3278 4358 3282 4362
rect 3310 4358 3314 4362
rect 3342 4358 3346 4362
rect 3254 4208 3258 4212
rect 3174 4168 3178 4172
rect 3222 4168 3226 4172
rect 3246 4168 3250 4172
rect 3134 4138 3138 4142
rect 3070 4128 3074 4132
rect 3102 4128 3106 4132
rect 3022 4118 3026 4122
rect 3030 4108 3034 4112
rect 2990 4098 2994 4102
rect 3006 4098 3010 4102
rect 2982 4088 2986 4092
rect 2934 4058 2938 4062
rect 3022 4078 3026 4082
rect 3014 4068 3018 4072
rect 3070 4108 3074 4112
rect 3054 4088 3058 4092
rect 3098 4103 3102 4107
rect 3105 4103 3109 4107
rect 3078 4088 3082 4092
rect 3086 4088 3090 4092
rect 3054 4068 3058 4072
rect 2958 4058 2962 4062
rect 3046 4058 3050 4062
rect 3094 4058 3098 4062
rect 2894 4048 2898 4052
rect 2918 4048 2922 4052
rect 2950 4048 2954 4052
rect 3014 4048 3018 4052
rect 2990 4018 2994 4022
rect 2974 4008 2978 4012
rect 2878 3998 2882 4002
rect 2974 3988 2978 3992
rect 2902 3978 2906 3982
rect 2870 3958 2874 3962
rect 2878 3958 2882 3962
rect 2806 3928 2810 3932
rect 2854 3928 2858 3932
rect 2790 3908 2794 3912
rect 2814 3888 2818 3892
rect 2782 3858 2786 3862
rect 2806 3858 2810 3862
rect 2726 3848 2730 3852
rect 2742 3848 2746 3852
rect 2742 3838 2746 3842
rect 2702 3828 2706 3832
rect 2662 3788 2666 3792
rect 2670 3758 2674 3762
rect 2646 3728 2650 3732
rect 2638 3708 2642 3712
rect 2766 3848 2770 3852
rect 2750 3828 2754 3832
rect 2790 3818 2794 3822
rect 2782 3778 2786 3782
rect 2694 3728 2698 3732
rect 2654 3688 2658 3692
rect 2622 3668 2626 3672
rect 2654 3668 2658 3672
rect 2614 3658 2618 3662
rect 2710 3658 2714 3662
rect 2646 3648 2650 3652
rect 2678 3648 2682 3652
rect 2550 3638 2554 3642
rect 2702 3618 2706 3622
rect 2558 3608 2562 3612
rect 2614 3608 2618 3612
rect 2550 3528 2554 3532
rect 2534 3518 2538 3522
rect 2550 3518 2554 3522
rect 2534 3488 2538 3492
rect 2526 3468 2530 3472
rect 2526 3458 2530 3462
rect 2518 3368 2522 3372
rect 2586 3603 2590 3607
rect 2593 3603 2597 3607
rect 2598 3588 2602 3592
rect 2582 3568 2586 3572
rect 2566 3528 2570 3532
rect 2694 3578 2698 3582
rect 2622 3548 2626 3552
rect 2662 3548 2666 3552
rect 2694 3548 2698 3552
rect 2638 3538 2642 3542
rect 2662 3538 2666 3542
rect 2646 3528 2650 3532
rect 2630 3518 2634 3522
rect 2654 3518 2658 3522
rect 2622 3488 2626 3492
rect 2630 3488 2634 3492
rect 2630 3468 2634 3472
rect 2614 3448 2618 3452
rect 2630 3448 2634 3452
rect 2646 3448 2650 3452
rect 2566 3438 2570 3442
rect 2586 3403 2590 3407
rect 2593 3403 2597 3407
rect 2550 3398 2554 3402
rect 2606 3388 2610 3392
rect 2534 3368 2538 3372
rect 2542 3368 2546 3372
rect 2558 3368 2562 3372
rect 2550 3358 2554 3362
rect 2526 3348 2530 3352
rect 2534 3348 2538 3352
rect 2526 3328 2530 3332
rect 2654 3438 2658 3442
rect 2614 3368 2618 3372
rect 2614 3358 2618 3362
rect 2566 3328 2570 3332
rect 2550 3288 2554 3292
rect 2566 3288 2570 3292
rect 2542 3248 2546 3252
rect 2534 3228 2538 3232
rect 2558 3188 2562 3192
rect 2518 3168 2522 3172
rect 2582 3278 2586 3282
rect 2614 3268 2618 3272
rect 2574 3258 2578 3262
rect 2630 3258 2634 3262
rect 2598 3248 2602 3252
rect 2622 3248 2626 3252
rect 2586 3203 2590 3207
rect 2593 3203 2597 3207
rect 2654 3268 2658 3272
rect 2654 3258 2658 3262
rect 2614 3168 2618 3172
rect 2638 3168 2642 3172
rect 2542 3148 2546 3152
rect 2566 3148 2570 3152
rect 2606 3148 2610 3152
rect 2518 3118 2522 3122
rect 2510 3108 2514 3112
rect 2534 3138 2538 3142
rect 2550 3138 2554 3142
rect 2526 3078 2530 3082
rect 2630 3138 2634 3142
rect 2654 3128 2658 3132
rect 2638 3118 2642 3122
rect 2574 3088 2578 3092
rect 2470 3068 2474 3072
rect 2502 3068 2506 3072
rect 2566 3078 2570 3082
rect 2614 3078 2618 3082
rect 2558 3068 2562 3072
rect 2582 3068 2586 3072
rect 2494 3058 2498 3062
rect 2510 3058 2514 3062
rect 2542 3058 2546 3062
rect 2414 3038 2418 3042
rect 2430 3038 2434 3042
rect 2462 3008 2466 3012
rect 2406 2998 2410 3002
rect 2422 2998 2426 3002
rect 2382 2958 2386 2962
rect 2422 2978 2426 2982
rect 2406 2948 2410 2952
rect 2342 2928 2346 2932
rect 2502 3038 2506 3042
rect 2526 3028 2530 3032
rect 2494 2978 2498 2982
rect 2470 2968 2474 2972
rect 2486 2968 2490 2972
rect 2494 2958 2498 2962
rect 2486 2948 2490 2952
rect 2518 2948 2522 2952
rect 2446 2938 2450 2942
rect 2502 2918 2506 2922
rect 2518 2908 2522 2912
rect 2486 2898 2490 2902
rect 2414 2868 2418 2872
rect 2422 2868 2426 2872
rect 2446 2868 2450 2872
rect 2470 2868 2474 2872
rect 2510 2868 2514 2872
rect 2334 2808 2338 2812
rect 2382 2848 2386 2852
rect 2430 2848 2434 2852
rect 2462 2848 2466 2852
rect 2302 2778 2306 2782
rect 2350 2778 2354 2782
rect 2470 2818 2474 2822
rect 2446 2768 2450 2772
rect 2550 3028 2554 3032
rect 2542 2968 2546 2972
rect 2670 3528 2674 3532
rect 2766 3738 2770 3742
rect 2782 3728 2786 3732
rect 2750 3678 2754 3682
rect 2846 3878 2850 3882
rect 2806 3698 2810 3702
rect 2838 3808 2842 3812
rect 2830 3788 2834 3792
rect 2822 3748 2826 3752
rect 2822 3698 2826 3702
rect 2814 3688 2818 3692
rect 2790 3678 2794 3682
rect 2782 3668 2786 3672
rect 2862 3918 2866 3922
rect 2854 3758 2858 3762
rect 2854 3738 2858 3742
rect 2862 3738 2866 3742
rect 2918 3968 2922 3972
rect 2982 3898 2986 3902
rect 2950 3878 2954 3882
rect 2918 3868 2922 3872
rect 2958 3868 2962 3872
rect 2974 3868 2978 3872
rect 2878 3778 2882 3782
rect 2950 3858 2954 3862
rect 3062 4008 3066 4012
rect 3118 4008 3122 4012
rect 3038 3958 3042 3962
rect 3070 3948 3074 3952
rect 3006 3918 3010 3922
rect 3046 3928 3050 3932
rect 3014 3908 3018 3912
rect 3014 3878 3018 3882
rect 2998 3868 3002 3872
rect 2990 3858 2994 3862
rect 3006 3858 3010 3862
rect 2990 3848 2994 3852
rect 3038 3868 3042 3872
rect 3062 3868 3066 3872
rect 3182 4118 3186 4122
rect 3142 4108 3146 4112
rect 3198 4108 3202 4112
rect 3254 4148 3258 4152
rect 3246 4138 3250 4142
rect 3270 4128 3274 4132
rect 3206 4098 3210 4102
rect 3214 4088 3218 4092
rect 3158 4068 3162 4072
rect 3246 4068 3250 4072
rect 3182 4058 3186 4062
rect 3214 4008 3218 4012
rect 3182 3948 3186 3952
rect 3246 3948 3250 3952
rect 3094 3918 3098 3922
rect 3134 3918 3138 3922
rect 3098 3903 3102 3907
rect 3105 3903 3109 3907
rect 3142 3898 3146 3902
rect 3254 3918 3258 3922
rect 3238 3898 3242 3902
rect 3222 3868 3226 3872
rect 3254 3868 3258 3872
rect 3294 4348 3298 4352
rect 3366 4338 3370 4342
rect 3310 4288 3314 4292
rect 3310 4278 3314 4282
rect 3310 4268 3314 4272
rect 3334 4298 3338 4302
rect 3438 4368 3442 4372
rect 3438 4358 3442 4362
rect 3446 4358 3450 4362
rect 3414 4348 3418 4352
rect 3462 4368 3466 4372
rect 3534 4558 3538 4562
rect 3510 4548 3514 4552
rect 3518 4548 3522 4552
rect 3534 4538 3538 4542
rect 3614 4618 3618 4622
rect 3646 4618 3650 4622
rect 3610 4603 3614 4607
rect 3617 4603 3621 4607
rect 3566 4558 3570 4562
rect 3590 4547 3594 4551
rect 3630 4548 3634 4552
rect 3750 4718 3754 4722
rect 3862 4748 3866 4752
rect 3838 4738 3842 4742
rect 3686 4668 3690 4672
rect 3726 4668 3730 4672
rect 3798 4668 3802 4672
rect 3670 4658 3674 4662
rect 3670 4648 3674 4652
rect 3662 4638 3666 4642
rect 3686 4588 3690 4592
rect 3734 4588 3738 4592
rect 3686 4558 3690 4562
rect 3534 4508 3538 4512
rect 3542 4508 3546 4512
rect 3606 4498 3610 4502
rect 3534 4488 3538 4492
rect 3590 4468 3594 4472
rect 3542 4458 3546 4462
rect 3566 4458 3570 4462
rect 3502 4448 3506 4452
rect 3534 4438 3538 4442
rect 3542 4428 3546 4432
rect 3526 4398 3530 4402
rect 3558 4448 3562 4452
rect 3590 4448 3594 4452
rect 3598 4448 3602 4452
rect 3550 4388 3554 4392
rect 3494 4378 3498 4382
rect 3550 4358 3554 4362
rect 3470 4348 3474 4352
rect 3502 4348 3506 4352
rect 3550 4348 3554 4352
rect 3398 4338 3402 4342
rect 3462 4338 3466 4342
rect 3478 4338 3482 4342
rect 3486 4328 3490 4332
rect 3502 4318 3506 4322
rect 3422 4278 3426 4282
rect 3454 4278 3458 4282
rect 3350 4268 3354 4272
rect 3342 4258 3346 4262
rect 3326 4248 3330 4252
rect 3342 4248 3346 4252
rect 3286 4188 3290 4192
rect 3302 4168 3306 4172
rect 3366 4238 3370 4242
rect 3398 4158 3402 4162
rect 3470 4268 3474 4272
rect 3478 4258 3482 4262
rect 3510 4288 3514 4292
rect 3510 4268 3514 4272
rect 3610 4403 3614 4407
rect 3617 4403 3621 4407
rect 3622 4378 3626 4382
rect 3718 4548 3722 4552
rect 3662 4538 3666 4542
rect 3670 4528 3674 4532
rect 3662 4438 3666 4442
rect 3798 4648 3802 4652
rect 3886 4728 3890 4732
rect 3878 4718 3882 4722
rect 3838 4708 3842 4712
rect 3822 4698 3826 4702
rect 3830 4698 3834 4702
rect 3878 4688 3882 4692
rect 3974 4758 3978 4762
rect 4070 4758 4074 4762
rect 3942 4748 3946 4752
rect 3926 4738 3930 4742
rect 3830 4678 3834 4682
rect 3910 4678 3914 4682
rect 3894 4668 3898 4672
rect 3878 4648 3882 4652
rect 3782 4638 3786 4642
rect 3814 4638 3818 4642
rect 3870 4628 3874 4632
rect 3806 4618 3810 4622
rect 3758 4548 3762 4552
rect 3766 4508 3770 4512
rect 3790 4508 3794 4512
rect 3766 4488 3770 4492
rect 3782 4488 3786 4492
rect 3782 4468 3786 4472
rect 3726 4458 3730 4462
rect 3678 4438 3682 4442
rect 3686 4388 3690 4392
rect 3670 4348 3674 4352
rect 3598 4338 3602 4342
rect 3590 4308 3594 4312
rect 3582 4278 3586 4282
rect 3606 4288 3610 4292
rect 3534 4268 3538 4272
rect 3558 4268 3562 4272
rect 3574 4268 3578 4272
rect 3582 4268 3586 4272
rect 3598 4268 3602 4272
rect 3478 4248 3482 4252
rect 3526 4248 3530 4252
rect 3566 4248 3570 4252
rect 3646 4318 3650 4322
rect 3598 4258 3602 4262
rect 3654 4258 3658 4262
rect 3630 4248 3634 4252
rect 3446 4218 3450 4222
rect 3462 4218 3466 4222
rect 3422 4178 3426 4182
rect 3414 4168 3418 4172
rect 3438 4168 3442 4172
rect 3526 4228 3530 4232
rect 3438 4148 3442 4152
rect 3326 4138 3330 4142
rect 3390 4128 3394 4132
rect 3358 4098 3362 4102
rect 3390 4108 3394 4112
rect 3334 4088 3338 4092
rect 3470 4148 3474 4152
rect 3454 4138 3458 4142
rect 3462 4138 3466 4142
rect 3446 4118 3450 4122
rect 3406 4088 3410 4092
rect 3446 4088 3450 4092
rect 3486 4138 3490 4142
rect 3478 4118 3482 4122
rect 3470 4108 3474 4112
rect 3374 4068 3378 4072
rect 3390 4068 3394 4072
rect 3406 4068 3410 4072
rect 3454 4068 3458 4072
rect 3278 4058 3282 4062
rect 3310 4048 3314 4052
rect 3334 4048 3338 4052
rect 3342 4008 3346 4012
rect 3366 4008 3370 4012
rect 3286 3998 3290 4002
rect 3270 3948 3274 3952
rect 3270 3878 3274 3882
rect 3270 3868 3274 3872
rect 3382 4058 3386 4062
rect 3390 4048 3394 4052
rect 3486 4068 3490 4072
rect 3502 4068 3506 4072
rect 3470 4048 3474 4052
rect 3414 4018 3418 4022
rect 3390 3988 3394 3992
rect 3430 3988 3434 3992
rect 3342 3958 3346 3962
rect 3406 3968 3410 3972
rect 3558 4218 3562 4222
rect 3534 4098 3538 4102
rect 3582 4208 3586 4212
rect 3630 4208 3634 4212
rect 3566 4148 3570 4152
rect 3610 4203 3614 4207
rect 3617 4203 3621 4207
rect 3582 4138 3586 4142
rect 3606 4138 3610 4142
rect 3654 4248 3658 4252
rect 3662 4248 3666 4252
rect 3646 4218 3650 4222
rect 3638 4178 3642 4182
rect 3646 4168 3650 4172
rect 3718 4268 3722 4272
rect 3694 4158 3698 4162
rect 3758 4458 3762 4462
rect 3742 4448 3746 4452
rect 3870 4598 3874 4602
rect 3814 4548 3818 4552
rect 3822 4508 3826 4512
rect 3798 4468 3802 4472
rect 3742 4398 3746 4402
rect 3758 4378 3762 4382
rect 3806 4428 3810 4432
rect 3798 4368 3802 4372
rect 3774 4348 3778 4352
rect 3782 4338 3786 4342
rect 3782 4278 3786 4282
rect 3790 4278 3794 4282
rect 3806 4278 3810 4282
rect 3758 4268 3762 4272
rect 3750 4258 3754 4262
rect 3766 4248 3770 4252
rect 3798 4258 3802 4262
rect 3790 4238 3794 4242
rect 3774 4198 3778 4202
rect 3790 4178 3794 4182
rect 3790 4168 3794 4172
rect 3750 4158 3754 4162
rect 3766 4148 3770 4152
rect 3742 4138 3746 4142
rect 3758 4138 3762 4142
rect 3782 4138 3786 4142
rect 3590 4118 3594 4122
rect 3630 4118 3634 4122
rect 3550 4068 3554 4072
rect 3542 4058 3546 4062
rect 3662 4108 3666 4112
rect 3638 4098 3642 4102
rect 3566 4088 3570 4092
rect 3574 4088 3578 4092
rect 3734 4108 3738 4112
rect 3742 4088 3746 4092
rect 3574 4068 3578 4072
rect 3686 4068 3690 4072
rect 3726 4068 3730 4072
rect 3654 4058 3658 4062
rect 3678 4058 3682 4062
rect 3550 4048 3554 4052
rect 3518 4038 3522 4042
rect 3518 4018 3522 4022
rect 3542 3998 3546 4002
rect 3510 3968 3514 3972
rect 3486 3958 3490 3962
rect 3246 3858 3250 3862
rect 3054 3848 3058 3852
rect 3070 3848 3074 3852
rect 3022 3828 3026 3832
rect 3086 3828 3090 3832
rect 3014 3768 3018 3772
rect 3022 3768 3026 3772
rect 2894 3758 2898 3762
rect 2910 3758 2914 3762
rect 2878 3748 2882 3752
rect 2918 3748 2922 3752
rect 2998 3748 3002 3752
rect 3110 3748 3114 3752
rect 3126 3748 3130 3752
rect 2894 3738 2898 3742
rect 2974 3738 2978 3742
rect 3078 3738 3082 3742
rect 2870 3718 2874 3722
rect 2894 3698 2898 3702
rect 3098 3703 3102 3707
rect 3105 3703 3109 3707
rect 3014 3698 3018 3702
rect 3102 3688 3106 3692
rect 3102 3678 3106 3682
rect 2910 3668 2914 3672
rect 2950 3668 2954 3672
rect 3094 3668 3098 3672
rect 2726 3598 2730 3602
rect 2710 3588 2714 3592
rect 2726 3578 2730 3582
rect 2790 3658 2794 3662
rect 2902 3658 2906 3662
rect 2958 3658 2962 3662
rect 2998 3659 3002 3663
rect 3070 3658 3074 3662
rect 2774 3648 2778 3652
rect 2734 3568 2738 3572
rect 2790 3568 2794 3572
rect 2766 3547 2770 3551
rect 2710 3518 2714 3522
rect 2678 3498 2682 3502
rect 2710 3488 2714 3492
rect 2830 3578 2834 3582
rect 2886 3578 2890 3582
rect 2838 3568 2842 3572
rect 2862 3548 2866 3552
rect 2830 3528 2834 3532
rect 2822 3498 2826 3502
rect 2814 3488 2818 3492
rect 2726 3478 2730 3482
rect 2790 3478 2794 3482
rect 2670 3468 2674 3472
rect 2678 3458 2682 3462
rect 2774 3448 2778 3452
rect 2710 3438 2714 3442
rect 2670 3428 2674 3432
rect 2758 3358 2762 3362
rect 2678 3348 2682 3352
rect 2678 3298 2682 3302
rect 2782 3428 2786 3432
rect 2750 3288 2754 3292
rect 2774 3288 2778 3292
rect 2734 3268 2738 3272
rect 2886 3538 2890 3542
rect 2870 3518 2874 3522
rect 2862 3508 2866 3512
rect 2894 3498 2898 3502
rect 2894 3468 2898 3472
rect 2870 3458 2874 3462
rect 2886 3448 2890 3452
rect 2838 3418 2842 3422
rect 2878 3418 2882 3422
rect 2870 3408 2874 3412
rect 2822 3368 2826 3372
rect 2854 3368 2858 3372
rect 2838 3358 2842 3362
rect 2862 3358 2866 3362
rect 2886 3358 2890 3362
rect 2830 3348 2834 3352
rect 2814 3338 2818 3342
rect 2798 3318 2802 3322
rect 2822 3308 2826 3312
rect 2694 3258 2698 3262
rect 2774 3258 2778 3262
rect 2798 3258 2802 3262
rect 2742 3248 2746 3252
rect 2766 3248 2770 3252
rect 2670 3238 2674 3242
rect 2758 3238 2762 3242
rect 2750 3218 2754 3222
rect 2718 3198 2722 3202
rect 2822 3248 2826 3252
rect 2782 3208 2786 3212
rect 2774 3198 2778 3202
rect 2726 3188 2730 3192
rect 2694 3148 2698 3152
rect 2806 3178 2810 3182
rect 2822 3178 2826 3182
rect 2878 3328 2882 3332
rect 2862 3298 2866 3302
rect 2886 3268 2890 3272
rect 2934 3648 2938 3652
rect 2934 3568 2938 3572
rect 2926 3547 2930 3551
rect 3046 3648 3050 3652
rect 3062 3638 3066 3642
rect 2990 3588 2994 3592
rect 3038 3588 3042 3592
rect 2974 3578 2978 3582
rect 2974 3568 2978 3572
rect 2942 3528 2946 3532
rect 2942 3518 2946 3522
rect 3006 3578 3010 3582
rect 3078 3628 3082 3632
rect 3030 3548 3034 3552
rect 3054 3548 3058 3552
rect 3086 3548 3090 3552
rect 3006 3538 3010 3542
rect 3038 3538 3042 3542
rect 3046 3538 3050 3542
rect 3022 3508 3026 3512
rect 3046 3478 3050 3482
rect 3054 3468 3058 3472
rect 2990 3458 2994 3462
rect 2926 3448 2930 3452
rect 2910 3418 2914 3422
rect 2902 3408 2906 3412
rect 3046 3438 3050 3442
rect 2942 3418 2946 3422
rect 2926 3368 2930 3372
rect 3054 3408 3058 3412
rect 2958 3378 2962 3382
rect 2934 3348 2938 3352
rect 2990 3368 2994 3372
rect 3046 3368 3050 3372
rect 2910 3338 2914 3342
rect 2974 3338 2978 3342
rect 2910 3288 2914 3292
rect 2902 3268 2906 3272
rect 2934 3268 2938 3272
rect 2846 3258 2850 3262
rect 2894 3248 2898 3252
rect 2910 3248 2914 3252
rect 2854 3198 2858 3202
rect 2790 3168 2794 3172
rect 2838 3168 2842 3172
rect 2766 3158 2770 3162
rect 2678 3128 2682 3132
rect 2662 3098 2666 3102
rect 2574 3048 2578 3052
rect 2598 3048 2602 3052
rect 2614 3008 2618 3012
rect 2586 3003 2590 3007
rect 2593 3003 2597 3007
rect 2574 2998 2578 3002
rect 2574 2968 2578 2972
rect 2630 2968 2634 2972
rect 2798 3148 2802 3152
rect 2758 3138 2762 3142
rect 2742 3108 2746 3112
rect 2806 3138 2810 3142
rect 2798 3118 2802 3122
rect 2718 3098 2722 3102
rect 2774 3098 2778 3102
rect 2710 3078 2714 3082
rect 2694 3058 2698 3062
rect 2710 3048 2714 3052
rect 2686 2968 2690 2972
rect 2710 2968 2714 2972
rect 2558 2948 2562 2952
rect 2622 2948 2626 2952
rect 2590 2938 2594 2942
rect 2542 2928 2546 2932
rect 2558 2868 2562 2872
rect 2502 2838 2506 2842
rect 2518 2838 2522 2842
rect 2526 2808 2530 2812
rect 2526 2788 2530 2792
rect 2358 2758 2362 2762
rect 2430 2758 2434 2762
rect 2486 2758 2490 2762
rect 2534 2758 2538 2762
rect 2598 2898 2602 2902
rect 2614 2928 2618 2932
rect 2606 2838 2610 2842
rect 2586 2803 2590 2807
rect 2593 2803 2597 2807
rect 2606 2768 2610 2772
rect 2334 2748 2338 2752
rect 2390 2748 2394 2752
rect 2542 2748 2546 2752
rect 2558 2748 2562 2752
rect 2606 2748 2610 2752
rect 2310 2738 2314 2742
rect 2334 2728 2338 2732
rect 2302 2668 2306 2672
rect 2150 2658 2154 2662
rect 2166 2658 2170 2662
rect 2222 2658 2226 2662
rect 2270 2658 2274 2662
rect 2262 2648 2266 2652
rect 2302 2648 2306 2652
rect 2102 2548 2106 2552
rect 2142 2548 2146 2552
rect 2158 2548 2162 2552
rect 2062 2508 2066 2512
rect 2074 2503 2078 2507
rect 2081 2503 2085 2507
rect 2110 2518 2114 2522
rect 2102 2508 2106 2512
rect 2134 2528 2138 2532
rect 2158 2518 2162 2522
rect 2118 2488 2122 2492
rect 2062 2478 2066 2482
rect 2094 2478 2098 2482
rect 2166 2508 2170 2512
rect 2198 2508 2202 2512
rect 2246 2628 2250 2632
rect 2270 2598 2274 2602
rect 2294 2598 2298 2602
rect 2238 2578 2242 2582
rect 2214 2528 2218 2532
rect 2214 2518 2218 2522
rect 2206 2498 2210 2502
rect 2302 2588 2306 2592
rect 2294 2548 2298 2552
rect 2382 2738 2386 2742
rect 2430 2728 2434 2732
rect 2350 2718 2354 2722
rect 2366 2698 2370 2702
rect 2422 2698 2426 2702
rect 2430 2698 2434 2702
rect 2358 2668 2362 2672
rect 2382 2668 2386 2672
rect 2414 2668 2418 2672
rect 2478 2738 2482 2742
rect 2566 2728 2570 2732
rect 2558 2718 2562 2722
rect 2478 2698 2482 2702
rect 2526 2698 2530 2702
rect 2542 2698 2546 2702
rect 2462 2668 2466 2672
rect 2350 2658 2354 2662
rect 2374 2658 2378 2662
rect 2406 2648 2410 2652
rect 2406 2628 2410 2632
rect 2374 2618 2378 2622
rect 2366 2588 2370 2592
rect 2318 2558 2322 2562
rect 2334 2558 2338 2562
rect 2262 2538 2266 2542
rect 2238 2518 2242 2522
rect 2262 2518 2266 2522
rect 2238 2498 2242 2502
rect 2222 2488 2226 2492
rect 2246 2478 2250 2482
rect 2254 2468 2258 2472
rect 2030 2448 2034 2452
rect 2014 2368 2018 2372
rect 2118 2458 2122 2462
rect 2126 2458 2130 2462
rect 2166 2458 2170 2462
rect 2070 2448 2074 2452
rect 2070 2438 2074 2442
rect 2046 2358 2050 2362
rect 2062 2358 2066 2362
rect 2014 2348 2018 2352
rect 2006 2338 2010 2342
rect 2038 2338 2042 2342
rect 1974 2328 1978 2332
rect 2030 2328 2034 2332
rect 2022 2318 2026 2322
rect 1990 2308 1994 2312
rect 2006 2308 2010 2312
rect 1998 2288 2002 2292
rect 2014 2278 2018 2282
rect 1942 2268 1946 2272
rect 1998 2268 2002 2272
rect 1886 2258 1890 2262
rect 1870 2218 1874 2222
rect 1934 2218 1938 2222
rect 1966 2218 1970 2222
rect 1910 2208 1914 2212
rect 1934 2208 1938 2212
rect 1862 2198 1866 2202
rect 1878 2198 1882 2202
rect 1926 2198 1930 2202
rect 1862 2158 1866 2162
rect 1830 2138 1834 2142
rect 1846 2138 1850 2142
rect 1814 2128 1818 2132
rect 1846 2098 1850 2102
rect 1870 2088 1874 2092
rect 1902 2168 1906 2172
rect 1950 2198 1954 2202
rect 1918 2158 1922 2162
rect 1886 2118 1890 2122
rect 1894 2108 1898 2112
rect 1958 2178 1962 2182
rect 1958 2158 1962 2162
rect 1918 2138 1922 2142
rect 1990 2188 1994 2192
rect 1990 2168 1994 2172
rect 1974 2148 1978 2152
rect 1990 2148 1994 2152
rect 2014 2248 2018 2252
rect 2006 2218 2010 2222
rect 2014 2218 2018 2222
rect 2014 2178 2018 2182
rect 2022 2158 2026 2162
rect 1934 2138 1938 2142
rect 1966 2138 1970 2142
rect 1998 2138 2002 2142
rect 1926 2108 1930 2112
rect 1902 2098 1906 2102
rect 1758 2058 1762 2062
rect 1830 2058 1834 2062
rect 1878 2058 1882 2062
rect 1774 2028 1778 2032
rect 1758 1998 1762 2002
rect 1750 1988 1754 1992
rect 1838 2048 1842 2052
rect 1854 2048 1858 2052
rect 1806 2028 1810 2032
rect 1790 2008 1794 2012
rect 1782 1998 1786 2002
rect 1774 1978 1778 1982
rect 1734 1958 1738 1962
rect 1718 1888 1722 1892
rect 1742 1868 1746 1872
rect 1758 1938 1762 1942
rect 1782 1938 1786 1942
rect 1766 1908 1770 1912
rect 1862 2018 1866 2022
rect 1862 1958 1866 1962
rect 1814 1868 1818 1872
rect 1830 1868 1834 1872
rect 1734 1858 1738 1862
rect 1750 1858 1754 1862
rect 1766 1858 1770 1862
rect 1814 1858 1818 1862
rect 1782 1848 1786 1852
rect 1718 1778 1722 1782
rect 1726 1778 1730 1782
rect 1758 1788 1762 1792
rect 1750 1758 1754 1762
rect 1718 1738 1722 1742
rect 1702 1728 1706 1732
rect 1734 1738 1738 1742
rect 1750 1748 1754 1752
rect 1726 1718 1730 1722
rect 1742 1718 1746 1722
rect 1742 1698 1746 1702
rect 1678 1668 1682 1672
rect 1678 1658 1682 1662
rect 1774 1758 1778 1762
rect 1790 1758 1794 1762
rect 1774 1748 1778 1752
rect 1726 1658 1730 1662
rect 1766 1658 1770 1662
rect 1702 1648 1706 1652
rect 1734 1648 1738 1652
rect 1750 1648 1754 1652
rect 1694 1628 1698 1632
rect 1718 1628 1722 1632
rect 1694 1598 1698 1602
rect 1678 1558 1682 1562
rect 1806 1728 1810 1732
rect 1798 1708 1802 1712
rect 1862 1938 1866 1942
rect 1846 1928 1850 1932
rect 1862 1908 1866 1912
rect 1878 1908 1882 1912
rect 1854 1868 1858 1872
rect 1862 1868 1866 1872
rect 1838 1858 1842 1862
rect 1838 1848 1842 1852
rect 1822 1688 1826 1692
rect 1806 1658 1810 1662
rect 1790 1628 1794 1632
rect 1758 1598 1762 1602
rect 1774 1598 1778 1602
rect 1790 1578 1794 1582
rect 1702 1558 1706 1562
rect 1830 1588 1834 1592
rect 1798 1558 1802 1562
rect 1926 2078 1930 2082
rect 1942 2128 1946 2132
rect 1958 2128 1962 2132
rect 2014 2128 2018 2132
rect 1990 2108 1994 2112
rect 1910 2018 1914 2022
rect 1902 1978 1906 1982
rect 1910 1968 1914 1972
rect 1918 1968 1922 1972
rect 1902 1958 1906 1962
rect 1894 1948 1898 1952
rect 1902 1928 1906 1932
rect 1910 1928 1914 1932
rect 1902 1898 1906 1902
rect 1926 1858 1930 1862
rect 1902 1848 1906 1852
rect 1910 1848 1914 1852
rect 1974 2018 1978 2022
rect 2022 2008 2026 2012
rect 2054 2328 2058 2332
rect 2038 2268 2042 2272
rect 2054 2288 2058 2292
rect 2070 2348 2074 2352
rect 2150 2438 2154 2442
rect 2110 2428 2114 2432
rect 2166 2438 2170 2442
rect 2158 2418 2162 2422
rect 2150 2408 2154 2412
rect 2134 2388 2138 2392
rect 2118 2368 2122 2372
rect 2094 2338 2098 2342
rect 2110 2338 2114 2342
rect 2078 2328 2082 2332
rect 2094 2328 2098 2332
rect 2102 2328 2106 2332
rect 2074 2303 2078 2307
rect 2081 2303 2085 2307
rect 2046 2258 2050 2262
rect 2054 2248 2058 2252
rect 2062 2248 2066 2252
rect 2070 2198 2074 2202
rect 2062 2188 2066 2192
rect 2046 2178 2050 2182
rect 2054 2178 2058 2182
rect 2062 2148 2066 2152
rect 2054 2138 2058 2142
rect 2046 2098 2050 2102
rect 2078 2148 2082 2152
rect 2086 2148 2090 2152
rect 2142 2368 2146 2372
rect 2158 2398 2162 2402
rect 2134 2308 2138 2312
rect 2126 2268 2130 2272
rect 2118 2248 2122 2252
rect 2110 2218 2114 2222
rect 2102 2198 2106 2202
rect 2118 2168 2122 2172
rect 2134 2228 2138 2232
rect 2230 2458 2234 2462
rect 2182 2418 2186 2422
rect 2174 2388 2178 2392
rect 2174 2348 2178 2352
rect 2206 2448 2210 2452
rect 2222 2448 2226 2452
rect 2214 2378 2218 2382
rect 2230 2348 2234 2352
rect 2278 2538 2282 2542
rect 2278 2518 2282 2522
rect 2302 2508 2306 2512
rect 2358 2548 2362 2552
rect 2334 2528 2338 2532
rect 2302 2478 2306 2482
rect 2342 2478 2346 2482
rect 2462 2608 2466 2612
rect 2390 2588 2394 2592
rect 2382 2558 2386 2562
rect 2398 2578 2402 2582
rect 2414 2558 2418 2562
rect 2438 2558 2442 2562
rect 2454 2558 2458 2562
rect 2366 2528 2370 2532
rect 2438 2518 2442 2522
rect 2446 2498 2450 2502
rect 2422 2478 2426 2482
rect 2430 2478 2434 2482
rect 2278 2468 2282 2472
rect 2366 2468 2370 2472
rect 2390 2468 2394 2472
rect 2406 2468 2410 2472
rect 2318 2458 2322 2462
rect 2358 2458 2362 2462
rect 2382 2458 2386 2462
rect 2430 2458 2434 2462
rect 2310 2448 2314 2452
rect 2294 2438 2298 2442
rect 2302 2438 2306 2442
rect 2294 2428 2298 2432
rect 2278 2408 2282 2412
rect 2286 2378 2290 2382
rect 2278 2358 2282 2362
rect 2262 2348 2266 2352
rect 2182 2328 2186 2332
rect 2198 2328 2202 2332
rect 2206 2328 2210 2332
rect 2190 2318 2194 2322
rect 2166 2308 2170 2312
rect 2198 2278 2202 2282
rect 2174 2268 2178 2272
rect 2286 2328 2290 2332
rect 2334 2448 2338 2452
rect 2326 2438 2330 2442
rect 2366 2438 2370 2442
rect 2334 2368 2338 2372
rect 2358 2368 2362 2372
rect 2342 2358 2346 2362
rect 2326 2348 2330 2352
rect 2318 2338 2322 2342
rect 2286 2308 2290 2312
rect 2302 2308 2306 2312
rect 2310 2288 2314 2292
rect 2358 2348 2362 2352
rect 2438 2448 2442 2452
rect 2534 2678 2538 2682
rect 2558 2678 2562 2682
rect 2526 2648 2530 2652
rect 2534 2618 2538 2622
rect 2502 2578 2506 2582
rect 2494 2488 2498 2492
rect 2462 2468 2466 2472
rect 2462 2458 2466 2462
rect 2486 2458 2490 2462
rect 2382 2428 2386 2432
rect 2430 2428 2434 2432
rect 2382 2358 2386 2362
rect 2414 2348 2418 2352
rect 2366 2338 2370 2342
rect 2358 2308 2362 2312
rect 2230 2278 2234 2282
rect 2262 2278 2266 2282
rect 2326 2278 2330 2282
rect 2238 2268 2242 2272
rect 2278 2268 2282 2272
rect 2302 2268 2306 2272
rect 2150 2258 2154 2262
rect 2214 2258 2218 2262
rect 2158 2248 2162 2252
rect 2142 2218 2146 2222
rect 2142 2158 2146 2162
rect 2110 2138 2114 2142
rect 2142 2138 2146 2142
rect 2062 2118 2066 2122
rect 2102 2128 2106 2132
rect 2054 2068 2058 2072
rect 2074 2103 2078 2107
rect 2081 2103 2085 2107
rect 2126 2128 2130 2132
rect 2206 2198 2210 2202
rect 2182 2178 2186 2182
rect 2198 2168 2202 2172
rect 2174 2158 2178 2162
rect 2182 2148 2186 2152
rect 2206 2138 2210 2142
rect 2254 2238 2258 2242
rect 2318 2248 2322 2252
rect 2350 2248 2354 2252
rect 2302 2228 2306 2232
rect 2230 2208 2234 2212
rect 2350 2218 2354 2222
rect 2294 2168 2298 2172
rect 2350 2158 2354 2162
rect 2110 2108 2114 2112
rect 2118 2068 2122 2072
rect 2086 2048 2090 2052
rect 2038 2018 2042 2022
rect 1974 1998 1978 2002
rect 1990 1998 1994 2002
rect 2014 1998 2018 2002
rect 1950 1958 1954 1962
rect 2134 2008 2138 2012
rect 2142 2008 2146 2012
rect 2110 1998 2114 2002
rect 2118 1998 2122 2002
rect 2054 1978 2058 1982
rect 2006 1968 2010 1972
rect 2022 1958 2026 1962
rect 2062 1948 2066 1952
rect 2086 1948 2090 1952
rect 1942 1858 1946 1862
rect 1894 1828 1898 1832
rect 1894 1808 1898 1812
rect 1886 1798 1890 1802
rect 1926 1828 1930 1832
rect 1934 1828 1938 1832
rect 1934 1798 1938 1802
rect 1958 1798 1962 1802
rect 1902 1778 1906 1782
rect 1958 1778 1962 1782
rect 1878 1768 1882 1772
rect 1862 1758 1866 1762
rect 1870 1758 1874 1762
rect 1862 1688 1866 1692
rect 1870 1688 1874 1692
rect 1918 1758 1922 1762
rect 1918 1738 1922 1742
rect 1926 1728 1930 1732
rect 1950 1708 1954 1712
rect 1870 1658 1874 1662
rect 1894 1658 1898 1662
rect 1926 1658 1930 1662
rect 1934 1648 1938 1652
rect 1878 1628 1882 1632
rect 1894 1628 1898 1632
rect 1670 1548 1674 1552
rect 1686 1548 1690 1552
rect 1742 1548 1746 1552
rect 1798 1548 1802 1552
rect 1846 1548 1850 1552
rect 1662 1538 1666 1542
rect 1638 1508 1642 1512
rect 1670 1508 1674 1512
rect 1622 1438 1626 1442
rect 1694 1528 1698 1532
rect 1702 1488 1706 1492
rect 1686 1468 1690 1472
rect 1734 1488 1738 1492
rect 1678 1438 1682 1442
rect 1638 1398 1642 1402
rect 1670 1378 1674 1382
rect 1702 1428 1706 1432
rect 1694 1368 1698 1372
rect 1582 1358 1586 1362
rect 1662 1358 1666 1362
rect 1750 1448 1754 1452
rect 1782 1538 1786 1542
rect 1846 1508 1850 1512
rect 1806 1498 1810 1502
rect 1814 1488 1818 1492
rect 1790 1468 1794 1472
rect 1766 1458 1770 1462
rect 1758 1438 1762 1442
rect 1814 1448 1818 1452
rect 1846 1448 1850 1452
rect 1822 1438 1826 1442
rect 1790 1428 1794 1432
rect 1758 1408 1762 1412
rect 1726 1398 1730 1402
rect 1742 1398 1746 1402
rect 1710 1378 1714 1382
rect 1710 1358 1714 1362
rect 1838 1368 1842 1372
rect 1830 1358 1834 1362
rect 1598 1348 1602 1352
rect 1630 1348 1634 1352
rect 1774 1348 1778 1352
rect 1790 1348 1794 1352
rect 1830 1348 1834 1352
rect 1550 1338 1554 1342
rect 1566 1338 1570 1342
rect 1550 1318 1554 1322
rect 1614 1298 1618 1302
rect 1574 1288 1578 1292
rect 1630 1288 1634 1292
rect 1542 1268 1546 1272
rect 1606 1268 1610 1272
rect 1398 1238 1402 1242
rect 1422 1238 1426 1242
rect 1438 1238 1442 1242
rect 1494 1238 1498 1242
rect 1454 1208 1458 1212
rect 1494 1198 1498 1202
rect 1390 1188 1394 1192
rect 1518 1188 1522 1192
rect 1470 1178 1474 1182
rect 1510 1178 1514 1182
rect 1422 1158 1426 1162
rect 1454 1158 1458 1162
rect 1382 1148 1386 1152
rect 1430 1148 1434 1152
rect 1438 1148 1442 1152
rect 1350 1128 1354 1132
rect 1406 1128 1410 1132
rect 1310 1058 1314 1062
rect 1222 978 1226 982
rect 1214 968 1218 972
rect 1198 938 1202 942
rect 1190 928 1194 932
rect 1166 918 1170 922
rect 1182 918 1186 922
rect 1166 878 1170 882
rect 1190 908 1194 912
rect 1142 858 1146 862
rect 1150 858 1154 862
rect 1166 858 1170 862
rect 1134 808 1138 812
rect 1150 768 1154 772
rect 1182 768 1186 772
rect 1062 758 1066 762
rect 1126 758 1130 762
rect 1062 748 1066 752
rect 1086 748 1090 752
rect 1046 738 1050 742
rect 1050 703 1054 707
rect 1057 703 1061 707
rect 1038 678 1042 682
rect 1030 668 1034 672
rect 1006 628 1010 632
rect 998 618 1002 622
rect 950 588 954 592
rect 926 578 930 582
rect 846 568 850 572
rect 886 568 890 572
rect 902 558 906 562
rect 926 558 930 562
rect 942 558 946 562
rect 1006 608 1010 612
rect 862 548 866 552
rect 878 548 882 552
rect 886 548 890 552
rect 918 548 922 552
rect 990 548 994 552
rect 846 538 850 542
rect 886 528 890 532
rect 838 518 842 522
rect 886 508 890 512
rect 926 538 930 542
rect 950 498 954 502
rect 1094 738 1098 742
rect 1070 618 1074 622
rect 1126 738 1130 742
rect 1126 728 1130 732
rect 1150 728 1154 732
rect 1110 668 1114 672
rect 1110 658 1114 662
rect 1166 708 1170 712
rect 1142 668 1146 672
rect 1142 658 1146 662
rect 1134 648 1138 652
rect 1078 568 1082 572
rect 1014 558 1018 562
rect 1014 528 1018 532
rect 1030 548 1034 552
rect 1062 548 1066 552
rect 1142 548 1146 552
rect 1038 538 1042 542
rect 1030 528 1034 532
rect 902 488 906 492
rect 790 478 794 482
rect 830 478 834 482
rect 766 468 770 472
rect 694 448 698 452
rect 662 338 666 342
rect 606 288 610 292
rect 638 278 642 282
rect 614 268 618 272
rect 606 248 610 252
rect 638 248 642 252
rect 774 458 778 462
rect 766 438 770 442
rect 758 408 762 412
rect 734 338 738 342
rect 670 268 674 272
rect 686 268 690 272
rect 726 308 730 312
rect 718 288 722 292
rect 734 278 738 282
rect 806 468 810 472
rect 838 468 842 472
rect 934 468 938 472
rect 942 468 946 472
rect 806 458 810 462
rect 782 438 786 442
rect 806 438 810 442
rect 790 418 794 422
rect 822 448 826 452
rect 822 418 826 422
rect 814 388 818 392
rect 806 368 810 372
rect 838 438 842 442
rect 870 458 874 462
rect 902 448 906 452
rect 854 418 858 422
rect 870 418 874 422
rect 846 408 850 412
rect 854 408 858 412
rect 782 348 786 352
rect 822 338 826 342
rect 870 338 874 342
rect 798 328 802 332
rect 798 268 802 272
rect 710 258 714 262
rect 782 258 786 262
rect 598 238 602 242
rect 614 238 618 242
rect 630 238 634 242
rect 638 168 642 172
rect 582 158 586 162
rect 630 158 634 162
rect 646 158 650 162
rect 598 148 602 152
rect 550 128 554 132
rect 574 118 578 122
rect 542 108 546 112
rect 534 98 538 102
rect 566 78 570 82
rect 502 68 506 72
rect 670 198 674 202
rect 718 248 722 252
rect 694 218 698 222
rect 686 178 690 182
rect 702 158 706 162
rect 710 148 714 152
rect 686 118 690 122
rect 654 98 658 102
rect 566 58 570 62
rect 758 218 762 222
rect 758 208 762 212
rect 734 168 738 172
rect 798 248 802 252
rect 814 248 818 252
rect 798 238 802 242
rect 790 198 794 202
rect 774 158 778 162
rect 750 148 754 152
rect 774 148 778 152
rect 742 138 746 142
rect 750 98 754 102
rect 758 68 762 72
rect 766 68 770 72
rect 710 59 714 63
rect 830 218 834 222
rect 934 448 938 452
rect 926 428 930 432
rect 966 458 970 462
rect 998 458 1002 462
rect 950 438 954 442
rect 910 368 914 372
rect 910 338 914 342
rect 886 288 890 292
rect 950 328 954 332
rect 918 278 922 282
rect 918 268 922 272
rect 894 248 898 252
rect 910 248 914 252
rect 878 208 882 212
rect 846 188 850 192
rect 838 158 842 162
rect 854 158 858 162
rect 974 308 978 312
rect 1014 438 1018 442
rect 1014 428 1018 432
rect 1158 538 1162 542
rect 1070 518 1074 522
rect 1102 518 1106 522
rect 1050 503 1054 507
rect 1057 503 1061 507
rect 1086 478 1090 482
rect 1046 468 1050 472
rect 1078 468 1082 472
rect 1078 448 1082 452
rect 1030 408 1034 412
rect 1062 418 1066 422
rect 1214 908 1218 912
rect 1206 898 1210 902
rect 1238 958 1242 962
rect 1254 958 1258 962
rect 1254 948 1258 952
rect 1286 1048 1290 1052
rect 1294 1038 1298 1042
rect 1302 947 1306 951
rect 1246 928 1250 932
rect 1230 888 1234 892
rect 1262 888 1266 892
rect 1254 868 1258 872
rect 1302 868 1306 872
rect 1198 858 1202 862
rect 1246 858 1250 862
rect 1350 1048 1354 1052
rect 1326 1008 1330 1012
rect 1390 1118 1394 1122
rect 1414 1118 1418 1122
rect 1374 1098 1378 1102
rect 1406 1098 1410 1102
rect 1454 1148 1458 1152
rect 1446 1128 1450 1132
rect 1486 1158 1490 1162
rect 1502 1148 1506 1152
rect 1478 1138 1482 1142
rect 1502 1138 1506 1142
rect 1462 1128 1466 1132
rect 1518 1128 1522 1132
rect 1478 1088 1482 1092
rect 1454 1068 1458 1072
rect 1422 1048 1426 1052
rect 1438 1048 1442 1052
rect 1406 1018 1410 1022
rect 1398 978 1402 982
rect 1486 1038 1490 1042
rect 1502 1038 1506 1042
rect 1398 968 1402 972
rect 1462 968 1466 972
rect 1366 958 1370 962
rect 1446 958 1450 962
rect 1470 958 1474 962
rect 1438 948 1442 952
rect 1358 928 1362 932
rect 1382 918 1386 922
rect 1358 908 1362 912
rect 1318 898 1322 902
rect 1350 878 1354 882
rect 1374 898 1378 902
rect 1382 888 1386 892
rect 1334 858 1338 862
rect 1310 848 1314 852
rect 1334 808 1338 812
rect 1238 778 1242 782
rect 1294 778 1298 782
rect 1254 768 1258 772
rect 1246 758 1250 762
rect 1270 758 1274 762
rect 1286 758 1290 762
rect 1302 758 1306 762
rect 1238 748 1242 752
rect 1262 738 1266 742
rect 1270 678 1274 682
rect 1230 658 1234 662
rect 1246 658 1250 662
rect 1326 738 1330 742
rect 1302 728 1306 732
rect 1222 648 1226 652
rect 1278 648 1282 652
rect 1294 648 1298 652
rect 1182 548 1186 552
rect 1182 528 1186 532
rect 1190 528 1194 532
rect 1206 478 1210 482
rect 1166 458 1170 462
rect 1118 448 1122 452
rect 1102 428 1106 432
rect 1102 398 1106 402
rect 1070 368 1074 372
rect 1094 368 1098 372
rect 1054 328 1058 332
rect 1070 328 1074 332
rect 1006 308 1010 312
rect 966 288 970 292
rect 982 288 986 292
rect 982 278 986 282
rect 998 258 1002 262
rect 1030 248 1034 252
rect 926 198 930 202
rect 942 168 946 172
rect 790 148 794 152
rect 822 148 826 152
rect 846 148 850 152
rect 998 148 1002 152
rect 814 138 818 142
rect 894 138 898 142
rect 798 128 802 132
rect 790 118 794 122
rect 830 118 834 122
rect 798 108 802 112
rect 806 88 810 92
rect 806 68 810 72
rect 918 98 922 102
rect 910 88 914 92
rect 910 78 914 82
rect 966 88 970 92
rect 934 68 938 72
rect 790 58 794 62
rect 854 58 858 62
rect 926 58 930 62
rect 958 58 962 62
rect 982 78 986 82
rect 1006 78 1010 82
rect 1050 303 1054 307
rect 1057 303 1061 307
rect 1062 288 1066 292
rect 1126 388 1130 392
rect 1182 388 1186 392
rect 1118 368 1122 372
rect 1270 618 1274 622
rect 1230 608 1234 612
rect 1278 578 1282 582
rect 1262 568 1266 572
rect 1246 558 1250 562
rect 1238 508 1242 512
rect 1398 918 1402 922
rect 1430 908 1434 912
rect 1462 898 1466 902
rect 1422 888 1426 892
rect 1430 878 1434 882
rect 1454 878 1458 882
rect 1430 858 1434 862
rect 1390 848 1394 852
rect 1406 848 1410 852
rect 1430 818 1434 822
rect 1390 808 1394 812
rect 1342 768 1346 772
rect 1358 768 1362 772
rect 1406 768 1410 772
rect 1318 638 1322 642
rect 1326 628 1330 632
rect 1422 758 1426 762
rect 1462 768 1466 772
rect 1478 928 1482 932
rect 1646 1328 1650 1332
rect 1598 1258 1602 1262
rect 1630 1258 1634 1262
rect 1686 1278 1690 1282
rect 1662 1268 1666 1272
rect 1638 1208 1642 1212
rect 1562 1203 1566 1207
rect 1569 1203 1573 1207
rect 1598 1188 1602 1192
rect 1582 1168 1586 1172
rect 1534 1158 1538 1162
rect 1566 1158 1570 1162
rect 1566 1148 1570 1152
rect 1558 1138 1562 1142
rect 1566 1088 1570 1092
rect 1534 1068 1538 1072
rect 1646 1158 1650 1162
rect 1678 1248 1682 1252
rect 1798 1338 1802 1342
rect 1806 1338 1810 1342
rect 1734 1328 1738 1332
rect 1702 1318 1706 1322
rect 1710 1288 1714 1292
rect 1726 1288 1730 1292
rect 1726 1278 1730 1282
rect 1750 1278 1754 1282
rect 1702 1258 1706 1262
rect 1782 1258 1786 1262
rect 1766 1238 1770 1242
rect 1758 1218 1762 1222
rect 1750 1168 1754 1172
rect 1702 1148 1706 1152
rect 1726 1138 1730 1142
rect 1686 1128 1690 1132
rect 1790 1148 1794 1152
rect 1782 1138 1786 1142
rect 1662 1098 1666 1102
rect 1670 1098 1674 1102
rect 1718 1098 1722 1102
rect 1734 1098 1738 1102
rect 1654 1088 1658 1092
rect 1638 1078 1642 1082
rect 1646 1078 1650 1082
rect 1614 1068 1618 1072
rect 1622 1068 1626 1072
rect 1686 1068 1690 1072
rect 1598 1038 1602 1042
rect 1614 1038 1618 1042
rect 1606 1028 1610 1032
rect 1630 1028 1634 1032
rect 1562 1003 1566 1007
rect 1569 1003 1573 1007
rect 1630 988 1634 992
rect 1566 968 1570 972
rect 1614 968 1618 972
rect 1526 958 1530 962
rect 1598 958 1602 962
rect 1494 948 1498 952
rect 1582 948 1586 952
rect 1518 938 1522 942
rect 1526 928 1530 932
rect 1502 888 1506 892
rect 1478 868 1482 872
rect 1502 868 1506 872
rect 1358 748 1362 752
rect 1374 748 1378 752
rect 1406 738 1410 742
rect 1350 728 1354 732
rect 1390 728 1394 732
rect 1350 678 1354 682
rect 1390 718 1394 722
rect 1446 748 1450 752
rect 1454 738 1458 742
rect 1446 728 1450 732
rect 1406 708 1410 712
rect 1438 708 1442 712
rect 1430 698 1434 702
rect 1414 678 1418 682
rect 1454 698 1458 702
rect 1462 678 1466 682
rect 1422 658 1426 662
rect 1334 598 1338 602
rect 1318 558 1322 562
rect 1382 648 1386 652
rect 1374 638 1378 642
rect 1350 568 1354 572
rect 1286 538 1290 542
rect 1334 538 1338 542
rect 1518 828 1522 832
rect 1606 938 1610 942
rect 1534 918 1538 922
rect 1598 908 1602 912
rect 1534 898 1538 902
rect 1550 898 1554 902
rect 1542 888 1546 892
rect 1566 888 1570 892
rect 1574 858 1578 862
rect 1662 1058 1666 1062
rect 1710 1038 1714 1042
rect 1654 998 1658 1002
rect 1638 938 1642 942
rect 1734 1088 1738 1092
rect 1766 1078 1770 1082
rect 1678 958 1682 962
rect 1702 948 1706 952
rect 1758 1018 1762 1022
rect 1774 1008 1778 1012
rect 1774 958 1778 962
rect 1734 938 1738 942
rect 1726 908 1730 912
rect 1678 898 1682 902
rect 1606 888 1610 892
rect 1614 878 1618 882
rect 1622 868 1626 872
rect 1638 868 1642 872
rect 1710 868 1714 872
rect 1542 848 1546 852
rect 1534 748 1538 752
rect 1502 738 1506 742
rect 1494 668 1498 672
rect 1502 658 1506 662
rect 1478 638 1482 642
rect 1446 628 1450 632
rect 1494 628 1498 632
rect 1478 618 1482 622
rect 1470 568 1474 572
rect 1406 548 1410 552
rect 1398 528 1402 532
rect 1414 528 1418 532
rect 1398 518 1402 522
rect 1350 488 1354 492
rect 1278 478 1282 482
rect 1366 478 1370 482
rect 1350 468 1354 472
rect 1222 398 1226 402
rect 1166 368 1170 372
rect 1110 338 1114 342
rect 1174 338 1178 342
rect 1110 328 1114 332
rect 1102 288 1106 292
rect 1086 268 1090 272
rect 1150 268 1154 272
rect 1214 368 1218 372
rect 1230 368 1234 372
rect 1342 438 1346 442
rect 1342 428 1346 432
rect 1270 418 1274 422
rect 1246 368 1250 372
rect 1286 368 1290 372
rect 1326 368 1330 372
rect 1206 328 1210 332
rect 1222 318 1226 322
rect 1206 298 1210 302
rect 1070 258 1074 262
rect 1062 238 1066 242
rect 1046 198 1050 202
rect 1078 198 1082 202
rect 1070 188 1074 192
rect 1062 158 1066 162
rect 1102 248 1106 252
rect 1110 218 1114 222
rect 1086 148 1090 152
rect 1062 128 1066 132
rect 1070 108 1074 112
rect 1050 103 1054 107
rect 1057 103 1061 107
rect 1238 268 1242 272
rect 1222 258 1226 262
rect 1238 258 1242 262
rect 1214 228 1218 232
rect 1206 198 1210 202
rect 1198 178 1202 182
rect 1302 328 1306 332
rect 1262 308 1266 312
rect 1270 278 1274 282
rect 1326 278 1330 282
rect 1278 268 1282 272
rect 1302 268 1306 272
rect 1358 268 1362 272
rect 1270 258 1274 262
rect 1334 258 1338 262
rect 1358 258 1362 262
rect 1286 248 1290 252
rect 1302 248 1306 252
rect 1294 238 1298 242
rect 1254 228 1258 232
rect 1254 208 1258 212
rect 1222 178 1226 182
rect 1246 178 1250 182
rect 1214 168 1218 172
rect 1142 148 1146 152
rect 1198 118 1202 122
rect 1150 98 1154 102
rect 1326 218 1330 222
rect 1310 198 1314 202
rect 1254 158 1258 162
rect 1270 158 1274 162
rect 1230 148 1234 152
rect 1262 148 1266 152
rect 1334 178 1338 182
rect 1358 168 1362 172
rect 1310 148 1314 152
rect 1350 148 1354 152
rect 1334 138 1338 142
rect 1318 118 1322 122
rect 1294 108 1298 112
rect 1302 108 1306 112
rect 1246 88 1250 92
rect 1358 128 1362 132
rect 1358 108 1362 112
rect 1342 98 1346 102
rect 1270 78 1274 82
rect 1326 78 1330 82
rect 1382 468 1386 472
rect 1550 838 1554 842
rect 1598 838 1602 842
rect 1550 818 1554 822
rect 1562 803 1566 807
rect 1569 803 1573 807
rect 1558 788 1562 792
rect 1574 778 1578 782
rect 1542 718 1546 722
rect 1542 658 1546 662
rect 1510 608 1514 612
rect 1526 598 1530 602
rect 1502 588 1506 592
rect 1486 548 1490 552
rect 1478 518 1482 522
rect 1510 518 1514 522
rect 1462 478 1466 482
rect 1494 478 1498 482
rect 1542 548 1546 552
rect 1534 508 1538 512
rect 1414 468 1418 472
rect 1502 468 1506 472
rect 1518 468 1522 472
rect 1430 388 1434 392
rect 1438 388 1442 392
rect 1398 378 1402 382
rect 1390 368 1394 372
rect 1414 368 1418 372
rect 1470 438 1474 442
rect 1486 438 1490 442
rect 1446 378 1450 382
rect 1462 368 1466 372
rect 1430 348 1434 352
rect 1462 348 1466 352
rect 1422 338 1426 342
rect 1414 328 1418 332
rect 1398 268 1402 272
rect 1374 248 1378 252
rect 1382 218 1386 222
rect 1462 328 1466 332
rect 1518 448 1522 452
rect 1502 438 1506 442
rect 1502 398 1506 402
rect 1510 378 1514 382
rect 1494 338 1498 342
rect 1502 328 1506 332
rect 1478 318 1482 322
rect 1430 308 1434 312
rect 1542 408 1546 412
rect 1526 388 1530 392
rect 1566 688 1570 692
rect 1590 738 1594 742
rect 1590 698 1594 702
rect 1614 848 1618 852
rect 1718 858 1722 862
rect 1646 848 1650 852
rect 1694 848 1698 852
rect 1638 838 1642 842
rect 1662 828 1666 832
rect 1654 778 1658 782
rect 1654 768 1658 772
rect 1710 798 1714 802
rect 1702 778 1706 782
rect 1718 768 1722 772
rect 1686 758 1690 762
rect 1694 758 1698 762
rect 1774 918 1778 922
rect 1766 898 1770 902
rect 1742 868 1746 872
rect 1750 868 1754 872
rect 1830 1328 1834 1332
rect 1814 1258 1818 1262
rect 1926 1588 1930 1592
rect 1918 1578 1922 1582
rect 1950 1558 1954 1562
rect 1878 1538 1882 1542
rect 1902 1538 1906 1542
rect 1918 1538 1922 1542
rect 1918 1528 1922 1532
rect 1942 1548 1946 1552
rect 1942 1528 1946 1532
rect 2030 1928 2034 1932
rect 2074 1903 2078 1907
rect 2081 1903 2085 1907
rect 2054 1898 2058 1902
rect 2094 1898 2098 1902
rect 2110 1898 2114 1902
rect 2038 1878 2042 1882
rect 2022 1858 2026 1862
rect 2062 1858 2066 1862
rect 1982 1768 1986 1772
rect 1974 1698 1978 1702
rect 2046 1768 2050 1772
rect 2022 1738 2026 1742
rect 2030 1738 2034 1742
rect 2022 1688 2026 1692
rect 1998 1678 2002 1682
rect 1982 1658 1986 1662
rect 1966 1558 1970 1562
rect 1974 1548 1978 1552
rect 1974 1518 1978 1522
rect 1990 1518 1994 1522
rect 1958 1508 1962 1512
rect 1990 1508 1994 1512
rect 1870 1448 1874 1452
rect 1862 1438 1866 1442
rect 1854 1408 1858 1412
rect 1846 1318 1850 1322
rect 1902 1348 1906 1352
rect 1894 1328 1898 1332
rect 1854 1288 1858 1292
rect 1854 1268 1858 1272
rect 1838 1198 1842 1202
rect 1894 1198 1898 1202
rect 1838 1178 1842 1182
rect 1814 1168 1818 1172
rect 1830 1168 1834 1172
rect 1878 1168 1882 1172
rect 1806 1158 1810 1162
rect 1854 1148 1858 1152
rect 1798 1118 1802 1122
rect 1838 1118 1842 1122
rect 1830 1088 1834 1092
rect 1838 1078 1842 1082
rect 1814 1068 1818 1072
rect 1798 1048 1802 1052
rect 1822 1048 1826 1052
rect 1814 1038 1818 1042
rect 1806 968 1810 972
rect 1838 968 1842 972
rect 1830 958 1834 962
rect 1830 948 1834 952
rect 1790 928 1794 932
rect 1806 928 1810 932
rect 1830 928 1834 932
rect 1798 908 1802 912
rect 1790 898 1794 902
rect 1806 868 1810 872
rect 1814 868 1818 872
rect 1750 838 1754 842
rect 1814 828 1818 832
rect 1734 788 1738 792
rect 1814 788 1818 792
rect 1758 758 1762 762
rect 1678 748 1682 752
rect 1702 748 1706 752
rect 1726 748 1730 752
rect 1622 738 1626 742
rect 1606 678 1610 682
rect 1590 668 1594 672
rect 1590 638 1594 642
rect 1606 648 1610 652
rect 1606 628 1610 632
rect 1562 603 1566 607
rect 1569 603 1573 607
rect 1566 528 1570 532
rect 1598 538 1602 542
rect 1646 728 1650 732
rect 1654 728 1658 732
rect 1670 728 1674 732
rect 1638 708 1642 712
rect 1630 698 1634 702
rect 1798 738 1802 742
rect 1822 738 1826 742
rect 1662 668 1666 672
rect 1670 668 1674 672
rect 1694 668 1698 672
rect 1622 658 1626 662
rect 1630 638 1634 642
rect 1646 638 1650 642
rect 1614 488 1618 492
rect 1678 658 1682 662
rect 1702 598 1706 602
rect 1654 588 1658 592
rect 1702 588 1706 592
rect 1678 558 1682 562
rect 1694 558 1698 562
rect 1678 548 1682 552
rect 1670 538 1674 542
rect 1646 528 1650 532
rect 1558 468 1562 472
rect 1606 468 1610 472
rect 1622 438 1626 442
rect 1562 403 1566 407
rect 1569 403 1573 407
rect 1550 378 1554 382
rect 1526 368 1530 372
rect 1542 358 1546 362
rect 1542 338 1546 342
rect 1526 318 1530 322
rect 1542 318 1546 322
rect 1534 308 1538 312
rect 1542 298 1546 302
rect 1502 278 1506 282
rect 1526 278 1530 282
rect 1534 278 1538 282
rect 1446 268 1450 272
rect 1486 268 1490 272
rect 1430 188 1434 192
rect 1478 258 1482 262
rect 1502 258 1506 262
rect 1454 158 1458 162
rect 1462 158 1466 162
rect 1478 158 1482 162
rect 1406 148 1410 152
rect 1462 148 1466 152
rect 1502 147 1506 151
rect 1374 138 1378 142
rect 1414 138 1418 142
rect 1446 138 1450 142
rect 1326 68 1330 72
rect 1342 68 1346 72
rect 1030 58 1034 62
rect 1070 58 1074 62
rect 1126 58 1130 62
rect 1222 58 1226 62
rect 1302 58 1306 62
rect 1510 128 1514 132
rect 1406 118 1410 122
rect 1470 98 1474 102
rect 1494 78 1498 82
rect 1422 58 1426 62
rect 1446 58 1450 62
rect 1702 538 1706 542
rect 1766 688 1770 692
rect 1726 658 1730 662
rect 1742 658 1746 662
rect 1750 658 1754 662
rect 1718 648 1722 652
rect 1734 648 1738 652
rect 1766 648 1770 652
rect 1766 638 1770 642
rect 1766 558 1770 562
rect 1726 548 1730 552
rect 1718 538 1722 542
rect 1710 518 1714 522
rect 1686 498 1690 502
rect 1678 478 1682 482
rect 1742 528 1746 532
rect 1758 528 1762 532
rect 1758 498 1762 502
rect 1742 488 1746 492
rect 1766 478 1770 482
rect 1774 478 1778 482
rect 1718 458 1722 462
rect 1710 448 1714 452
rect 1734 448 1738 452
rect 1726 438 1730 442
rect 1694 418 1698 422
rect 1782 418 1786 422
rect 1718 408 1722 412
rect 1822 648 1826 652
rect 1814 568 1818 572
rect 1806 548 1810 552
rect 1934 1468 1938 1472
rect 1966 1458 1970 1462
rect 1982 1368 1986 1372
rect 1974 1358 1978 1362
rect 1990 1358 1994 1362
rect 1942 1328 1946 1332
rect 1950 1298 1954 1302
rect 1910 1288 1914 1292
rect 1926 1278 1930 1282
rect 1926 1268 1930 1272
rect 1926 1208 1930 1212
rect 1902 1188 1906 1192
rect 1926 1168 1930 1172
rect 1934 1148 1938 1152
rect 1870 1128 1874 1132
rect 1870 1088 1874 1092
rect 1894 1088 1898 1092
rect 1910 1108 1914 1112
rect 1902 1078 1906 1082
rect 2038 1678 2042 1682
rect 2030 1658 2034 1662
rect 2022 1648 2026 1652
rect 2046 1648 2050 1652
rect 2006 1528 2010 1532
rect 2054 1558 2058 1562
rect 2046 1548 2050 1552
rect 2030 1528 2034 1532
rect 2038 1488 2042 1492
rect 2014 1448 2018 1452
rect 2006 1358 2010 1362
rect 2014 1358 2018 1362
rect 2078 1728 2082 1732
rect 2074 1703 2078 1707
rect 2081 1703 2085 1707
rect 2086 1658 2090 1662
rect 2102 1858 2106 1862
rect 2118 1848 2122 1852
rect 2142 1878 2146 1882
rect 2142 1848 2146 1852
rect 2126 1838 2130 1842
rect 2102 1738 2106 1742
rect 2134 1738 2138 1742
rect 2110 1728 2114 1732
rect 2094 1638 2098 1642
rect 2134 1678 2138 1682
rect 2126 1668 2130 1672
rect 2158 2078 2162 2082
rect 2278 2148 2282 2152
rect 2286 2148 2290 2152
rect 2246 2098 2250 2102
rect 2262 2098 2266 2102
rect 2222 2068 2226 2072
rect 2230 2068 2234 2072
rect 2278 2068 2282 2072
rect 2174 2038 2178 2042
rect 2158 2018 2162 2022
rect 2158 1998 2162 2002
rect 2182 2018 2186 2022
rect 2214 1978 2218 1982
rect 2206 1958 2210 1962
rect 2198 1938 2202 1942
rect 2158 1928 2162 1932
rect 2190 1898 2194 1902
rect 2166 1848 2170 1852
rect 2214 1858 2218 1862
rect 2182 1808 2186 1812
rect 2206 1778 2210 1782
rect 2166 1738 2170 1742
rect 2246 2038 2250 2042
rect 2302 2138 2306 2142
rect 2294 2118 2298 2122
rect 2318 2098 2322 2102
rect 2318 2088 2322 2092
rect 2382 2298 2386 2302
rect 2446 2398 2450 2402
rect 2438 2338 2442 2342
rect 2382 2288 2386 2292
rect 2374 2268 2378 2272
rect 2406 2268 2410 2272
rect 2374 2158 2378 2162
rect 2342 2078 2346 2082
rect 2358 2078 2362 2082
rect 2310 2068 2314 2072
rect 2350 2068 2354 2072
rect 2374 2068 2378 2072
rect 2374 2048 2378 2052
rect 2310 2018 2314 2022
rect 2230 1998 2234 2002
rect 2286 1998 2290 2002
rect 2238 1978 2242 1982
rect 2294 1988 2298 1992
rect 2382 2018 2386 2022
rect 2430 2178 2434 2182
rect 2446 2258 2450 2262
rect 2446 2178 2450 2182
rect 2438 2138 2442 2142
rect 2470 2388 2474 2392
rect 2470 2378 2474 2382
rect 2478 2358 2482 2362
rect 2510 2518 2514 2522
rect 2534 2508 2538 2512
rect 2598 2668 2602 2672
rect 2590 2628 2594 2632
rect 2566 2618 2570 2622
rect 2558 2558 2562 2562
rect 2586 2603 2590 2607
rect 2593 2603 2597 2607
rect 2598 2558 2602 2562
rect 2558 2548 2562 2552
rect 2534 2488 2538 2492
rect 2526 2478 2530 2482
rect 2542 2468 2546 2472
rect 2510 2458 2514 2462
rect 2502 2408 2506 2412
rect 2534 2378 2538 2382
rect 2574 2528 2578 2532
rect 2574 2518 2578 2522
rect 2590 2518 2594 2522
rect 2582 2478 2586 2482
rect 2582 2468 2586 2472
rect 2598 2468 2602 2472
rect 2566 2458 2570 2462
rect 2574 2448 2578 2452
rect 2586 2403 2590 2407
rect 2593 2403 2597 2407
rect 2606 2378 2610 2382
rect 2622 2918 2626 2922
rect 2662 2918 2666 2922
rect 2702 2938 2706 2942
rect 2694 2928 2698 2932
rect 2678 2908 2682 2912
rect 2638 2888 2642 2892
rect 2622 2798 2626 2802
rect 2654 2868 2658 2872
rect 2662 2868 2666 2872
rect 2686 2868 2690 2872
rect 2630 2778 2634 2782
rect 2622 2758 2626 2762
rect 2630 2748 2634 2752
rect 2710 2758 2714 2762
rect 2686 2698 2690 2702
rect 2662 2658 2666 2662
rect 2694 2658 2698 2662
rect 2806 3078 2810 3082
rect 2766 3068 2770 3072
rect 2822 3068 2826 3072
rect 2854 3068 2858 3072
rect 2774 3058 2778 3062
rect 2750 2998 2754 3002
rect 2822 3028 2826 3032
rect 2846 3028 2850 3032
rect 2782 2968 2786 2972
rect 2774 2958 2778 2962
rect 2790 2958 2794 2962
rect 2814 2958 2818 2962
rect 2742 2948 2746 2952
rect 2726 2928 2730 2932
rect 2758 2928 2762 2932
rect 2766 2918 2770 2922
rect 2766 2898 2770 2902
rect 2806 2948 2810 2952
rect 2830 2938 2834 2942
rect 2886 3188 2890 3192
rect 3046 3318 3050 3322
rect 3006 3298 3010 3302
rect 3038 3298 3042 3302
rect 3046 3298 3050 3302
rect 3030 3288 3034 3292
rect 2982 3268 2986 3272
rect 2990 3268 2994 3272
rect 2958 3258 2962 3262
rect 2990 3258 2994 3262
rect 2958 3248 2962 3252
rect 2950 3198 2954 3202
rect 3014 3228 3018 3232
rect 2910 3178 2914 3182
rect 2942 3178 2946 3182
rect 2982 3178 2986 3182
rect 2934 3148 2938 3152
rect 2902 3138 2906 3142
rect 2942 3138 2946 3142
rect 2958 3138 2962 3142
rect 2982 3138 2986 3142
rect 2894 3078 2898 3082
rect 2966 3128 2970 3132
rect 2998 3128 3002 3132
rect 3230 3848 3234 3852
rect 3254 3848 3258 3852
rect 3206 3838 3210 3842
rect 3246 3838 3250 3842
rect 3262 3808 3266 3812
rect 3246 3758 3250 3762
rect 3206 3748 3210 3752
rect 3230 3748 3234 3752
rect 3158 3738 3162 3742
rect 3142 3708 3146 3712
rect 3134 3688 3138 3692
rect 3126 3668 3130 3672
rect 3118 3628 3122 3632
rect 3070 3538 3074 3542
rect 3078 3458 3082 3462
rect 3070 3438 3074 3442
rect 3098 3503 3102 3507
rect 3105 3503 3109 3507
rect 3102 3478 3106 3482
rect 3094 3428 3098 3432
rect 3086 3378 3090 3382
rect 3094 3368 3098 3372
rect 3078 3348 3082 3352
rect 3086 3348 3090 3352
rect 3030 3268 3034 3272
rect 3098 3303 3102 3307
rect 3105 3303 3109 3307
rect 3126 3528 3130 3532
rect 3126 3478 3130 3482
rect 3134 3468 3138 3472
rect 3134 3438 3138 3442
rect 3126 3348 3130 3352
rect 3118 3278 3122 3282
rect 3094 3268 3098 3272
rect 3262 3748 3266 3752
rect 3398 3948 3402 3952
rect 3422 3938 3426 3942
rect 3510 3938 3514 3942
rect 3398 3928 3402 3932
rect 3382 3908 3386 3912
rect 3398 3908 3402 3912
rect 3374 3898 3378 3902
rect 3342 3858 3346 3862
rect 3374 3858 3378 3862
rect 3382 3858 3386 3862
rect 3334 3848 3338 3852
rect 3326 3768 3330 3772
rect 3334 3758 3338 3762
rect 3278 3728 3282 3732
rect 3198 3718 3202 3722
rect 3214 3718 3218 3722
rect 3230 3718 3234 3722
rect 3190 3708 3194 3712
rect 3334 3708 3338 3712
rect 3270 3668 3274 3672
rect 3294 3668 3298 3672
rect 3238 3658 3242 3662
rect 3246 3658 3250 3662
rect 3182 3648 3186 3652
rect 3238 3588 3242 3592
rect 3254 3588 3258 3592
rect 3190 3568 3194 3572
rect 3222 3568 3226 3572
rect 3150 3558 3154 3562
rect 3310 3628 3314 3632
rect 3302 3588 3306 3592
rect 3286 3558 3290 3562
rect 3270 3548 3274 3552
rect 3262 3528 3266 3532
rect 3150 3518 3154 3522
rect 3166 3518 3170 3522
rect 3262 3508 3266 3512
rect 3206 3498 3210 3502
rect 3262 3498 3266 3502
rect 3326 3558 3330 3562
rect 3414 3868 3418 3872
rect 3446 3928 3450 3932
rect 3510 3928 3514 3932
rect 3486 3918 3490 3922
rect 3430 3878 3434 3882
rect 3446 3868 3450 3872
rect 3470 3868 3474 3872
rect 3502 3908 3506 3912
rect 3494 3858 3498 3862
rect 3526 3858 3530 3862
rect 3350 3838 3354 3842
rect 3414 3828 3418 3832
rect 3358 3818 3362 3822
rect 3382 3808 3386 3812
rect 3366 3788 3370 3792
rect 3374 3768 3378 3772
rect 3390 3778 3394 3782
rect 3398 3748 3402 3752
rect 3358 3738 3362 3742
rect 3406 3718 3410 3722
rect 3374 3698 3378 3702
rect 3398 3698 3402 3702
rect 3398 3688 3402 3692
rect 3414 3708 3418 3712
rect 3430 3708 3434 3712
rect 3422 3698 3426 3702
rect 3430 3688 3434 3692
rect 3398 3668 3402 3672
rect 3486 3838 3490 3842
rect 3446 3788 3450 3792
rect 3470 3688 3474 3692
rect 3446 3668 3450 3672
rect 3462 3668 3466 3672
rect 3390 3658 3394 3662
rect 3406 3658 3410 3662
rect 3422 3648 3426 3652
rect 3534 3778 3538 3782
rect 3542 3768 3546 3772
rect 3510 3748 3514 3752
rect 3526 3748 3530 3752
rect 3630 4038 3634 4042
rect 3670 4018 3674 4022
rect 3590 4008 3594 4012
rect 3610 4003 3614 4007
rect 3617 4003 3621 4007
rect 3590 3988 3594 3992
rect 3574 3968 3578 3972
rect 3662 3958 3666 3962
rect 3574 3948 3578 3952
rect 3598 3948 3602 3952
rect 3630 3948 3634 3952
rect 3558 3898 3562 3902
rect 3670 3938 3674 3942
rect 3662 3888 3666 3892
rect 3614 3868 3618 3872
rect 3582 3838 3586 3842
rect 3574 3828 3578 3832
rect 3574 3788 3578 3792
rect 3638 3838 3642 3842
rect 3654 3838 3658 3842
rect 3598 3828 3602 3832
rect 3574 3748 3578 3752
rect 3526 3728 3530 3732
rect 3558 3728 3562 3732
rect 3494 3718 3498 3722
rect 3526 3718 3530 3722
rect 3534 3708 3538 3712
rect 3510 3668 3514 3672
rect 3534 3668 3538 3672
rect 3438 3658 3442 3662
rect 3470 3658 3474 3662
rect 3454 3648 3458 3652
rect 3430 3638 3434 3642
rect 3350 3608 3354 3612
rect 3374 3608 3378 3612
rect 3390 3608 3394 3612
rect 3438 3558 3442 3562
rect 3414 3548 3418 3552
rect 3334 3538 3338 3542
rect 3342 3538 3346 3542
rect 3286 3488 3290 3492
rect 3294 3488 3298 3492
rect 3270 3468 3274 3472
rect 3158 3458 3162 3462
rect 3190 3458 3194 3462
rect 3238 3458 3242 3462
rect 3174 3428 3178 3432
rect 3254 3448 3258 3452
rect 3286 3448 3290 3452
rect 3262 3418 3266 3422
rect 3246 3408 3250 3412
rect 3142 3398 3146 3402
rect 3166 3378 3170 3382
rect 3150 3338 3154 3342
rect 3142 3318 3146 3322
rect 3142 3278 3146 3282
rect 3134 3268 3138 3272
rect 3110 3258 3114 3262
rect 3118 3258 3122 3262
rect 3126 3258 3130 3262
rect 3086 3198 3090 3202
rect 3094 3188 3098 3192
rect 3046 3178 3050 3182
rect 3094 3178 3098 3182
rect 3070 3168 3074 3172
rect 3022 3148 3026 3152
rect 3150 3148 3154 3152
rect 3030 3138 3034 3142
rect 3062 3138 3066 3142
rect 2886 3058 2890 3062
rect 2918 3058 2922 3062
rect 2878 3048 2882 3052
rect 2870 3038 2874 3042
rect 2886 3038 2890 3042
rect 2950 3048 2954 3052
rect 2902 3038 2906 3042
rect 2854 2918 2858 2922
rect 2870 2898 2874 2902
rect 2934 3008 2938 3012
rect 2958 2998 2962 3002
rect 2894 2958 2898 2962
rect 2918 2958 2922 2962
rect 2982 2958 2986 2962
rect 3014 3098 3018 3102
rect 3070 3098 3074 3102
rect 3062 3088 3066 3092
rect 3046 3078 3050 3082
rect 3062 3078 3066 3082
rect 3030 3068 3034 3072
rect 3014 3058 3018 3062
rect 3022 3058 3026 3062
rect 3134 3118 3138 3122
rect 3098 3103 3102 3107
rect 3105 3103 3109 3107
rect 3078 3088 3082 3092
rect 3142 3068 3146 3072
rect 3318 3528 3322 3532
rect 3350 3518 3354 3522
rect 3358 3468 3362 3472
rect 3358 3458 3362 3462
rect 3318 3448 3322 3452
rect 3342 3448 3346 3452
rect 3358 3438 3362 3442
rect 3382 3458 3386 3462
rect 3414 3528 3418 3532
rect 3430 3528 3434 3532
rect 3422 3508 3426 3512
rect 3454 3548 3458 3552
rect 3518 3658 3522 3662
rect 3502 3608 3506 3612
rect 3494 3568 3498 3572
rect 3478 3558 3482 3562
rect 3526 3558 3530 3562
rect 3478 3548 3482 3552
rect 3510 3538 3514 3542
rect 3518 3538 3522 3542
rect 3446 3518 3450 3522
rect 3438 3488 3442 3492
rect 3406 3478 3410 3482
rect 3454 3478 3458 3482
rect 3414 3468 3418 3472
rect 3430 3468 3434 3472
rect 3398 3448 3402 3452
rect 3406 3448 3410 3452
rect 3374 3428 3378 3432
rect 3302 3388 3306 3392
rect 3318 3388 3322 3392
rect 3310 3378 3314 3382
rect 3278 3368 3282 3372
rect 3278 3358 3282 3362
rect 3326 3358 3330 3362
rect 3262 3348 3266 3352
rect 3182 3268 3186 3272
rect 3222 3328 3226 3332
rect 3310 3338 3314 3342
rect 3270 3318 3274 3322
rect 3270 3288 3274 3292
rect 3254 3278 3258 3282
rect 3214 3268 3218 3272
rect 3206 3258 3210 3262
rect 3198 3208 3202 3212
rect 3214 3198 3218 3202
rect 3222 3188 3226 3192
rect 3214 3148 3218 3152
rect 3182 3128 3186 3132
rect 3214 3068 3218 3072
rect 3094 3058 3098 3062
rect 3110 3048 3114 3052
rect 3102 3038 3106 3042
rect 3142 3048 3146 3052
rect 3134 2998 3138 3002
rect 3022 2988 3026 2992
rect 2950 2948 2954 2952
rect 2998 2948 3002 2952
rect 2974 2938 2978 2942
rect 2998 2938 3002 2942
rect 2950 2918 2954 2922
rect 2902 2908 2906 2912
rect 2782 2868 2786 2872
rect 2790 2868 2794 2872
rect 2814 2868 2818 2872
rect 2846 2868 2850 2872
rect 2854 2868 2858 2872
rect 2886 2868 2890 2872
rect 2750 2838 2754 2842
rect 2798 2838 2802 2842
rect 2814 2828 2818 2832
rect 2766 2768 2770 2772
rect 2798 2768 2802 2772
rect 2782 2758 2786 2762
rect 2838 2858 2842 2862
rect 2838 2838 2842 2842
rect 2822 2788 2826 2792
rect 2830 2788 2834 2792
rect 2758 2738 2762 2742
rect 2830 2768 2834 2772
rect 2846 2758 2850 2762
rect 2774 2728 2778 2732
rect 2846 2728 2850 2732
rect 2854 2728 2858 2732
rect 2766 2718 2770 2722
rect 2822 2698 2826 2702
rect 2806 2668 2810 2672
rect 2726 2658 2730 2662
rect 2718 2648 2722 2652
rect 2790 2648 2794 2652
rect 2622 2588 2626 2592
rect 2654 2598 2658 2602
rect 2662 2588 2666 2592
rect 2702 2588 2706 2592
rect 2646 2568 2650 2572
rect 2630 2558 2634 2562
rect 2694 2558 2698 2562
rect 2662 2548 2666 2552
rect 2622 2538 2626 2542
rect 2630 2528 2634 2532
rect 2654 2528 2658 2532
rect 2654 2488 2658 2492
rect 2638 2478 2642 2482
rect 2638 2468 2642 2472
rect 2630 2428 2634 2432
rect 2654 2398 2658 2402
rect 2686 2518 2690 2522
rect 2710 2508 2714 2512
rect 2694 2498 2698 2502
rect 2702 2498 2706 2502
rect 2678 2488 2682 2492
rect 2686 2468 2690 2472
rect 2702 2468 2706 2472
rect 2710 2458 2714 2462
rect 2694 2448 2698 2452
rect 2678 2418 2682 2422
rect 2646 2378 2650 2382
rect 2550 2368 2554 2372
rect 2614 2368 2618 2372
rect 2518 2348 2522 2352
rect 2590 2348 2594 2352
rect 2614 2348 2618 2352
rect 2494 2338 2498 2342
rect 2502 2338 2506 2342
rect 2502 2328 2506 2332
rect 2486 2318 2490 2322
rect 2510 2318 2514 2322
rect 2534 2328 2538 2332
rect 2574 2338 2578 2342
rect 2614 2338 2618 2342
rect 2550 2278 2554 2282
rect 2566 2278 2570 2282
rect 2534 2258 2538 2262
rect 2534 2218 2538 2222
rect 2502 2208 2506 2212
rect 2518 2208 2522 2212
rect 2478 2188 2482 2192
rect 2510 2188 2514 2192
rect 2470 2168 2474 2172
rect 2502 2148 2506 2152
rect 2486 2138 2490 2142
rect 2502 2108 2506 2112
rect 2398 2088 2402 2092
rect 2422 2088 2426 2092
rect 2526 2158 2530 2162
rect 2542 2148 2546 2152
rect 2526 2128 2530 2132
rect 2534 2108 2538 2112
rect 2430 2078 2434 2082
rect 2510 2078 2514 2082
rect 2462 2068 2466 2072
rect 2438 2038 2442 2042
rect 2406 2028 2410 2032
rect 2398 2018 2402 2022
rect 2390 1998 2394 2002
rect 2350 1947 2354 1951
rect 2294 1938 2298 1942
rect 2334 1938 2338 1942
rect 2390 1938 2394 1942
rect 2270 1898 2274 1902
rect 2382 1888 2386 1892
rect 2230 1878 2234 1882
rect 2294 1878 2298 1882
rect 2358 1878 2362 1882
rect 2414 1948 2418 1952
rect 2406 1938 2410 1942
rect 2422 1938 2426 1942
rect 2438 1938 2442 1942
rect 2414 1918 2418 1922
rect 2350 1868 2354 1872
rect 2430 1928 2434 1932
rect 2438 1888 2442 1892
rect 2422 1868 2426 1872
rect 2278 1858 2282 1862
rect 2366 1858 2370 1862
rect 2382 1858 2386 1862
rect 2406 1858 2410 1862
rect 2382 1848 2386 1852
rect 2246 1838 2250 1842
rect 2430 1838 2434 1842
rect 2222 1808 2226 1812
rect 2606 2238 2610 2242
rect 2590 2218 2594 2222
rect 2606 2208 2610 2212
rect 2586 2203 2590 2207
rect 2593 2203 2597 2207
rect 2590 2188 2594 2192
rect 2590 2108 2594 2112
rect 2542 2088 2546 2092
rect 2550 2078 2554 2082
rect 2486 2048 2490 2052
rect 2486 2028 2490 2032
rect 2462 1988 2466 1992
rect 2454 1928 2458 1932
rect 2454 1858 2458 1862
rect 2478 1958 2482 1962
rect 2582 2068 2586 2072
rect 2630 2308 2634 2312
rect 2630 2148 2634 2152
rect 2694 2368 2698 2372
rect 2678 2308 2682 2312
rect 2654 2268 2658 2272
rect 2678 2268 2682 2272
rect 2646 2248 2650 2252
rect 2646 2148 2650 2152
rect 2614 2058 2618 2062
rect 2606 2038 2610 2042
rect 2542 2008 2546 2012
rect 2586 2003 2590 2007
rect 2593 2003 2597 2007
rect 2502 1968 2506 1972
rect 2494 1958 2498 1962
rect 2542 1958 2546 1962
rect 2558 1958 2562 1962
rect 2470 1938 2474 1942
rect 2526 1938 2530 1942
rect 2582 1948 2586 1952
rect 2566 1938 2570 1942
rect 2494 1898 2498 1902
rect 2486 1858 2490 1862
rect 2478 1838 2482 1842
rect 2486 1838 2490 1842
rect 2518 1778 2522 1782
rect 2310 1768 2314 1772
rect 2414 1768 2418 1772
rect 2430 1768 2434 1772
rect 2462 1768 2466 1772
rect 2262 1758 2266 1762
rect 2230 1748 2234 1752
rect 2230 1738 2234 1742
rect 2198 1728 2202 1732
rect 2214 1728 2218 1732
rect 2278 1728 2282 1732
rect 2166 1688 2170 1692
rect 2174 1688 2178 1692
rect 2182 1678 2186 1682
rect 2150 1658 2154 1662
rect 2174 1658 2178 1662
rect 2150 1638 2154 1642
rect 2158 1638 2162 1642
rect 2110 1618 2114 1622
rect 2078 1588 2082 1592
rect 2078 1578 2082 1582
rect 2102 1578 2106 1582
rect 2094 1548 2098 1552
rect 2074 1503 2078 1507
rect 2081 1503 2085 1507
rect 2110 1558 2114 1562
rect 2110 1518 2114 1522
rect 2150 1598 2154 1602
rect 2150 1578 2154 1582
rect 2142 1558 2146 1562
rect 2150 1548 2154 1552
rect 2126 1528 2130 1532
rect 2158 1528 2162 1532
rect 2142 1518 2146 1522
rect 2158 1518 2162 1522
rect 2118 1498 2122 1502
rect 2126 1488 2130 1492
rect 2174 1558 2178 1562
rect 2182 1558 2186 1562
rect 2214 1718 2218 1722
rect 2390 1748 2394 1752
rect 2374 1728 2378 1732
rect 2222 1688 2226 1692
rect 2318 1688 2322 1692
rect 2246 1678 2250 1682
rect 2262 1678 2266 1682
rect 2350 1678 2354 1682
rect 2222 1658 2226 1662
rect 2254 1658 2258 1662
rect 2230 1588 2234 1592
rect 2198 1558 2202 1562
rect 2166 1478 2170 1482
rect 2102 1468 2106 1472
rect 2110 1468 2114 1472
rect 2126 1468 2130 1472
rect 2158 1468 2162 1472
rect 2038 1408 2042 1412
rect 2062 1408 2066 1412
rect 2094 1448 2098 1452
rect 2102 1448 2106 1452
rect 2118 1438 2122 1442
rect 2142 1438 2146 1442
rect 2102 1418 2106 1422
rect 2070 1368 2074 1372
rect 2086 1368 2090 1372
rect 2062 1358 2066 1362
rect 2086 1328 2090 1332
rect 2094 1308 2098 1312
rect 2074 1303 2078 1307
rect 2081 1303 2085 1307
rect 2126 1368 2130 1372
rect 2110 1358 2114 1362
rect 2142 1328 2146 1332
rect 2022 1288 2026 1292
rect 2046 1288 2050 1292
rect 2054 1288 2058 1292
rect 2094 1288 2098 1292
rect 1998 1278 2002 1282
rect 1974 1268 1978 1272
rect 2030 1268 2034 1272
rect 1982 1258 1986 1262
rect 1958 1078 1962 1082
rect 1886 1068 1890 1072
rect 1894 1068 1898 1072
rect 1918 1068 1922 1072
rect 1854 1028 1858 1032
rect 1846 908 1850 912
rect 1838 888 1842 892
rect 1838 838 1842 842
rect 1910 1058 1914 1062
rect 1902 1048 1906 1052
rect 1926 1048 1930 1052
rect 1870 898 1874 902
rect 1870 878 1874 882
rect 1942 988 1946 992
rect 1902 968 1906 972
rect 1854 808 1858 812
rect 1862 798 1866 802
rect 1862 568 1866 572
rect 1894 848 1898 852
rect 1894 788 1898 792
rect 1894 698 1898 702
rect 1910 948 1914 952
rect 1982 1138 1986 1142
rect 1974 1108 1978 1112
rect 2046 1238 2050 1242
rect 2006 1218 2010 1222
rect 2030 1188 2034 1192
rect 1998 1138 2002 1142
rect 1990 1128 1994 1132
rect 2006 1088 2010 1092
rect 2022 1078 2026 1082
rect 2038 1138 2042 1142
rect 2062 1248 2066 1252
rect 2054 1208 2058 1212
rect 2054 1158 2058 1162
rect 2022 1058 2026 1062
rect 2030 1038 2034 1042
rect 1982 1028 1986 1032
rect 1974 1008 1978 1012
rect 2022 998 2026 1002
rect 1966 988 1970 992
rect 1982 978 1986 982
rect 2014 968 2018 972
rect 1998 958 2002 962
rect 1918 938 1922 942
rect 1910 908 1914 912
rect 1910 888 1914 892
rect 2094 1258 2098 1262
rect 2094 1248 2098 1252
rect 2078 1238 2082 1242
rect 2110 1228 2114 1232
rect 2126 1298 2130 1302
rect 2158 1338 2162 1342
rect 2150 1298 2154 1302
rect 2222 1548 2226 1552
rect 2230 1548 2234 1552
rect 2270 1628 2274 1632
rect 2286 1588 2290 1592
rect 2294 1578 2298 1582
rect 2262 1538 2266 1542
rect 2206 1528 2210 1532
rect 2278 1548 2282 1552
rect 2286 1538 2290 1542
rect 2254 1528 2258 1532
rect 2270 1528 2274 1532
rect 2190 1518 2194 1522
rect 2214 1518 2218 1522
rect 2214 1508 2218 1512
rect 2206 1498 2210 1502
rect 2198 1468 2202 1472
rect 2246 1478 2250 1482
rect 2190 1448 2194 1452
rect 2182 1438 2186 1442
rect 2206 1438 2210 1442
rect 2190 1418 2194 1422
rect 2174 1358 2178 1362
rect 2158 1258 2162 1262
rect 2142 1238 2146 1242
rect 2126 1208 2130 1212
rect 2118 1198 2122 1202
rect 2118 1168 2122 1172
rect 2110 1158 2114 1162
rect 2070 1138 2074 1142
rect 2074 1103 2078 1107
rect 2081 1103 2085 1107
rect 2046 1088 2050 1092
rect 2078 1068 2082 1072
rect 2182 1298 2186 1302
rect 2238 1448 2242 1452
rect 2246 1448 2250 1452
rect 2230 1438 2234 1442
rect 2198 1368 2202 1372
rect 2214 1368 2218 1372
rect 2222 1368 2226 1372
rect 2222 1348 2226 1352
rect 2198 1318 2202 1322
rect 2214 1318 2218 1322
rect 2214 1308 2218 1312
rect 2286 1478 2290 1482
rect 2262 1448 2266 1452
rect 2302 1548 2306 1552
rect 2438 1758 2442 1762
rect 2462 1758 2466 1762
rect 2566 1848 2570 1852
rect 2550 1778 2554 1782
rect 2558 1758 2562 1762
rect 2590 1878 2594 1882
rect 2586 1803 2590 1807
rect 2593 1803 2597 1807
rect 2406 1748 2410 1752
rect 2478 1748 2482 1752
rect 2486 1748 2490 1752
rect 2502 1748 2506 1752
rect 2542 1748 2546 1752
rect 2566 1748 2570 1752
rect 2422 1728 2426 1732
rect 2430 1728 2434 1732
rect 2414 1718 2418 1722
rect 2510 1728 2514 1732
rect 2438 1688 2442 1692
rect 2478 1688 2482 1692
rect 2406 1678 2410 1682
rect 2502 1678 2506 1682
rect 2390 1668 2394 1672
rect 2454 1668 2458 1672
rect 2430 1658 2434 1662
rect 2350 1648 2354 1652
rect 2318 1638 2322 1642
rect 2318 1608 2322 1612
rect 2342 1598 2346 1602
rect 2334 1538 2338 1542
rect 2342 1538 2346 1542
rect 2318 1498 2322 1502
rect 2342 1478 2346 1482
rect 2334 1448 2338 1452
rect 2294 1438 2298 1442
rect 2254 1418 2258 1422
rect 2286 1408 2290 1412
rect 2302 1358 2306 1362
rect 2318 1358 2322 1362
rect 2334 1358 2338 1362
rect 2366 1638 2370 1642
rect 2422 1638 2426 1642
rect 2430 1638 2434 1642
rect 2398 1608 2402 1612
rect 2422 1608 2426 1612
rect 2390 1588 2394 1592
rect 2414 1588 2418 1592
rect 2358 1548 2362 1552
rect 2374 1538 2378 1542
rect 2358 1518 2362 1522
rect 2350 1418 2354 1422
rect 2358 1408 2362 1412
rect 2246 1348 2250 1352
rect 2326 1348 2330 1352
rect 2270 1338 2274 1342
rect 2326 1338 2330 1342
rect 2350 1338 2354 1342
rect 2326 1328 2330 1332
rect 2246 1318 2250 1322
rect 2230 1288 2234 1292
rect 2286 1288 2290 1292
rect 2278 1268 2282 1272
rect 2310 1268 2314 1272
rect 2246 1258 2250 1262
rect 2270 1258 2274 1262
rect 2206 1238 2210 1242
rect 2198 1218 2202 1222
rect 2190 1188 2194 1192
rect 2182 1178 2186 1182
rect 2174 1158 2178 1162
rect 2102 1138 2106 1142
rect 2190 1138 2194 1142
rect 2118 1098 2122 1102
rect 2102 1078 2106 1082
rect 2094 1058 2098 1062
rect 2118 1058 2122 1062
rect 2086 1048 2090 1052
rect 2110 1038 2114 1042
rect 2150 1048 2154 1052
rect 2150 1028 2154 1032
rect 2118 998 2122 1002
rect 2046 978 2050 982
rect 2110 958 2114 962
rect 1966 908 1970 912
rect 2006 908 2010 912
rect 2022 908 2026 912
rect 1958 888 1962 892
rect 1958 878 1962 882
rect 1966 868 1970 872
rect 2022 898 2026 902
rect 2014 848 2018 852
rect 2094 938 2098 942
rect 2074 903 2078 907
rect 2081 903 2085 907
rect 2078 888 2082 892
rect 2038 878 2042 882
rect 2070 868 2074 872
rect 2054 848 2058 852
rect 2078 808 2082 812
rect 2070 788 2074 792
rect 2126 908 2130 912
rect 2102 888 2106 892
rect 2134 888 2138 892
rect 2174 958 2178 962
rect 2238 1198 2242 1202
rect 2270 1248 2274 1252
rect 2254 1218 2258 1222
rect 2302 1248 2306 1252
rect 2294 1208 2298 1212
rect 2318 1158 2322 1162
rect 2342 1158 2346 1162
rect 2262 1148 2266 1152
rect 2278 1138 2282 1142
rect 2302 1118 2306 1122
rect 2246 1108 2250 1112
rect 2270 1108 2274 1112
rect 2286 1108 2290 1112
rect 2238 1098 2242 1102
rect 2302 1098 2306 1102
rect 2206 1088 2210 1092
rect 2270 1088 2274 1092
rect 2230 1068 2234 1072
rect 2254 1068 2258 1072
rect 2246 1058 2250 1062
rect 2262 1058 2266 1062
rect 2214 1048 2218 1052
rect 2222 1028 2226 1032
rect 2206 998 2210 1002
rect 2190 948 2194 952
rect 2358 1258 2362 1262
rect 2398 1518 2402 1522
rect 2414 1518 2418 1522
rect 2406 1508 2410 1512
rect 2390 1488 2394 1492
rect 2406 1468 2410 1472
rect 2454 1518 2458 1522
rect 2430 1508 2434 1512
rect 2422 1498 2426 1502
rect 2422 1488 2426 1492
rect 2454 1498 2458 1502
rect 2446 1488 2450 1492
rect 2486 1518 2490 1522
rect 2430 1468 2434 1472
rect 2462 1468 2466 1472
rect 2414 1418 2418 1422
rect 2398 1398 2402 1402
rect 2414 1358 2418 1362
rect 2390 1328 2394 1332
rect 2454 1458 2458 1462
rect 2550 1688 2554 1692
rect 2526 1558 2530 1562
rect 2566 1648 2570 1652
rect 2590 1618 2594 1622
rect 2586 1603 2590 1607
rect 2593 1603 2597 1607
rect 2566 1588 2570 1592
rect 2510 1508 2514 1512
rect 2502 1478 2506 1482
rect 2550 1518 2554 1522
rect 2550 1458 2554 1462
rect 2622 1998 2626 2002
rect 2622 1978 2626 1982
rect 2622 1968 2626 1972
rect 2614 1928 2618 1932
rect 2654 2008 2658 2012
rect 2646 1998 2650 2002
rect 2670 2128 2674 2132
rect 2694 2298 2698 2302
rect 2742 2628 2746 2632
rect 2790 2588 2794 2592
rect 2774 2558 2778 2562
rect 2830 2668 2834 2672
rect 2822 2648 2826 2652
rect 2846 2708 2850 2712
rect 2886 2828 2890 2832
rect 2942 2888 2946 2892
rect 2918 2858 2922 2862
rect 2894 2808 2898 2812
rect 2902 2778 2906 2782
rect 2894 2768 2898 2772
rect 2886 2758 2890 2762
rect 2878 2738 2882 2742
rect 2886 2738 2890 2742
rect 2878 2718 2882 2722
rect 2870 2698 2874 2702
rect 2854 2678 2858 2682
rect 2870 2668 2874 2672
rect 2966 2868 2970 2872
rect 2990 2868 2994 2872
rect 3046 2978 3050 2982
rect 3030 2898 3034 2902
rect 3054 2958 3058 2962
rect 3070 2958 3074 2962
rect 3134 2958 3138 2962
rect 3118 2948 3122 2952
rect 3102 2938 3106 2942
rect 3150 2948 3154 2952
rect 3078 2908 3082 2912
rect 3062 2888 3066 2892
rect 3098 2903 3102 2907
rect 3105 2903 3109 2907
rect 3054 2868 3058 2872
rect 3142 2868 3146 2872
rect 2982 2858 2986 2862
rect 3038 2858 3042 2862
rect 2894 2668 2898 2672
rect 2918 2668 2922 2672
rect 2886 2658 2890 2662
rect 2862 2648 2866 2652
rect 2894 2648 2898 2652
rect 2910 2648 2914 2652
rect 2862 2598 2866 2602
rect 2846 2568 2850 2572
rect 2814 2558 2818 2562
rect 2830 2558 2834 2562
rect 2750 2548 2754 2552
rect 2758 2548 2762 2552
rect 2774 2548 2778 2552
rect 2822 2548 2826 2552
rect 2854 2548 2858 2552
rect 2750 2528 2754 2532
rect 2758 2528 2762 2532
rect 2726 2518 2730 2522
rect 2742 2498 2746 2502
rect 2734 2478 2738 2482
rect 2742 2458 2746 2462
rect 2782 2508 2786 2512
rect 2798 2478 2802 2482
rect 2774 2448 2778 2452
rect 2782 2448 2786 2452
rect 2758 2438 2762 2442
rect 2734 2378 2738 2382
rect 2718 2288 2722 2292
rect 2702 2278 2706 2282
rect 2702 2258 2706 2262
rect 2838 2518 2842 2522
rect 2846 2518 2850 2522
rect 2814 2468 2818 2472
rect 2870 2588 2874 2592
rect 2886 2568 2890 2572
rect 2894 2548 2898 2552
rect 2910 2528 2914 2532
rect 2926 2658 2930 2662
rect 2966 2728 2970 2732
rect 3014 2848 3018 2852
rect 3030 2788 3034 2792
rect 3022 2738 3026 2742
rect 2998 2728 3002 2732
rect 2974 2688 2978 2692
rect 2998 2658 3002 2662
rect 3046 2768 3050 2772
rect 3110 2858 3114 2862
rect 3078 2848 3082 2852
rect 3094 2848 3098 2852
rect 3086 2768 3090 2772
rect 3054 2738 3058 2742
rect 3086 2738 3090 2742
rect 3142 2778 3146 2782
rect 3062 2698 3066 2702
rect 3070 2678 3074 2682
rect 3126 2728 3130 2732
rect 3118 2708 3122 2712
rect 3098 2703 3102 2707
rect 3105 2703 3109 2707
rect 3126 2678 3130 2682
rect 3110 2668 3114 2672
rect 3086 2658 3090 2662
rect 2966 2608 2970 2612
rect 2982 2608 2986 2612
rect 2958 2588 2962 2592
rect 2934 2558 2938 2562
rect 2950 2548 2954 2552
rect 2966 2548 2970 2552
rect 2974 2548 2978 2552
rect 3214 2978 3218 2982
rect 3198 2948 3202 2952
rect 3182 2938 3186 2942
rect 3174 2918 3178 2922
rect 3166 2898 3170 2902
rect 3166 2888 3170 2892
rect 3190 2888 3194 2892
rect 3206 2888 3210 2892
rect 3206 2858 3210 2862
rect 3246 3178 3250 3182
rect 3398 3408 3402 3412
rect 3382 3378 3386 3382
rect 3438 3438 3442 3442
rect 3454 3438 3458 3442
rect 3462 3438 3466 3442
rect 3422 3428 3426 3432
rect 3374 3368 3378 3372
rect 3414 3368 3418 3372
rect 3358 3338 3362 3342
rect 3406 3308 3410 3312
rect 3318 3298 3322 3302
rect 3334 3298 3338 3302
rect 3374 3288 3378 3292
rect 3350 3278 3354 3282
rect 3262 3268 3266 3272
rect 3310 3258 3314 3262
rect 3326 3258 3330 3262
rect 3270 3248 3274 3252
rect 3278 3178 3282 3182
rect 3230 3148 3234 3152
rect 3246 3148 3250 3152
rect 3238 3128 3242 3132
rect 3238 2978 3242 2982
rect 3246 2968 3250 2972
rect 3286 3138 3290 3142
rect 3294 3128 3298 3132
rect 3334 3228 3338 3232
rect 3310 3118 3314 3122
rect 3342 3198 3346 3202
rect 3318 3068 3322 3072
rect 3334 3068 3338 3072
rect 3406 3288 3410 3292
rect 3422 3278 3426 3282
rect 3454 3338 3458 3342
rect 3374 3258 3378 3262
rect 3398 3258 3402 3262
rect 3438 3258 3442 3262
rect 3454 3258 3458 3262
rect 3374 3228 3378 3232
rect 3398 3218 3402 3222
rect 3390 3198 3394 3202
rect 3390 3178 3394 3182
rect 3350 3148 3354 3152
rect 3366 3148 3370 3152
rect 3414 3148 3418 3152
rect 3358 3138 3362 3142
rect 3398 3138 3402 3142
rect 3358 3088 3362 3092
rect 3350 3078 3354 3082
rect 3310 3058 3314 3062
rect 3342 3058 3346 3062
rect 3270 2998 3274 3002
rect 3238 2918 3242 2922
rect 3238 2888 3242 2892
rect 3206 2848 3210 2852
rect 3174 2788 3178 2792
rect 3166 2778 3170 2782
rect 3262 2938 3266 2942
rect 3286 2958 3290 2962
rect 3342 2968 3346 2972
rect 3326 2938 3330 2942
rect 3318 2878 3322 2882
rect 3246 2828 3250 2832
rect 3254 2828 3258 2832
rect 3222 2768 3226 2772
rect 3262 2768 3266 2772
rect 3246 2748 3250 2752
rect 3198 2708 3202 2712
rect 3182 2698 3186 2702
rect 3166 2648 3170 2652
rect 3158 2638 3162 2642
rect 3142 2628 3146 2632
rect 3110 2618 3114 2622
rect 3174 2608 3178 2612
rect 3198 2608 3202 2612
rect 3078 2598 3082 2602
rect 3030 2588 3034 2592
rect 3014 2578 3018 2582
rect 3006 2538 3010 2542
rect 2966 2528 2970 2532
rect 2918 2518 2922 2522
rect 2918 2508 2922 2512
rect 2902 2498 2906 2502
rect 2806 2418 2810 2422
rect 2782 2408 2786 2412
rect 2798 2408 2802 2412
rect 2950 2498 2954 2502
rect 2966 2488 2970 2492
rect 2934 2458 2938 2462
rect 2950 2458 2954 2462
rect 2830 2448 2834 2452
rect 2902 2428 2906 2432
rect 2838 2408 2842 2412
rect 2822 2378 2826 2382
rect 2814 2358 2818 2362
rect 2742 2348 2746 2352
rect 2726 2268 2730 2272
rect 2734 2168 2738 2172
rect 2734 2108 2738 2112
rect 2710 2078 2714 2082
rect 2734 2078 2738 2082
rect 2710 2068 2714 2072
rect 2734 2058 2738 2062
rect 2702 2048 2706 2052
rect 2726 2038 2730 2042
rect 2662 1988 2666 1992
rect 2646 1978 2650 1982
rect 2638 1968 2642 1972
rect 2718 1968 2722 1972
rect 2670 1958 2674 1962
rect 2702 1938 2706 1942
rect 2726 1928 2730 1932
rect 2710 1918 2714 1922
rect 2646 1908 2650 1912
rect 2638 1898 2642 1902
rect 2702 1878 2706 1882
rect 2630 1868 2634 1872
rect 2678 1868 2682 1872
rect 2614 1858 2618 1862
rect 2614 1828 2618 1832
rect 2718 1828 2722 1832
rect 2622 1768 2626 1772
rect 2774 2338 2778 2342
rect 2790 2328 2794 2332
rect 2758 2308 2762 2312
rect 2750 2298 2754 2302
rect 2750 2248 2754 2252
rect 2822 2348 2826 2352
rect 2886 2348 2890 2352
rect 2822 2298 2826 2302
rect 2774 2268 2778 2272
rect 2806 2268 2810 2272
rect 2766 2258 2770 2262
rect 2886 2338 2890 2342
rect 2854 2308 2858 2312
rect 2862 2308 2866 2312
rect 2854 2278 2858 2282
rect 2838 2248 2842 2252
rect 2846 2238 2850 2242
rect 2798 2228 2802 2232
rect 2790 2198 2794 2202
rect 2758 2178 2762 2182
rect 2774 2158 2778 2162
rect 2766 2088 2770 2092
rect 2766 2058 2770 2062
rect 2790 2148 2794 2152
rect 2790 2078 2794 2082
rect 2926 2388 2930 2392
rect 2982 2498 2986 2502
rect 3022 2538 3026 2542
rect 3086 2558 3090 2562
rect 3126 2547 3130 2551
rect 3190 2548 3194 2552
rect 3150 2528 3154 2532
rect 3046 2518 3050 2522
rect 3166 2518 3170 2522
rect 3182 2518 3186 2522
rect 3086 2508 3090 2512
rect 3046 2498 3050 2502
rect 3098 2503 3102 2507
rect 3105 2503 3109 2507
rect 3158 2498 3162 2502
rect 3070 2488 3074 2492
rect 3062 2468 3066 2472
rect 3198 2498 3202 2502
rect 3214 2698 3218 2702
rect 3278 2838 3282 2842
rect 3358 2888 3362 2892
rect 3342 2878 3346 2882
rect 3358 2878 3362 2882
rect 3326 2868 3330 2872
rect 3334 2858 3338 2862
rect 3342 2858 3346 2862
rect 3406 3128 3410 3132
rect 3702 4058 3706 4062
rect 3694 3918 3698 3922
rect 3702 3888 3706 3892
rect 3686 3858 3690 3862
rect 3662 3808 3666 3812
rect 3610 3803 3614 3807
rect 3617 3803 3621 3807
rect 3638 3768 3642 3772
rect 3686 3768 3690 3772
rect 3606 3758 3610 3762
rect 3678 3758 3682 3762
rect 3598 3738 3602 3742
rect 3590 3708 3594 3712
rect 3670 3748 3674 3752
rect 3614 3738 3618 3742
rect 3654 3728 3658 3732
rect 3662 3728 3666 3732
rect 3638 3698 3642 3702
rect 3550 3688 3554 3692
rect 3566 3688 3570 3692
rect 3630 3688 3634 3692
rect 3566 3668 3570 3672
rect 3566 3658 3570 3662
rect 3534 3528 3538 3532
rect 3542 3528 3546 3532
rect 3534 3478 3538 3482
rect 3542 3478 3546 3482
rect 3478 3368 3482 3372
rect 3534 3428 3538 3432
rect 3518 3398 3522 3402
rect 3574 3648 3578 3652
rect 3598 3638 3602 3642
rect 3582 3618 3586 3622
rect 3646 3608 3650 3612
rect 3610 3603 3614 3607
rect 3617 3603 3621 3607
rect 3582 3598 3586 3602
rect 3662 3688 3666 3692
rect 3766 4058 3770 4062
rect 3814 4268 3818 4272
rect 3886 4528 3890 4532
rect 3878 4488 3882 4492
rect 3838 4438 3842 4442
rect 3846 4428 3850 4432
rect 3830 4378 3834 4382
rect 3830 4338 3834 4342
rect 3862 4448 3866 4452
rect 3854 4398 3858 4402
rect 3854 4378 3858 4382
rect 3846 4268 3850 4272
rect 3822 4228 3826 4232
rect 3830 4228 3834 4232
rect 3814 4218 3818 4222
rect 3878 4458 3882 4462
rect 3998 4718 4002 4722
rect 4030 4718 4034 4722
rect 4006 4698 4010 4702
rect 4006 4678 4010 4682
rect 3958 4668 3962 4672
rect 3974 4668 3978 4672
rect 3926 4648 3930 4652
rect 3926 4628 3930 4632
rect 3942 4658 3946 4662
rect 3982 4658 3986 4662
rect 4006 4658 4010 4662
rect 3982 4648 3986 4652
rect 3942 4638 3946 4642
rect 3910 4618 3914 4622
rect 3934 4618 3938 4622
rect 3926 4558 3930 4562
rect 3902 4538 3906 4542
rect 3918 4528 3922 4532
rect 3974 4608 3978 4612
rect 3934 4508 3938 4512
rect 3902 4488 3906 4492
rect 3982 4548 3986 4552
rect 4166 4808 4170 4812
rect 4110 4778 4114 4782
rect 4158 4768 4162 4772
rect 4094 4718 4098 4722
rect 4110 4728 4114 4732
rect 4078 4688 4082 4692
rect 4054 4648 4058 4652
rect 4014 4568 4018 4572
rect 4006 4558 4010 4562
rect 3966 4508 3970 4512
rect 3950 4468 3954 4472
rect 3902 4448 3906 4452
rect 3910 4438 3914 4442
rect 3982 4528 3986 4532
rect 3974 4498 3978 4502
rect 3998 4468 4002 4472
rect 3934 4458 3938 4462
rect 3966 4458 3970 4462
rect 3926 4408 3930 4412
rect 3894 4348 3898 4352
rect 3918 4338 3922 4342
rect 3886 4328 3890 4332
rect 3894 4318 3898 4322
rect 3886 4308 3890 4312
rect 3926 4308 3930 4312
rect 3870 4278 3874 4282
rect 3862 4268 3866 4272
rect 3862 4258 3866 4262
rect 3878 4258 3882 4262
rect 3846 4208 3850 4212
rect 3854 4208 3858 4212
rect 3846 4188 3850 4192
rect 3846 4158 3850 4162
rect 3814 4128 3818 4132
rect 3878 4248 3882 4252
rect 3870 4218 3874 4222
rect 3798 4058 3802 4062
rect 3854 4058 3858 4062
rect 3758 4048 3762 4052
rect 3790 4048 3794 4052
rect 3806 4048 3810 4052
rect 3758 4038 3762 4042
rect 3838 4038 3842 4042
rect 3814 4028 3818 4032
rect 3718 3988 3722 3992
rect 3846 3978 3850 3982
rect 3854 3958 3858 3962
rect 3766 3948 3770 3952
rect 3814 3948 3818 3952
rect 3734 3908 3738 3912
rect 3758 3908 3762 3912
rect 3750 3878 3754 3882
rect 3710 3868 3714 3872
rect 3774 3868 3778 3872
rect 3718 3848 3722 3852
rect 3718 3798 3722 3802
rect 3710 3768 3714 3772
rect 3710 3748 3714 3752
rect 3718 3748 3722 3752
rect 3742 3748 3746 3752
rect 3750 3748 3754 3752
rect 3694 3708 3698 3712
rect 3694 3688 3698 3692
rect 3694 3658 3698 3662
rect 3694 3638 3698 3642
rect 3662 3578 3666 3582
rect 3598 3548 3602 3552
rect 3630 3548 3634 3552
rect 3574 3508 3578 3512
rect 3582 3478 3586 3482
rect 3638 3478 3642 3482
rect 3574 3468 3578 3472
rect 3622 3468 3626 3472
rect 3590 3448 3594 3452
rect 3638 3448 3642 3452
rect 3610 3403 3614 3407
rect 3617 3403 3621 3407
rect 3686 3538 3690 3542
rect 3670 3508 3674 3512
rect 3694 3508 3698 3512
rect 3662 3488 3666 3492
rect 3718 3708 3722 3712
rect 3718 3668 3722 3672
rect 3734 3608 3738 3612
rect 3790 3928 3794 3932
rect 3830 3928 3834 3932
rect 3806 3888 3810 3892
rect 3838 3878 3842 3882
rect 3782 3828 3786 3832
rect 3790 3798 3794 3802
rect 3822 3848 3826 3852
rect 3910 4298 3914 4302
rect 3942 4418 3946 4422
rect 4086 4638 4090 4642
rect 4078 4628 4082 4632
rect 4062 4578 4066 4582
rect 4030 4548 4034 4552
rect 4062 4528 4066 4532
rect 4014 4518 4018 4522
rect 4030 4478 4034 4482
rect 4014 4468 4018 4472
rect 4006 4408 4010 4412
rect 3966 4378 3970 4382
rect 3974 4358 3978 4362
rect 3966 4348 3970 4352
rect 3942 4338 3946 4342
rect 3958 4338 3962 4342
rect 4062 4478 4066 4482
rect 4046 4448 4050 4452
rect 4046 4418 4050 4422
rect 4030 4378 4034 4382
rect 4054 4408 4058 4412
rect 4030 4368 4034 4372
rect 4062 4398 4066 4402
rect 3990 4338 3994 4342
rect 4014 4338 4018 4342
rect 4022 4338 4026 4342
rect 4054 4338 4058 4342
rect 3974 4318 3978 4322
rect 4006 4308 4010 4312
rect 3990 4298 3994 4302
rect 3958 4288 3962 4292
rect 3934 4268 3938 4272
rect 3894 4248 3898 4252
rect 3918 4258 3922 4262
rect 3926 4248 3930 4252
rect 3950 4248 3954 4252
rect 4022 4268 4026 4272
rect 4046 4288 4050 4292
rect 4022 4248 4026 4252
rect 3982 4238 3986 4242
rect 3910 4228 3914 4232
rect 4014 4228 4018 4232
rect 3894 4208 3898 4212
rect 3950 4178 3954 4182
rect 3974 4178 3978 4182
rect 3998 4178 4002 4182
rect 3918 4168 3922 4172
rect 4006 4168 4010 4172
rect 3966 4158 3970 4162
rect 3974 4158 3978 4162
rect 3950 4148 3954 4152
rect 3966 4138 3970 4142
rect 3958 4118 3962 4122
rect 3982 4118 3986 4122
rect 3934 4088 3938 4092
rect 3950 4068 3954 4072
rect 3902 4058 3906 4062
rect 3878 3898 3882 3902
rect 3846 3828 3850 3832
rect 3862 3828 3866 3832
rect 3870 3828 3874 3832
rect 3814 3758 3818 3762
rect 3798 3748 3802 3752
rect 3766 3698 3770 3702
rect 3806 3747 3810 3751
rect 3830 3748 3834 3752
rect 3854 3738 3858 3742
rect 3870 3728 3874 3732
rect 3846 3718 3850 3722
rect 3878 3708 3882 3712
rect 3854 3688 3858 3692
rect 3854 3678 3858 3682
rect 3758 3638 3762 3642
rect 3750 3618 3754 3622
rect 3814 3668 3818 3672
rect 3830 3668 3834 3672
rect 3942 4028 3946 4032
rect 3926 3988 3930 3992
rect 3950 3978 3954 3982
rect 3934 3948 3938 3952
rect 3974 4058 3978 4062
rect 4006 4108 4010 4112
rect 3998 4068 4002 4072
rect 4014 4068 4018 4072
rect 4030 4088 4034 4092
rect 4114 4703 4118 4707
rect 4121 4703 4125 4707
rect 4150 4698 4154 4702
rect 4110 4678 4114 4682
rect 4134 4678 4138 4682
rect 4286 4868 4290 4872
rect 4366 4868 4370 4872
rect 4510 4868 4514 4872
rect 4574 4868 4578 4872
rect 5038 4868 5042 4872
rect 4246 4858 4250 4862
rect 4222 4818 4226 4822
rect 4198 4808 4202 4812
rect 4206 4788 4210 4792
rect 4190 4778 4194 4782
rect 4190 4748 4194 4752
rect 4190 4728 4194 4732
rect 4158 4688 4162 4692
rect 4174 4688 4178 4692
rect 4158 4678 4162 4682
rect 4190 4668 4194 4672
rect 4110 4658 4114 4662
rect 4150 4658 4154 4662
rect 4134 4628 4138 4632
rect 4150 4628 4154 4632
rect 4174 4658 4178 4662
rect 4166 4638 4170 4642
rect 4158 4618 4162 4622
rect 4094 4598 4098 4602
rect 4150 4598 4154 4602
rect 4110 4588 4114 4592
rect 4078 4558 4082 4562
rect 4094 4548 4098 4552
rect 4142 4578 4146 4582
rect 4126 4568 4130 4572
rect 4102 4508 4106 4512
rect 4086 4458 4090 4462
rect 4114 4503 4118 4507
rect 4121 4503 4125 4507
rect 4118 4478 4122 4482
rect 4102 4408 4106 4412
rect 4094 4388 4098 4392
rect 4110 4388 4114 4392
rect 4078 4358 4082 4362
rect 4078 4348 4082 4352
rect 4094 4348 4098 4352
rect 4246 4688 4250 4692
rect 4318 4828 4322 4832
rect 4358 4818 4362 4822
rect 4278 4758 4282 4762
rect 4318 4738 4322 4742
rect 4302 4698 4306 4702
rect 4278 4688 4282 4692
rect 4254 4668 4258 4672
rect 4262 4668 4266 4672
rect 4206 4638 4210 4642
rect 4206 4618 4210 4622
rect 4246 4618 4250 4622
rect 4190 4588 4194 4592
rect 4318 4678 4322 4682
rect 4326 4668 4330 4672
rect 4286 4638 4290 4642
rect 4278 4578 4282 4582
rect 4326 4638 4330 4642
rect 4358 4688 4362 4692
rect 4358 4668 4362 4672
rect 4350 4658 4354 4662
rect 4342 4638 4346 4642
rect 4358 4638 4362 4642
rect 4310 4628 4314 4632
rect 4294 4618 4298 4622
rect 4326 4578 4330 4582
rect 4278 4568 4282 4572
rect 4182 4548 4186 4552
rect 4214 4548 4218 4552
rect 4310 4548 4314 4552
rect 4270 4538 4274 4542
rect 4294 4538 4298 4542
rect 4214 4518 4218 4522
rect 4198 4498 4202 4502
rect 4166 4458 4170 4462
rect 4134 4388 4138 4392
rect 4142 4348 4146 4352
rect 4126 4318 4130 4322
rect 4142 4318 4146 4322
rect 4114 4303 4118 4307
rect 4121 4303 4125 4307
rect 4102 4298 4106 4302
rect 4070 4288 4074 4292
rect 4158 4448 4162 4452
rect 4158 4438 4162 4442
rect 4158 4408 4162 4412
rect 4166 4358 4170 4362
rect 4158 4328 4162 4332
rect 4166 4328 4170 4332
rect 4150 4298 4154 4302
rect 4158 4298 4162 4302
rect 4206 4448 4210 4452
rect 4254 4488 4258 4492
rect 4278 4458 4282 4462
rect 4278 4448 4282 4452
rect 4262 4408 4266 4412
rect 4278 4408 4282 4412
rect 4230 4388 4234 4392
rect 4246 4378 4250 4382
rect 4214 4368 4218 4372
rect 4230 4348 4234 4352
rect 4294 4478 4298 4482
rect 4294 4448 4298 4452
rect 4334 4438 4338 4442
rect 4606 4858 4610 4862
rect 4606 4848 4610 4852
rect 4558 4828 4562 4832
rect 4374 4698 4378 4702
rect 4446 4758 4450 4762
rect 4526 4758 4530 4762
rect 4542 4748 4546 4752
rect 4462 4728 4466 4732
rect 4446 4698 4450 4702
rect 4422 4688 4426 4692
rect 4382 4678 4386 4682
rect 4414 4678 4418 4682
rect 4406 4668 4410 4672
rect 4382 4658 4386 4662
rect 4390 4638 4394 4642
rect 4374 4628 4378 4632
rect 4438 4658 4442 4662
rect 4510 4728 4514 4732
rect 4486 4668 4490 4672
rect 4534 4738 4538 4742
rect 4574 4738 4578 4742
rect 4598 4728 4602 4732
rect 4582 4718 4586 4722
rect 4534 4708 4538 4712
rect 4526 4678 4530 4682
rect 4574 4668 4578 4672
rect 4510 4658 4514 4662
rect 4494 4648 4498 4652
rect 4414 4598 4418 4602
rect 4414 4578 4418 4582
rect 4382 4568 4386 4572
rect 4406 4568 4410 4572
rect 4550 4658 4554 4662
rect 4518 4628 4522 4632
rect 4446 4568 4450 4572
rect 4478 4548 4482 4552
rect 4558 4628 4562 4632
rect 4526 4608 4530 4612
rect 4566 4578 4570 4582
rect 4518 4568 4522 4572
rect 4542 4558 4546 4562
rect 4566 4558 4570 4562
rect 4510 4548 4514 4552
rect 4430 4538 4434 4542
rect 4494 4538 4498 4542
rect 4534 4538 4538 4542
rect 4542 4538 4546 4542
rect 4558 4538 4562 4542
rect 4366 4528 4370 4532
rect 4398 4528 4402 4532
rect 4454 4528 4458 4532
rect 4398 4518 4402 4522
rect 4486 4518 4490 4522
rect 4462 4498 4466 4502
rect 4454 4488 4458 4492
rect 4446 4468 4450 4472
rect 4390 4448 4394 4452
rect 4374 4378 4378 4382
rect 4310 4358 4314 4362
rect 4318 4358 4322 4362
rect 4326 4348 4330 4352
rect 4262 4338 4266 4342
rect 4382 4358 4386 4362
rect 4358 4348 4362 4352
rect 4374 4348 4378 4352
rect 4278 4328 4282 4332
rect 4286 4328 4290 4332
rect 4350 4328 4354 4332
rect 4278 4308 4282 4312
rect 4254 4278 4258 4282
rect 4174 4268 4178 4272
rect 4230 4268 4234 4272
rect 4270 4268 4274 4272
rect 4086 4258 4090 4262
rect 4206 4258 4210 4262
rect 4070 4248 4074 4252
rect 4078 4168 4082 4172
rect 4062 4148 4066 4152
rect 4086 4138 4090 4142
rect 4054 4108 4058 4112
rect 4062 4088 4066 4092
rect 4078 4088 4082 4092
rect 4070 4068 4074 4072
rect 4022 4038 4026 4042
rect 3998 3998 4002 4002
rect 3990 3978 3994 3982
rect 3974 3948 3978 3952
rect 3990 3948 3994 3952
rect 4022 3948 4026 3952
rect 3974 3938 3978 3942
rect 3958 3928 3962 3932
rect 3918 3918 3922 3922
rect 3982 3928 3986 3932
rect 3990 3928 3994 3932
rect 3974 3898 3978 3902
rect 3942 3868 3946 3872
rect 3982 3868 3986 3872
rect 3990 3858 3994 3862
rect 3902 3818 3906 3822
rect 3958 3818 3962 3822
rect 3950 3798 3954 3802
rect 3894 3778 3898 3782
rect 3998 3848 4002 3852
rect 3998 3838 4002 3842
rect 3990 3768 3994 3772
rect 3894 3748 3898 3752
rect 3966 3748 3970 3752
rect 3934 3728 3938 3732
rect 3918 3688 3922 3692
rect 3910 3668 3914 3672
rect 3942 3678 3946 3682
rect 3846 3658 3850 3662
rect 3870 3658 3874 3662
rect 3926 3658 3930 3662
rect 3854 3648 3858 3652
rect 3886 3638 3890 3642
rect 3942 3648 3946 3652
rect 3934 3608 3938 3612
rect 3774 3598 3778 3602
rect 3798 3598 3802 3602
rect 3902 3598 3906 3602
rect 3902 3568 3906 3572
rect 3750 3558 3754 3562
rect 3862 3558 3866 3562
rect 3910 3558 3914 3562
rect 3934 3558 3938 3562
rect 3942 3558 3946 3562
rect 3742 3548 3746 3552
rect 3838 3548 3842 3552
rect 3710 3498 3714 3502
rect 3678 3488 3682 3492
rect 3670 3468 3674 3472
rect 3662 3438 3666 3442
rect 3646 3398 3650 3402
rect 3614 3378 3618 3382
rect 3542 3368 3546 3372
rect 3566 3368 3570 3372
rect 3582 3368 3586 3372
rect 3598 3368 3602 3372
rect 3550 3358 3554 3362
rect 3574 3358 3578 3362
rect 3574 3348 3578 3352
rect 3566 3338 3570 3342
rect 3582 3338 3586 3342
rect 3486 3288 3490 3292
rect 3486 3278 3490 3282
rect 3502 3278 3506 3282
rect 3502 3258 3506 3262
rect 3438 3248 3442 3252
rect 3470 3248 3474 3252
rect 3430 3218 3434 3222
rect 3446 3158 3450 3162
rect 3470 3148 3474 3152
rect 3430 3138 3434 3142
rect 3462 3138 3466 3142
rect 3438 3128 3442 3132
rect 3398 3058 3402 3062
rect 3414 3038 3418 3042
rect 3446 3088 3450 3092
rect 3462 3078 3466 3082
rect 3478 3098 3482 3102
rect 3510 3228 3514 3232
rect 3550 3328 3554 3332
rect 3542 3298 3546 3302
rect 3534 3278 3538 3282
rect 3590 3318 3594 3322
rect 3558 3308 3562 3312
rect 3630 3348 3634 3352
rect 3654 3328 3658 3332
rect 3574 3298 3578 3302
rect 3542 3258 3546 3262
rect 3526 3218 3530 3222
rect 3542 3208 3546 3212
rect 3566 3178 3570 3182
rect 3582 3268 3586 3272
rect 3582 3238 3586 3242
rect 3574 3158 3578 3162
rect 3534 3138 3538 3142
rect 3582 3138 3586 3142
rect 3494 3088 3498 3092
rect 3470 3068 3474 3072
rect 3454 3058 3458 3062
rect 3494 3078 3498 3082
rect 3502 3068 3506 3072
rect 3526 3068 3530 3072
rect 3510 3058 3514 3062
rect 3518 3058 3522 3062
rect 3486 3048 3490 3052
rect 3502 3028 3506 3032
rect 3430 3018 3434 3022
rect 3406 3008 3410 3012
rect 3390 2958 3394 2962
rect 3462 2958 3466 2962
rect 3494 2948 3498 2952
rect 3542 3048 3546 3052
rect 3534 3038 3538 3042
rect 3582 3108 3586 3112
rect 3566 3068 3570 3072
rect 3574 3048 3578 3052
rect 3558 2998 3562 3002
rect 3566 2998 3570 3002
rect 3518 2978 3522 2982
rect 3534 2968 3538 2972
rect 3542 2958 3546 2962
rect 3430 2938 3434 2942
rect 3534 2938 3538 2942
rect 3398 2888 3402 2892
rect 3462 2888 3466 2892
rect 3478 2888 3482 2892
rect 3494 2888 3498 2892
rect 3446 2878 3450 2882
rect 3422 2868 3426 2872
rect 3518 2928 3522 2932
rect 3478 2868 3482 2872
rect 3510 2868 3514 2872
rect 3534 2918 3538 2922
rect 3614 3288 3618 3292
rect 3894 3548 3898 3552
rect 3926 3548 3930 3552
rect 3750 3538 3754 3542
rect 3790 3538 3794 3542
rect 3982 3738 3986 3742
rect 3974 3678 3978 3682
rect 4126 4208 4130 4212
rect 4114 4103 4118 4107
rect 4121 4103 4125 4107
rect 4046 4048 4050 4052
rect 4086 4048 4090 4052
rect 4046 3998 4050 4002
rect 4038 3908 4042 3912
rect 4238 4258 4242 4262
rect 4342 4318 4346 4322
rect 4366 4308 4370 4312
rect 4334 4288 4338 4292
rect 4286 4268 4290 4272
rect 4238 4248 4242 4252
rect 4222 4238 4226 4242
rect 4198 4228 4202 4232
rect 4158 4218 4162 4222
rect 4214 4178 4218 4182
rect 4190 4168 4194 4172
rect 4198 4168 4202 4172
rect 4150 4147 4154 4151
rect 4222 4168 4226 4172
rect 4238 4158 4242 4162
rect 4230 4148 4234 4152
rect 4246 4148 4250 4152
rect 4206 4128 4210 4132
rect 4262 4128 4266 4132
rect 4206 4108 4210 4112
rect 4190 4068 4194 4072
rect 4222 4068 4226 4072
rect 4238 4068 4242 4072
rect 4166 4048 4170 4052
rect 4150 4038 4154 4042
rect 4182 4038 4186 4042
rect 4150 4028 4154 4032
rect 4134 4018 4138 4022
rect 4126 3998 4130 4002
rect 4142 3998 4146 4002
rect 4118 3988 4122 3992
rect 4102 3978 4106 3982
rect 4110 3958 4114 3962
rect 4014 3858 4018 3862
rect 4022 3848 4026 3852
rect 4014 3818 4018 3822
rect 4006 3798 4010 3802
rect 3998 3698 4002 3702
rect 4014 3688 4018 3692
rect 3990 3668 3994 3672
rect 3990 3658 3994 3662
rect 3958 3618 3962 3622
rect 3958 3568 3962 3572
rect 3902 3528 3906 3532
rect 3942 3528 3946 3532
rect 3950 3528 3954 3532
rect 3750 3498 3754 3502
rect 3742 3448 3746 3452
rect 3718 3388 3722 3392
rect 3702 3368 3706 3372
rect 3814 3508 3818 3512
rect 3782 3478 3786 3482
rect 3806 3468 3810 3472
rect 3950 3518 3954 3522
rect 3902 3498 3906 3502
rect 3870 3478 3874 3482
rect 3910 3478 3914 3482
rect 3822 3468 3826 3472
rect 3894 3468 3898 3472
rect 3926 3458 3930 3462
rect 3766 3448 3770 3452
rect 3798 3448 3802 3452
rect 3846 3448 3850 3452
rect 3790 3438 3794 3442
rect 3910 3448 3914 3452
rect 3926 3448 3930 3452
rect 3982 3518 3986 3522
rect 3966 3508 3970 3512
rect 3966 3498 3970 3502
rect 4134 3948 4138 3952
rect 4118 3938 4122 3942
rect 4054 3888 4058 3892
rect 4062 3888 4066 3892
rect 4102 3918 4106 3922
rect 4114 3903 4118 3907
rect 4121 3903 4125 3907
rect 4134 3898 4138 3902
rect 4086 3878 4090 3882
rect 4134 3878 4138 3882
rect 4070 3858 4074 3862
rect 4102 3848 4106 3852
rect 4086 3818 4090 3822
rect 4126 3798 4130 3802
rect 4126 3758 4130 3762
rect 4054 3738 4058 3742
rect 4078 3738 4082 3742
rect 4118 3738 4122 3742
rect 4046 3678 4050 3682
rect 4070 3668 4074 3672
rect 4062 3658 4066 3662
rect 4006 3648 4010 3652
rect 4022 3588 4026 3592
rect 4094 3638 4098 3642
rect 4086 3628 4090 3632
rect 4114 3703 4118 3707
rect 4121 3703 4125 3707
rect 4190 4018 4194 4022
rect 4214 4018 4218 4022
rect 4278 4058 4282 4062
rect 4270 4018 4274 4022
rect 4318 4268 4322 4272
rect 4414 4458 4418 4462
rect 4462 4458 4466 4462
rect 4422 4448 4426 4452
rect 4414 4438 4418 4442
rect 4446 4408 4450 4412
rect 4430 4358 4434 4362
rect 4398 4258 4402 4262
rect 4318 4248 4322 4252
rect 4366 4248 4370 4252
rect 4438 4228 4442 4232
rect 4302 4218 4306 4222
rect 4438 4218 4442 4222
rect 4454 4338 4458 4342
rect 4358 4198 4362 4202
rect 4382 4198 4386 4202
rect 4446 4198 4450 4202
rect 4350 4158 4354 4162
rect 4286 4008 4290 4012
rect 4254 3998 4258 4002
rect 4262 3998 4266 4002
rect 4278 3988 4282 3992
rect 4166 3968 4170 3972
rect 4182 3968 4186 3972
rect 4150 3868 4154 3872
rect 4158 3858 4162 3862
rect 4174 3908 4178 3912
rect 4174 3898 4178 3902
rect 4190 3958 4194 3962
rect 4238 3958 4242 3962
rect 4198 3948 4202 3952
rect 4190 3918 4194 3922
rect 4198 3918 4202 3922
rect 4246 3948 4250 3952
rect 4222 3888 4226 3892
rect 4214 3878 4218 3882
rect 4166 3848 4170 3852
rect 4142 3838 4146 3842
rect 4174 3818 4178 3822
rect 4214 3858 4218 3862
rect 4254 3938 4258 3942
rect 4262 3938 4266 3942
rect 4238 3918 4242 3922
rect 4230 3878 4234 3882
rect 4254 3888 4258 3892
rect 4246 3868 4250 3872
rect 4302 4108 4306 4112
rect 4334 4108 4338 4112
rect 4318 4088 4322 4092
rect 4302 4068 4306 4072
rect 4318 4068 4322 4072
rect 4334 4058 4338 4062
rect 4310 4048 4314 4052
rect 4302 3948 4306 3952
rect 4510 4488 4514 4492
rect 4494 4468 4498 4472
rect 4518 4428 4522 4432
rect 4494 4418 4498 4422
rect 4518 4418 4522 4422
rect 4534 4418 4538 4422
rect 4518 4388 4522 4392
rect 4478 4358 4482 4362
rect 4502 4358 4506 4362
rect 4510 4358 4514 4362
rect 4502 4348 4506 4352
rect 4590 4638 4594 4642
rect 4678 4838 4682 4842
rect 4634 4803 4638 4807
rect 4641 4803 4645 4807
rect 4702 4858 4706 4862
rect 4862 4858 4866 4862
rect 4918 4858 4922 4862
rect 5030 4858 5034 4862
rect 4774 4848 4778 4852
rect 4846 4848 4850 4852
rect 4934 4848 4938 4852
rect 5070 4848 5074 4852
rect 5102 4848 5106 4852
rect 4750 4838 4754 4842
rect 5006 4838 5010 4842
rect 4686 4828 4690 4832
rect 4694 4818 4698 4822
rect 4814 4818 4818 4822
rect 4622 4788 4626 4792
rect 4622 4778 4626 4782
rect 4902 4808 4906 4812
rect 5038 4808 5042 4812
rect 5022 4798 5026 4802
rect 4750 4778 4754 4782
rect 4902 4778 4906 4782
rect 4622 4748 4626 4752
rect 4614 4708 4618 4712
rect 4638 4708 4642 4712
rect 4830 4768 4834 4772
rect 4854 4768 4858 4772
rect 4686 4748 4690 4752
rect 4838 4748 4842 4752
rect 4686 4698 4690 4702
rect 4654 4688 4658 4692
rect 4630 4668 4634 4672
rect 4678 4668 4682 4672
rect 4702 4668 4706 4672
rect 4638 4648 4642 4652
rect 4678 4648 4682 4652
rect 4606 4638 4610 4642
rect 4582 4618 4586 4622
rect 4598 4618 4602 4622
rect 4654 4638 4658 4642
rect 4678 4638 4682 4642
rect 4634 4603 4638 4607
rect 4641 4603 4645 4607
rect 4614 4568 4618 4572
rect 4630 4568 4634 4572
rect 4614 4558 4618 4562
rect 4590 4508 4594 4512
rect 4574 4478 4578 4482
rect 4582 4468 4586 4472
rect 4542 4408 4546 4412
rect 4550 4408 4554 4412
rect 4542 4398 4546 4402
rect 4494 4328 4498 4332
rect 4558 4328 4562 4332
rect 4478 4288 4482 4292
rect 4678 4578 4682 4582
rect 4606 4448 4610 4452
rect 4654 4438 4658 4442
rect 4606 4408 4610 4412
rect 4598 4358 4602 4362
rect 4634 4403 4638 4407
rect 4641 4403 4645 4407
rect 4686 4518 4690 4522
rect 4678 4488 4682 4492
rect 4694 4488 4698 4492
rect 4678 4468 4682 4472
rect 4710 4648 4714 4652
rect 4710 4608 4714 4612
rect 4862 4758 4866 4762
rect 4998 4758 5002 4762
rect 5014 4758 5018 4762
rect 4918 4748 4922 4752
rect 4982 4748 4986 4752
rect 4814 4718 4818 4722
rect 4862 4718 4866 4722
rect 4950 4718 4954 4722
rect 4862 4678 4866 4682
rect 4942 4678 4946 4682
rect 4814 4668 4818 4672
rect 4742 4658 4746 4662
rect 4790 4658 4794 4662
rect 4750 4648 4754 4652
rect 4774 4648 4778 4652
rect 4726 4568 4730 4572
rect 4742 4558 4746 4562
rect 4726 4538 4730 4542
rect 4710 4518 4714 4522
rect 4734 4518 4738 4522
rect 4670 4448 4674 4452
rect 4694 4438 4698 4442
rect 4718 4458 4722 4462
rect 4710 4438 4714 4442
rect 4782 4618 4786 4622
rect 4814 4638 4818 4642
rect 4814 4598 4818 4602
rect 4966 4698 4970 4702
rect 4846 4658 4850 4662
rect 4854 4658 4858 4662
rect 4870 4658 4874 4662
rect 4886 4658 4890 4662
rect 4838 4598 4842 4602
rect 4830 4588 4834 4592
rect 4798 4558 4802 4562
rect 4798 4547 4802 4551
rect 4846 4548 4850 4552
rect 4822 4528 4826 4532
rect 4862 4638 4866 4642
rect 4862 4588 4866 4592
rect 4878 4648 4882 4652
rect 4886 4638 4890 4642
rect 4894 4568 4898 4572
rect 4926 4568 4930 4572
rect 4902 4548 4906 4552
rect 4862 4528 4866 4532
rect 4854 4498 4858 4502
rect 4862 4498 4866 4502
rect 4854 4488 4858 4492
rect 4798 4478 4802 4482
rect 4814 4468 4818 4472
rect 4750 4458 4754 4462
rect 4806 4458 4810 4462
rect 4838 4458 4842 4462
rect 4846 4448 4850 4452
rect 4830 4438 4834 4442
rect 4814 4428 4818 4432
rect 4734 4408 4738 4412
rect 4702 4398 4706 4402
rect 4750 4398 4754 4402
rect 4694 4358 4698 4362
rect 4734 4358 4738 4362
rect 4638 4318 4642 4322
rect 4574 4308 4578 4312
rect 4566 4288 4570 4292
rect 4526 4278 4530 4282
rect 4494 4268 4498 4272
rect 4526 4268 4530 4272
rect 4462 4248 4466 4252
rect 4502 4258 4506 4262
rect 4486 4248 4490 4252
rect 4478 4238 4482 4242
rect 4494 4228 4498 4232
rect 4510 4228 4514 4232
rect 4462 4218 4466 4222
rect 4454 4178 4458 4182
rect 4478 4198 4482 4202
rect 4454 4168 4458 4172
rect 4422 4158 4426 4162
rect 4374 4148 4378 4152
rect 4398 4138 4402 4142
rect 4406 4128 4410 4132
rect 4422 4128 4426 4132
rect 4430 4128 4434 4132
rect 4486 4188 4490 4192
rect 4518 4208 4522 4212
rect 4558 4258 4562 4262
rect 4526 4178 4530 4182
rect 4566 4178 4570 4182
rect 4574 4158 4578 4162
rect 4542 4148 4546 4152
rect 4566 4148 4570 4152
rect 4534 4138 4538 4142
rect 4558 4138 4562 4142
rect 4478 4128 4482 4132
rect 4486 4128 4490 4132
rect 4510 4128 4514 4132
rect 4446 4118 4450 4122
rect 4414 4108 4418 4112
rect 4438 4088 4442 4092
rect 4430 4078 4434 4082
rect 4446 4068 4450 4072
rect 4390 4048 4394 4052
rect 4398 4048 4402 4052
rect 4558 4098 4562 4102
rect 4486 4068 4490 4072
rect 4478 4058 4482 4062
rect 4430 4038 4434 4042
rect 4446 4038 4450 4042
rect 4406 3998 4410 4002
rect 4350 3958 4354 3962
rect 4382 3958 4386 3962
rect 4398 3958 4402 3962
rect 4358 3948 4362 3952
rect 4374 3948 4378 3952
rect 4318 3938 4322 3942
rect 4390 3938 4394 3942
rect 4350 3928 4354 3932
rect 4334 3908 4338 3912
rect 4342 3908 4346 3912
rect 4198 3838 4202 3842
rect 4190 3808 4194 3812
rect 4254 3848 4258 3852
rect 4254 3828 4258 3832
rect 4238 3798 4242 3802
rect 4238 3768 4242 3772
rect 4222 3758 4226 3762
rect 4198 3748 4202 3752
rect 4150 3738 4154 3742
rect 4182 3678 4186 3682
rect 4206 3738 4210 3742
rect 4222 3688 4226 3692
rect 4150 3658 4154 3662
rect 4318 3848 4322 3852
rect 4326 3768 4330 3772
rect 4294 3758 4298 3762
rect 4310 3758 4314 3762
rect 4310 3748 4314 3752
rect 4262 3738 4266 3742
rect 4366 3898 4370 3902
rect 4414 3968 4418 3972
rect 4510 4028 4514 4032
rect 4526 4018 4530 4022
rect 4486 3988 4490 3992
rect 4478 3958 4482 3962
rect 4438 3948 4442 3952
rect 4462 3948 4466 3952
rect 4414 3928 4418 3932
rect 4670 4318 4674 4322
rect 4726 4318 4730 4322
rect 4662 4288 4666 4292
rect 4702 4308 4706 4312
rect 4782 4408 4786 4412
rect 4758 4378 4762 4382
rect 4766 4358 4770 4362
rect 4766 4348 4770 4352
rect 4758 4338 4762 4342
rect 4750 4328 4754 4332
rect 4798 4358 4802 4362
rect 4806 4358 4810 4362
rect 4782 4338 4786 4342
rect 4774 4318 4778 4322
rect 4790 4308 4794 4312
rect 4766 4298 4770 4302
rect 4742 4268 4746 4272
rect 4798 4278 4802 4282
rect 4622 4258 4626 4262
rect 4678 4258 4682 4262
rect 4622 4248 4626 4252
rect 4670 4248 4674 4252
rect 4694 4248 4698 4252
rect 4718 4238 4722 4242
rect 4630 4228 4634 4232
rect 4670 4218 4674 4222
rect 4838 4408 4842 4412
rect 4846 4378 4850 4382
rect 4822 4348 4826 4352
rect 4822 4298 4826 4302
rect 4814 4288 4818 4292
rect 4814 4268 4818 4272
rect 4830 4268 4834 4272
rect 4798 4258 4802 4262
rect 4878 4498 4882 4502
rect 4966 4538 4970 4542
rect 4990 4678 4994 4682
rect 4990 4648 4994 4652
rect 5038 4748 5042 4752
rect 5030 4718 5034 4722
rect 5126 4718 5130 4722
rect 5046 4668 5050 4672
rect 5022 4658 5026 4662
rect 5070 4658 5074 4662
rect 4998 4618 5002 4622
rect 5014 4618 5018 4622
rect 5030 4648 5034 4652
rect 4982 4548 4986 4552
rect 5054 4648 5058 4652
rect 5046 4628 5050 4632
rect 5046 4558 5050 4562
rect 4926 4528 4930 4532
rect 4974 4528 4978 4532
rect 4918 4488 4922 4492
rect 5070 4648 5074 4652
rect 5078 4628 5082 4632
rect 5078 4618 5082 4622
rect 5150 4848 5154 4852
rect 5150 4818 5154 4822
rect 5134 4668 5138 4672
rect 5126 4658 5130 4662
rect 5142 4618 5146 4622
rect 5094 4558 5098 4562
rect 5158 4558 5162 4562
rect 5174 4538 5178 4542
rect 5086 4508 5090 4512
rect 5062 4488 5066 4492
rect 5078 4488 5082 4492
rect 5022 4478 5026 4482
rect 5062 4478 5066 4482
rect 5078 4478 5082 4482
rect 4926 4468 4930 4472
rect 5094 4468 5098 4472
rect 4862 4428 4866 4432
rect 4862 4398 4866 4402
rect 4862 4358 4866 4362
rect 4918 4448 4922 4452
rect 4902 4418 4906 4422
rect 4990 4448 4994 4452
rect 4950 4418 4954 4422
rect 4966 4398 4970 4402
rect 4926 4368 4930 4372
rect 4934 4368 4938 4372
rect 4910 4358 4914 4362
rect 4878 4348 4882 4352
rect 4894 4348 4898 4352
rect 4854 4328 4858 4332
rect 4870 4328 4874 4332
rect 4862 4268 4866 4272
rect 4846 4258 4850 4262
rect 4782 4228 4786 4232
rect 4822 4218 4826 4222
rect 4854 4218 4858 4222
rect 4634 4203 4638 4207
rect 4641 4203 4645 4207
rect 4622 4148 4626 4152
rect 4654 4108 4658 4112
rect 4646 4098 4650 4102
rect 4582 4078 4586 4082
rect 4582 4058 4586 4062
rect 4606 4058 4610 4062
rect 4598 4028 4602 4032
rect 4566 3998 4570 4002
rect 4590 3998 4594 4002
rect 4534 3988 4538 3992
rect 4526 3968 4530 3972
rect 4502 3928 4506 3932
rect 4462 3888 4466 3892
rect 4478 3888 4482 3892
rect 4494 3888 4498 3892
rect 4398 3868 4402 3872
rect 4430 3868 4434 3872
rect 4374 3858 4378 3862
rect 4430 3858 4434 3862
rect 4462 3858 4466 3862
rect 4478 3858 4482 3862
rect 4486 3858 4490 3862
rect 4390 3848 4394 3852
rect 4422 3838 4426 3842
rect 4382 3828 4386 3832
rect 4358 3818 4362 3822
rect 4342 3758 4346 3762
rect 4286 3728 4290 3732
rect 4270 3698 4274 3702
rect 4270 3688 4274 3692
rect 4238 3668 4242 3672
rect 4254 3668 4258 3672
rect 4262 3658 4266 3662
rect 4254 3648 4258 3652
rect 4110 3628 4114 3632
rect 4094 3588 4098 3592
rect 4054 3568 4058 3572
rect 4078 3568 4082 3572
rect 4046 3548 4050 3552
rect 3998 3528 4002 3532
rect 3998 3508 4002 3512
rect 4094 3528 4098 3532
rect 4086 3518 4090 3522
rect 3990 3478 3994 3482
rect 4030 3459 4034 3463
rect 4190 3628 4194 3632
rect 4134 3598 4138 3602
rect 4118 3568 4122 3572
rect 4110 3528 4114 3532
rect 4114 3503 4118 3507
rect 4121 3503 4125 3507
rect 4102 3498 4106 3502
rect 4182 3568 4186 3572
rect 4206 3568 4210 3572
rect 4222 3568 4226 3572
rect 4158 3548 4162 3552
rect 4174 3548 4178 3552
rect 4142 3528 4146 3532
rect 4142 3518 4146 3522
rect 4094 3468 4098 3472
rect 4094 3458 4098 3462
rect 4150 3458 4154 3462
rect 3974 3448 3978 3452
rect 4094 3448 4098 3452
rect 4118 3448 4122 3452
rect 3910 3438 3914 3442
rect 3942 3438 3946 3442
rect 3902 3418 3906 3422
rect 3830 3408 3834 3412
rect 3830 3398 3834 3402
rect 3782 3388 3786 3392
rect 3678 3348 3682 3352
rect 3710 3348 3714 3352
rect 3718 3348 3722 3352
rect 3742 3348 3746 3352
rect 3734 3328 3738 3332
rect 3718 3308 3722 3312
rect 3598 3278 3602 3282
rect 3726 3268 3730 3272
rect 3654 3258 3658 3262
rect 3670 3248 3674 3252
rect 3686 3248 3690 3252
rect 3610 3203 3614 3207
rect 3617 3203 3621 3207
rect 3614 3148 3618 3152
rect 3622 3138 3626 3142
rect 3734 3248 3738 3252
rect 3694 3228 3698 3232
rect 3638 3188 3642 3192
rect 3630 3128 3634 3132
rect 3622 3078 3626 3082
rect 3590 3068 3594 3072
rect 3614 3068 3618 3072
rect 3646 3048 3650 3052
rect 3630 3038 3634 3042
rect 3582 2978 3586 2982
rect 3590 2947 3594 2951
rect 3630 3008 3634 3012
rect 3610 3003 3614 3007
rect 3617 3003 3621 3007
rect 3630 2988 3634 2992
rect 3614 2928 3618 2932
rect 3558 2868 3562 2872
rect 3502 2858 3506 2862
rect 3550 2858 3554 2862
rect 3366 2838 3370 2842
rect 3446 2848 3450 2852
rect 3310 2828 3314 2832
rect 3390 2828 3394 2832
rect 3398 2828 3402 2832
rect 3350 2808 3354 2812
rect 3286 2788 3290 2792
rect 3342 2788 3346 2792
rect 3286 2738 3290 2742
rect 3302 2698 3306 2702
rect 3334 2678 3338 2682
rect 3294 2648 3298 2652
rect 3318 2648 3322 2652
rect 3270 2578 3274 2582
rect 3222 2548 3226 2552
rect 3214 2528 3218 2532
rect 3334 2628 3338 2632
rect 3318 2588 3322 2592
rect 3374 2768 3378 2772
rect 3366 2728 3370 2732
rect 3358 2668 3362 2672
rect 3430 2748 3434 2752
rect 3430 2708 3434 2712
rect 3390 2668 3394 2672
rect 3382 2658 3386 2662
rect 3366 2648 3370 2652
rect 3430 2648 3434 2652
rect 3390 2638 3394 2642
rect 3358 2598 3362 2602
rect 3390 2568 3394 2572
rect 3382 2558 3386 2562
rect 3318 2548 3322 2552
rect 3326 2538 3330 2542
rect 3358 2538 3362 2542
rect 3374 2538 3378 2542
rect 3286 2528 3290 2532
rect 3294 2528 3298 2532
rect 3334 2528 3338 2532
rect 3326 2518 3330 2522
rect 3310 2508 3314 2512
rect 3350 2508 3354 2512
rect 3334 2498 3338 2502
rect 3206 2488 3210 2492
rect 3262 2488 3266 2492
rect 3278 2488 3282 2492
rect 3294 2488 3298 2492
rect 3126 2468 3130 2472
rect 3150 2468 3154 2472
rect 3174 2468 3178 2472
rect 3182 2468 3186 2472
rect 3246 2468 3250 2472
rect 3014 2458 3018 2462
rect 3038 2458 3042 2462
rect 3078 2458 3082 2462
rect 2990 2388 2994 2392
rect 3022 2448 3026 2452
rect 3062 2448 3066 2452
rect 3014 2408 3018 2412
rect 3022 2388 3026 2392
rect 2998 2368 3002 2372
rect 3014 2368 3018 2372
rect 2942 2348 2946 2352
rect 2958 2348 2962 2352
rect 2974 2348 2978 2352
rect 2886 2228 2890 2232
rect 2982 2338 2986 2342
rect 2958 2278 2962 2282
rect 3006 2278 3010 2282
rect 2974 2268 2978 2272
rect 3014 2268 3018 2272
rect 2918 2258 2922 2262
rect 2990 2258 2994 2262
rect 2942 2238 2946 2242
rect 2958 2228 2962 2232
rect 3006 2228 3010 2232
rect 2902 2218 2906 2222
rect 2926 2168 2930 2172
rect 2894 2158 2898 2162
rect 2966 2178 2970 2182
rect 2998 2168 3002 2172
rect 3006 2168 3010 2172
rect 3014 2168 3018 2172
rect 2982 2158 2986 2162
rect 2894 2148 2898 2152
rect 2910 2148 2914 2152
rect 2942 2148 2946 2152
rect 2950 2148 2954 2152
rect 2838 2138 2842 2142
rect 2886 2138 2890 2142
rect 2862 2128 2866 2132
rect 2878 2118 2882 2122
rect 2822 2088 2826 2092
rect 2830 2068 2834 2072
rect 2814 2058 2818 2062
rect 2862 2058 2866 2062
rect 2838 2048 2842 2052
rect 2862 2048 2866 2052
rect 2878 2048 2882 2052
rect 2910 2048 2914 2052
rect 2750 2038 2754 2042
rect 2758 2008 2762 2012
rect 2782 2008 2786 2012
rect 2830 2008 2834 2012
rect 2878 1978 2882 1982
rect 2814 1968 2818 1972
rect 2774 1958 2778 1962
rect 2870 1958 2874 1962
rect 2758 1948 2762 1952
rect 2838 1938 2842 1942
rect 2926 2138 2930 2142
rect 2974 2128 2978 2132
rect 2982 2118 2986 2122
rect 2934 2108 2938 2112
rect 2934 2078 2938 2082
rect 2990 2108 2994 2112
rect 3006 2108 3010 2112
rect 2926 2058 2930 2062
rect 3030 2328 3034 2332
rect 3054 2318 3058 2322
rect 3030 2308 3034 2312
rect 3046 2308 3050 2312
rect 3046 2258 3050 2262
rect 3086 2398 3090 2402
rect 3150 2458 3154 2462
rect 3198 2458 3202 2462
rect 3102 2448 3106 2452
rect 3142 2438 3146 2442
rect 3142 2418 3146 2422
rect 3094 2368 3098 2372
rect 3182 2438 3186 2442
rect 3206 2438 3210 2442
rect 3190 2408 3194 2412
rect 3206 2408 3210 2412
rect 3190 2398 3194 2402
rect 3166 2358 3170 2362
rect 3070 2338 3074 2342
rect 3174 2338 3178 2342
rect 3118 2308 3122 2312
rect 3098 2303 3102 2307
rect 3105 2303 3109 2307
rect 3070 2298 3074 2302
rect 3062 2278 3066 2282
rect 3070 2268 3074 2272
rect 3094 2268 3098 2272
rect 3062 2228 3066 2232
rect 3046 2188 3050 2192
rect 3030 2168 3034 2172
rect 3054 2158 3058 2162
rect 3054 2118 3058 2122
rect 3022 2078 3026 2082
rect 3102 2248 3106 2252
rect 3086 2238 3090 2242
rect 3078 2168 3082 2172
rect 3190 2268 3194 2272
rect 3142 2248 3146 2252
rect 3126 2218 3130 2222
rect 3134 2218 3138 2222
rect 3078 2148 3082 2152
rect 3110 2148 3114 2152
rect 3118 2148 3122 2152
rect 3078 2128 3082 2132
rect 3070 2068 3074 2072
rect 3030 2048 3034 2052
rect 3014 2038 3018 2042
rect 2998 1988 3002 1992
rect 2998 1968 3002 1972
rect 2990 1958 2994 1962
rect 2894 1948 2898 1952
rect 2910 1948 2914 1952
rect 2950 1948 2954 1952
rect 2966 1948 2970 1952
rect 2982 1948 2986 1952
rect 2886 1938 2890 1942
rect 2910 1938 2914 1942
rect 2806 1898 2810 1902
rect 2750 1888 2754 1892
rect 2790 1888 2794 1892
rect 2806 1878 2810 1882
rect 2798 1868 2802 1872
rect 2870 1868 2874 1872
rect 2886 1868 2890 1872
rect 2750 1828 2754 1832
rect 2734 1778 2738 1782
rect 2662 1758 2666 1762
rect 2718 1748 2722 1752
rect 2742 1748 2746 1752
rect 2710 1738 2714 1742
rect 2614 1708 2618 1712
rect 2670 1688 2674 1692
rect 2630 1678 2634 1682
rect 2646 1678 2650 1682
rect 2630 1558 2634 1562
rect 2638 1558 2642 1562
rect 2686 1658 2690 1662
rect 2734 1688 2738 1692
rect 2854 1848 2858 1852
rect 2838 1798 2842 1802
rect 2862 1748 2866 1752
rect 2814 1738 2818 1742
rect 2806 1718 2810 1722
rect 2782 1708 2786 1712
rect 2766 1688 2770 1692
rect 2750 1678 2754 1682
rect 2790 1668 2794 1672
rect 2734 1658 2738 1662
rect 2718 1648 2722 1652
rect 2726 1648 2730 1652
rect 2694 1608 2698 1612
rect 2750 1588 2754 1592
rect 2790 1578 2794 1582
rect 2782 1558 2786 1562
rect 2726 1548 2730 1552
rect 2622 1538 2626 1542
rect 2638 1538 2642 1542
rect 2638 1498 2642 1502
rect 2638 1468 2642 1472
rect 2670 1538 2674 1542
rect 2670 1498 2674 1502
rect 2662 1468 2666 1472
rect 2614 1458 2618 1462
rect 2646 1458 2650 1462
rect 2654 1448 2658 1452
rect 2574 1428 2578 1432
rect 2606 1428 2610 1432
rect 2654 1428 2658 1432
rect 2486 1408 2490 1412
rect 2470 1388 2474 1392
rect 2478 1368 2482 1372
rect 2558 1368 2562 1372
rect 2422 1348 2426 1352
rect 2438 1348 2442 1352
rect 2470 1338 2474 1342
rect 2478 1338 2482 1342
rect 2494 1338 2498 1342
rect 2510 1338 2514 1342
rect 2454 1328 2458 1332
rect 2462 1288 2466 1292
rect 2414 1258 2418 1262
rect 2390 1218 2394 1222
rect 2374 1168 2378 1172
rect 2414 1208 2418 1212
rect 2430 1258 2434 1262
rect 2446 1238 2450 1242
rect 2406 1168 2410 1172
rect 2454 1178 2458 1182
rect 2422 1168 2426 1172
rect 2446 1158 2450 1162
rect 2430 1148 2434 1152
rect 2406 1138 2410 1142
rect 2342 1128 2346 1132
rect 2286 1058 2290 1062
rect 2254 1038 2258 1042
rect 2278 1038 2282 1042
rect 2286 1008 2290 1012
rect 2230 948 2234 952
rect 2182 938 2186 942
rect 2174 928 2178 932
rect 2166 908 2170 912
rect 2126 868 2130 872
rect 2142 868 2146 872
rect 2134 848 2138 852
rect 2126 808 2130 812
rect 2094 788 2098 792
rect 1926 748 1930 752
rect 2030 748 2034 752
rect 1942 738 1946 742
rect 1974 738 1978 742
rect 1966 728 1970 732
rect 1958 708 1962 712
rect 1902 668 1906 672
rect 1942 668 1946 672
rect 1902 658 1906 662
rect 1918 648 1922 652
rect 1862 558 1866 562
rect 1886 578 1890 582
rect 1830 538 1834 542
rect 1798 508 1802 512
rect 1822 488 1826 492
rect 1846 478 1850 482
rect 1574 368 1578 372
rect 1654 368 1658 372
rect 1662 368 1666 372
rect 1750 368 1754 372
rect 1758 368 1762 372
rect 1766 368 1770 372
rect 1566 358 1570 362
rect 1670 358 1674 362
rect 1694 358 1698 362
rect 1734 358 1738 362
rect 1710 338 1714 342
rect 1734 338 1738 342
rect 1750 338 1754 342
rect 1606 328 1610 332
rect 1606 308 1610 312
rect 1606 288 1610 292
rect 1582 278 1586 282
rect 1550 268 1554 272
rect 1598 268 1602 272
rect 1598 238 1602 242
rect 1582 228 1586 232
rect 1614 238 1618 242
rect 1606 218 1610 222
rect 1562 203 1566 207
rect 1569 203 1573 207
rect 1550 188 1554 192
rect 1726 278 1730 282
rect 1662 268 1666 272
rect 1630 248 1634 252
rect 1766 318 1770 322
rect 1854 468 1858 472
rect 1926 558 1930 562
rect 1902 548 1906 552
rect 1878 528 1882 532
rect 1998 718 2002 722
rect 1990 688 1994 692
rect 1974 678 1978 682
rect 2006 708 2010 712
rect 2014 708 2018 712
rect 2006 668 2010 672
rect 1950 648 1954 652
rect 1966 638 1970 642
rect 1982 628 1986 632
rect 2030 688 2034 692
rect 2126 758 2130 762
rect 2126 748 2130 752
rect 2214 928 2218 932
rect 2206 898 2210 902
rect 2254 918 2258 922
rect 2262 918 2266 922
rect 2222 888 2226 892
rect 2278 888 2282 892
rect 2254 878 2258 882
rect 2190 748 2194 752
rect 2166 738 2170 742
rect 2094 728 2098 732
rect 2150 728 2154 732
rect 2054 708 2058 712
rect 2074 703 2078 707
rect 2081 703 2085 707
rect 2174 698 2178 702
rect 2126 688 2130 692
rect 2038 678 2042 682
rect 2086 678 2090 682
rect 2126 678 2130 682
rect 2038 658 2042 662
rect 2022 578 2026 582
rect 2022 568 2026 572
rect 2006 558 2010 562
rect 2014 558 2018 562
rect 2070 648 2074 652
rect 2054 638 2058 642
rect 2086 638 2090 642
rect 2046 578 2050 582
rect 2030 548 2034 552
rect 1990 538 1994 542
rect 1934 518 1938 522
rect 1966 528 1970 532
rect 1886 478 1890 482
rect 1934 468 1938 472
rect 1878 428 1882 432
rect 1910 418 1914 422
rect 2014 518 2018 522
rect 1990 488 1994 492
rect 2006 478 2010 482
rect 2094 568 2098 572
rect 2054 558 2058 562
rect 2118 558 2122 562
rect 2270 858 2274 862
rect 2262 828 2266 832
rect 2254 808 2258 812
rect 2238 758 2242 762
rect 2334 1048 2338 1052
rect 2294 998 2298 1002
rect 2406 1118 2410 1122
rect 2406 1098 2410 1102
rect 2390 1088 2394 1092
rect 2382 1078 2386 1082
rect 2462 1168 2466 1172
rect 2470 1158 2474 1162
rect 2438 1068 2442 1072
rect 2382 1048 2386 1052
rect 2406 1048 2410 1052
rect 2430 1038 2434 1042
rect 2414 1028 2418 1032
rect 2406 998 2410 1002
rect 2382 958 2386 962
rect 2326 948 2330 952
rect 2342 948 2346 952
rect 2350 938 2354 942
rect 2390 928 2394 932
rect 2350 918 2354 922
rect 2366 918 2370 922
rect 2310 898 2314 902
rect 2318 888 2322 892
rect 2302 858 2306 862
rect 2342 858 2346 862
rect 2326 808 2330 812
rect 2342 808 2346 812
rect 2318 798 2322 802
rect 2406 888 2410 892
rect 2470 1108 2474 1112
rect 2462 1048 2466 1052
rect 2446 1038 2450 1042
rect 2510 1328 2514 1332
rect 2534 1328 2538 1332
rect 2534 1278 2538 1282
rect 2526 1128 2530 1132
rect 2502 1058 2506 1062
rect 2502 1048 2506 1052
rect 2518 1028 2522 1032
rect 2486 988 2490 992
rect 2454 968 2458 972
rect 2486 958 2490 962
rect 2462 948 2466 952
rect 2454 938 2458 942
rect 2438 928 2442 932
rect 2438 918 2442 922
rect 2438 878 2442 882
rect 2550 1338 2554 1342
rect 2566 1328 2570 1332
rect 2586 1403 2590 1407
rect 2593 1403 2597 1407
rect 2606 1378 2610 1382
rect 2630 1368 2634 1372
rect 2606 1358 2610 1362
rect 2638 1358 2642 1362
rect 2614 1338 2618 1342
rect 2646 1338 2650 1342
rect 2590 1288 2594 1292
rect 2574 1268 2578 1272
rect 2574 1248 2578 1252
rect 2614 1248 2618 1252
rect 2566 1218 2570 1222
rect 2550 1208 2554 1212
rect 2550 1078 2554 1082
rect 2542 1068 2546 1072
rect 2606 1228 2610 1232
rect 2586 1203 2590 1207
rect 2593 1203 2597 1207
rect 2646 1298 2650 1302
rect 2630 1278 2634 1282
rect 2654 1238 2658 1242
rect 2734 1508 2738 1512
rect 2702 1488 2706 1492
rect 2678 1458 2682 1462
rect 2686 1438 2690 1442
rect 2678 1408 2682 1412
rect 2670 1358 2674 1362
rect 2662 1218 2666 1222
rect 2638 1198 2642 1202
rect 2702 1428 2706 1432
rect 2686 1368 2690 1372
rect 2734 1368 2738 1372
rect 2718 1358 2722 1362
rect 2694 1348 2698 1352
rect 2726 1348 2730 1352
rect 2734 1338 2738 1342
rect 2702 1308 2706 1312
rect 2822 1698 2826 1702
rect 2782 1528 2786 1532
rect 2790 1508 2794 1512
rect 2774 1468 2778 1472
rect 2758 1458 2762 1462
rect 2782 1358 2786 1362
rect 2750 1298 2754 1302
rect 2686 1288 2690 1292
rect 2702 1288 2706 1292
rect 2854 1698 2858 1702
rect 2910 1868 2914 1872
rect 2958 1938 2962 1942
rect 2926 1888 2930 1892
rect 2918 1848 2922 1852
rect 2902 1838 2906 1842
rect 2934 1778 2938 1782
rect 2934 1768 2938 1772
rect 2910 1758 2914 1762
rect 2942 1758 2946 1762
rect 2918 1748 2922 1752
rect 2958 1758 2962 1762
rect 2974 1848 2978 1852
rect 3006 1868 3010 1872
rect 3038 2008 3042 2012
rect 3046 1988 3050 1992
rect 3030 1978 3034 1982
rect 3038 1948 3042 1952
rect 3030 1898 3034 1902
rect 3022 1878 3026 1882
rect 3030 1868 3034 1872
rect 3022 1848 3026 1852
rect 3038 1848 3042 1852
rect 3014 1828 3018 1832
rect 3022 1828 3026 1832
rect 3062 2008 3066 2012
rect 3118 2128 3122 2132
rect 3098 2103 3102 2107
rect 3105 2103 3109 2107
rect 3158 2238 3162 2242
rect 3134 2128 3138 2132
rect 3166 2128 3170 2132
rect 3142 2108 3146 2112
rect 3190 2108 3194 2112
rect 3174 2098 3178 2102
rect 3118 2068 3122 2072
rect 3094 2058 3098 2062
rect 3118 2048 3122 2052
rect 3102 2008 3106 2012
rect 3086 1978 3090 1982
rect 3110 1948 3114 1952
rect 3054 1928 3058 1932
rect 3062 1908 3066 1912
rect 3054 1878 3058 1882
rect 3078 1898 3082 1902
rect 3098 1903 3102 1907
rect 3105 1903 3109 1907
rect 3086 1848 3090 1852
rect 3102 1848 3106 1852
rect 3110 1838 3114 1842
rect 3078 1828 3082 1832
rect 3102 1788 3106 1792
rect 3014 1778 3018 1782
rect 3046 1778 3050 1782
rect 3062 1778 3066 1782
rect 2982 1758 2986 1762
rect 2990 1758 2994 1762
rect 3070 1758 3074 1762
rect 2966 1748 2970 1752
rect 2990 1748 2994 1752
rect 2886 1728 2890 1732
rect 2942 1708 2946 1712
rect 2870 1678 2874 1682
rect 2982 1728 2986 1732
rect 3014 1728 3018 1732
rect 3022 1728 3026 1732
rect 2966 1698 2970 1702
rect 2974 1688 2978 1692
rect 2958 1678 2962 1682
rect 2910 1658 2914 1662
rect 2878 1648 2882 1652
rect 2838 1608 2842 1612
rect 2822 1528 2826 1532
rect 2814 1498 2818 1502
rect 2846 1558 2850 1562
rect 2998 1708 3002 1712
rect 3030 1708 3034 1712
rect 3062 1748 3066 1752
rect 3062 1728 3066 1732
rect 3098 1703 3102 1707
rect 3105 1703 3109 1707
rect 3110 1688 3114 1692
rect 3046 1678 3050 1682
rect 3070 1678 3074 1682
rect 3062 1668 3066 1672
rect 2990 1658 2994 1662
rect 3006 1658 3010 1662
rect 2942 1618 2946 1622
rect 2982 1618 2986 1622
rect 2926 1578 2930 1582
rect 2870 1558 2874 1562
rect 2870 1548 2874 1552
rect 2958 1548 2962 1552
rect 2870 1538 2874 1542
rect 2910 1538 2914 1542
rect 2926 1528 2930 1532
rect 2886 1518 2890 1522
rect 2902 1508 2906 1512
rect 2854 1498 2858 1502
rect 2870 1498 2874 1502
rect 2870 1488 2874 1492
rect 2846 1468 2850 1472
rect 2822 1458 2826 1462
rect 2798 1448 2802 1452
rect 3038 1648 3042 1652
rect 3062 1648 3066 1652
rect 3022 1608 3026 1612
rect 3142 2078 3146 2082
rect 3182 2068 3186 2072
rect 3142 2058 3146 2062
rect 3174 2048 3178 2052
rect 3158 1978 3162 1982
rect 3166 1978 3170 1982
rect 3142 1958 3146 1962
rect 3158 1938 3162 1942
rect 3142 1898 3146 1902
rect 3134 1888 3138 1892
rect 3134 1868 3138 1872
rect 3174 1868 3178 1872
rect 3150 1858 3154 1862
rect 3134 1848 3138 1852
rect 3150 1848 3154 1852
rect 3126 1778 3130 1782
rect 3206 2298 3210 2302
rect 3254 2458 3258 2462
rect 3270 2458 3274 2462
rect 3222 2448 3226 2452
rect 3238 2448 3242 2452
rect 3310 2458 3314 2462
rect 3342 2458 3346 2462
rect 3310 2448 3314 2452
rect 3270 2438 3274 2442
rect 3286 2438 3290 2442
rect 3318 2438 3322 2442
rect 3278 2408 3282 2412
rect 3254 2398 3258 2402
rect 3294 2398 3298 2402
rect 3270 2378 3274 2382
rect 3230 2358 3234 2362
rect 3254 2358 3258 2362
rect 3262 2358 3266 2362
rect 3230 2338 3234 2342
rect 3238 2328 3242 2332
rect 3246 2328 3250 2332
rect 3334 2398 3338 2402
rect 3310 2358 3314 2362
rect 3326 2358 3330 2362
rect 3334 2358 3338 2362
rect 3302 2348 3306 2352
rect 3358 2488 3362 2492
rect 3366 2398 3370 2402
rect 3366 2388 3370 2392
rect 3358 2348 3362 2352
rect 3310 2338 3314 2342
rect 3278 2328 3282 2332
rect 3262 2308 3266 2312
rect 3318 2308 3322 2312
rect 3326 2308 3330 2312
rect 3238 2298 3242 2302
rect 3230 2278 3234 2282
rect 3310 2278 3314 2282
rect 3302 2268 3306 2272
rect 3222 2188 3226 2192
rect 3262 2248 3266 2252
rect 3302 2238 3306 2242
rect 3294 2228 3298 2232
rect 3262 2158 3266 2162
rect 3478 2838 3482 2842
rect 3510 2838 3514 2842
rect 3462 2798 3466 2802
rect 3494 2788 3498 2792
rect 3526 2808 3530 2812
rect 3550 2768 3554 2772
rect 3470 2748 3474 2752
rect 3486 2748 3490 2752
rect 3518 2748 3522 2752
rect 3494 2738 3498 2742
rect 3534 2738 3538 2742
rect 3542 2728 3546 2732
rect 3526 2718 3530 2722
rect 3518 2668 3522 2672
rect 3558 2708 3562 2712
rect 3558 2698 3562 2702
rect 3486 2658 3490 2662
rect 3478 2648 3482 2652
rect 3462 2628 3466 2632
rect 3454 2548 3458 2552
rect 3574 2848 3578 2852
rect 3574 2818 3578 2822
rect 3582 2768 3586 2772
rect 3606 2888 3610 2892
rect 3782 3338 3786 3342
rect 3766 3328 3770 3332
rect 3878 3378 3882 3382
rect 3838 3348 3842 3352
rect 3862 3338 3866 3342
rect 3886 3338 3890 3342
rect 3822 3328 3826 3332
rect 3806 3308 3810 3312
rect 3846 3308 3850 3312
rect 3790 3298 3794 3302
rect 3766 3288 3770 3292
rect 3750 3268 3754 3272
rect 3902 3328 3906 3332
rect 3798 3268 3802 3272
rect 3790 3248 3794 3252
rect 3806 3248 3810 3252
rect 3766 3238 3770 3242
rect 3814 3238 3818 3242
rect 3846 3228 3850 3232
rect 3750 3218 3754 3222
rect 3742 3208 3746 3212
rect 3694 3178 3698 3182
rect 3694 3148 3698 3152
rect 3814 3198 3818 3202
rect 3766 3168 3770 3172
rect 3790 3168 3794 3172
rect 3822 3168 3826 3172
rect 3902 3248 3906 3252
rect 3878 3158 3882 3162
rect 3886 3158 3890 3162
rect 3806 3138 3810 3142
rect 3742 3128 3746 3132
rect 3734 3118 3738 3122
rect 3718 3078 3722 3082
rect 3750 3078 3754 3082
rect 3686 3058 3690 3062
rect 3686 3048 3690 3052
rect 3830 3138 3834 3142
rect 3814 3118 3818 3122
rect 3846 3098 3850 3102
rect 3830 3088 3834 3092
rect 3814 3078 3818 3082
rect 3774 3068 3778 3072
rect 3798 3068 3802 3072
rect 3870 3098 3874 3102
rect 3862 3068 3866 3072
rect 3894 3148 3898 3152
rect 3902 3098 3906 3102
rect 3854 3058 3858 3062
rect 3990 3438 3994 3442
rect 3966 3408 3970 3412
rect 3974 3408 3978 3412
rect 4086 3438 4090 3442
rect 4142 3438 4146 3442
rect 4174 3438 4178 3442
rect 4006 3408 4010 3412
rect 4070 3408 4074 3412
rect 3942 3378 3946 3382
rect 4102 3398 4106 3402
rect 3974 3368 3978 3372
rect 4070 3368 4074 3372
rect 4174 3368 4178 3372
rect 4206 3538 4210 3542
rect 4230 3538 4234 3542
rect 4198 3468 4202 3472
rect 4206 3458 4210 3462
rect 4198 3428 4202 3432
rect 4214 3408 4218 3412
rect 4206 3378 4210 3382
rect 4086 3358 4090 3362
rect 4190 3358 4194 3362
rect 3966 3348 3970 3352
rect 4166 3348 4170 3352
rect 4182 3348 4186 3352
rect 3926 3338 3930 3342
rect 3958 3338 3962 3342
rect 4030 3338 4034 3342
rect 4070 3338 4074 3342
rect 3990 3298 3994 3302
rect 3966 3268 3970 3272
rect 3990 3268 3994 3272
rect 3998 3258 4002 3262
rect 4062 3328 4066 3332
rect 4150 3328 4154 3332
rect 4158 3328 4162 3332
rect 4102 3318 4106 3322
rect 4118 3318 4122 3322
rect 4114 3303 4118 3307
rect 4121 3303 4125 3307
rect 4134 3298 4138 3302
rect 4046 3288 4050 3292
rect 4022 3278 4026 3282
rect 4054 3258 4058 3262
rect 4110 3258 4114 3262
rect 3974 3248 3978 3252
rect 4022 3248 4026 3252
rect 3934 3218 3938 3222
rect 3950 3208 3954 3212
rect 3950 3188 3954 3192
rect 3982 3188 3986 3192
rect 3926 3148 3930 3152
rect 3958 3148 3962 3152
rect 3926 3078 3930 3082
rect 3974 3118 3978 3122
rect 3982 3108 3986 3112
rect 3934 3068 3938 3072
rect 3990 3068 3994 3072
rect 3918 3058 3922 3062
rect 3950 3058 3954 3062
rect 3910 3038 3914 3042
rect 3886 3028 3890 3032
rect 3894 3028 3898 3032
rect 3774 3008 3778 3012
rect 3766 2998 3770 3002
rect 3718 2978 3722 2982
rect 3758 2978 3762 2982
rect 3678 2968 3682 2972
rect 3726 2958 3730 2962
rect 3686 2948 3690 2952
rect 3710 2948 3714 2952
rect 3726 2948 3730 2952
rect 3686 2938 3690 2942
rect 3702 2938 3706 2942
rect 3670 2888 3674 2892
rect 3654 2878 3658 2882
rect 3610 2803 3614 2807
rect 3617 2803 3621 2807
rect 3654 2818 3658 2822
rect 3638 2768 3642 2772
rect 3622 2758 3626 2762
rect 3590 2718 3594 2722
rect 3582 2678 3586 2682
rect 3598 2668 3602 2672
rect 3606 2658 3610 2662
rect 3566 2648 3570 2652
rect 3590 2628 3594 2632
rect 3566 2608 3570 2612
rect 3610 2603 3614 2607
rect 3617 2603 3621 2607
rect 3598 2598 3602 2602
rect 3534 2588 3538 2592
rect 3542 2588 3546 2592
rect 3526 2568 3530 2572
rect 3494 2558 3498 2562
rect 3518 2558 3522 2562
rect 3486 2548 3490 2552
rect 3486 2538 3490 2542
rect 3462 2528 3466 2532
rect 3430 2518 3434 2522
rect 3390 2508 3394 2512
rect 3398 2498 3402 2502
rect 3446 2478 3450 2482
rect 3414 2458 3418 2462
rect 3390 2438 3394 2442
rect 3382 2428 3386 2432
rect 3374 2368 3378 2372
rect 3398 2388 3402 2392
rect 3422 2448 3426 2452
rect 3414 2438 3418 2442
rect 3406 2378 3410 2382
rect 3382 2348 3386 2352
rect 3366 2338 3370 2342
rect 3374 2328 3378 2332
rect 3326 2298 3330 2302
rect 3334 2298 3338 2302
rect 3350 2298 3354 2302
rect 3382 2298 3386 2302
rect 3398 2298 3402 2302
rect 3334 2268 3338 2272
rect 3326 2258 3330 2262
rect 3342 2258 3346 2262
rect 3350 2258 3354 2262
rect 3406 2258 3410 2262
rect 3326 2228 3330 2232
rect 3326 2198 3330 2202
rect 3270 2148 3274 2152
rect 3310 2148 3314 2152
rect 3358 2248 3362 2252
rect 3366 2248 3370 2252
rect 3398 2248 3402 2252
rect 3438 2458 3442 2462
rect 3438 2448 3442 2452
rect 3470 2508 3474 2512
rect 3462 2488 3466 2492
rect 3478 2488 3482 2492
rect 3486 2488 3490 2492
rect 3462 2478 3466 2482
rect 3430 2408 3434 2412
rect 3422 2388 3426 2392
rect 3462 2368 3466 2372
rect 3422 2328 3426 2332
rect 3462 2238 3466 2242
rect 3446 2208 3450 2212
rect 3470 2208 3474 2212
rect 3414 2198 3418 2202
rect 3382 2178 3386 2182
rect 3398 2168 3402 2172
rect 3358 2148 3362 2152
rect 3406 2148 3410 2152
rect 3350 2138 3354 2142
rect 3302 2128 3306 2132
rect 3222 2118 3226 2122
rect 3270 2118 3274 2122
rect 3278 2108 3282 2112
rect 3326 2108 3330 2112
rect 3254 2088 3258 2092
rect 3206 2068 3210 2072
rect 3198 2028 3202 2032
rect 3222 1958 3226 1962
rect 3230 1938 3234 1942
rect 3230 1898 3234 1902
rect 3438 2168 3442 2172
rect 3502 2548 3506 2552
rect 3518 2548 3522 2552
rect 3550 2558 3554 2562
rect 3566 2558 3570 2562
rect 3542 2498 3546 2502
rect 3510 2458 3514 2462
rect 3534 2458 3538 2462
rect 3510 2388 3514 2392
rect 3494 2348 3498 2352
rect 3502 2298 3506 2302
rect 3494 2248 3498 2252
rect 3502 2248 3506 2252
rect 3478 2198 3482 2202
rect 3590 2488 3594 2492
rect 3646 2728 3650 2732
rect 3646 2678 3650 2682
rect 3638 2628 3642 2632
rect 3662 2758 3666 2762
rect 3662 2718 3666 2722
rect 3694 2868 3698 2872
rect 3694 2848 3698 2852
rect 3750 2908 3754 2912
rect 3782 2958 3786 2962
rect 3822 2958 3826 2962
rect 3838 2958 3842 2962
rect 3790 2948 3794 2952
rect 3822 2948 3826 2952
rect 3750 2858 3754 2862
rect 3766 2858 3770 2862
rect 3694 2738 3698 2742
rect 3678 2728 3682 2732
rect 3686 2728 3690 2732
rect 3694 2728 3698 2732
rect 3678 2688 3682 2692
rect 3654 2618 3658 2622
rect 3630 2568 3634 2572
rect 3646 2548 3650 2552
rect 3670 2678 3674 2682
rect 3678 2668 3682 2672
rect 3670 2658 3674 2662
rect 3694 2658 3698 2662
rect 3694 2628 3698 2632
rect 3670 2608 3674 2612
rect 3646 2538 3650 2542
rect 3678 2588 3682 2592
rect 3678 2578 3682 2582
rect 3718 2838 3722 2842
rect 3726 2768 3730 2772
rect 3710 2698 3714 2702
rect 3718 2678 3722 2682
rect 3758 2708 3762 2712
rect 3742 2678 3746 2682
rect 3726 2668 3730 2672
rect 3878 2947 3882 2951
rect 3854 2928 3858 2932
rect 3886 2888 3890 2892
rect 3830 2868 3834 2872
rect 3806 2858 3810 2862
rect 3846 2858 3850 2862
rect 3886 2858 3890 2862
rect 3870 2848 3874 2852
rect 3942 3048 3946 3052
rect 3934 3008 3938 3012
rect 3950 3038 3954 3042
rect 3974 2988 3978 2992
rect 3934 2958 3938 2962
rect 3958 2958 3962 2962
rect 3910 2868 3914 2872
rect 3918 2858 3922 2862
rect 3782 2838 3786 2842
rect 3822 2838 3826 2842
rect 3894 2838 3898 2842
rect 3830 2768 3834 2772
rect 3854 2768 3858 2772
rect 3886 2768 3890 2772
rect 3878 2758 3882 2762
rect 3782 2748 3786 2752
rect 3790 2747 3794 2751
rect 3854 2748 3858 2752
rect 3790 2738 3794 2742
rect 3830 2738 3834 2742
rect 3902 2808 3906 2812
rect 3910 2798 3914 2802
rect 3910 2768 3914 2772
rect 3910 2748 3914 2752
rect 3862 2738 3866 2742
rect 3870 2728 3874 2732
rect 3846 2718 3850 2722
rect 3782 2708 3786 2712
rect 3886 2708 3890 2712
rect 3806 2688 3810 2692
rect 3798 2678 3802 2682
rect 3774 2668 3778 2672
rect 3782 2658 3786 2662
rect 3894 2678 3898 2682
rect 3846 2658 3850 2662
rect 3790 2638 3794 2642
rect 3806 2638 3810 2642
rect 3718 2618 3722 2622
rect 3790 2618 3794 2622
rect 3750 2608 3754 2612
rect 3742 2598 3746 2602
rect 3710 2558 3714 2562
rect 3790 2598 3794 2602
rect 3814 2598 3818 2602
rect 3774 2578 3778 2582
rect 3806 2588 3810 2592
rect 3694 2548 3698 2552
rect 3718 2548 3722 2552
rect 3686 2538 3690 2542
rect 3670 2528 3674 2532
rect 3550 2458 3554 2462
rect 3630 2458 3634 2462
rect 3582 2448 3586 2452
rect 3598 2448 3602 2452
rect 3542 2368 3546 2372
rect 3526 2328 3530 2332
rect 3526 2308 3530 2312
rect 3542 2338 3546 2342
rect 3558 2438 3562 2442
rect 3582 2408 3586 2412
rect 3582 2348 3586 2352
rect 3542 2298 3546 2302
rect 3566 2298 3570 2302
rect 3574 2298 3578 2302
rect 3574 2278 3578 2282
rect 3550 2258 3554 2262
rect 3566 2228 3570 2232
rect 3534 2208 3538 2212
rect 3574 2208 3578 2212
rect 3478 2158 3482 2162
rect 3510 2158 3514 2162
rect 3422 2148 3426 2152
rect 3494 2148 3498 2152
rect 3414 2138 3418 2142
rect 3446 2138 3450 2142
rect 3422 2118 3426 2122
rect 3294 2088 3298 2092
rect 3366 2088 3370 2092
rect 3382 2088 3386 2092
rect 3398 2068 3402 2072
rect 3414 2068 3418 2072
rect 3438 2068 3442 2072
rect 3278 2048 3282 2052
rect 3262 1888 3266 1892
rect 3214 1878 3218 1882
rect 3198 1858 3202 1862
rect 3198 1788 3202 1792
rect 3134 1748 3138 1752
rect 3166 1748 3170 1752
rect 3222 1748 3226 1752
rect 3246 1858 3250 1862
rect 3270 1788 3274 1792
rect 3270 1758 3274 1762
rect 3238 1738 3242 1742
rect 3270 1738 3274 1742
rect 3206 1728 3210 1732
rect 3230 1728 3234 1732
rect 3142 1708 3146 1712
rect 3126 1678 3130 1682
rect 3118 1668 3122 1672
rect 3134 1618 3138 1622
rect 3118 1578 3122 1582
rect 3126 1578 3130 1582
rect 3046 1548 3050 1552
rect 3014 1538 3018 1542
rect 3030 1538 3034 1542
rect 3070 1538 3074 1542
rect 2950 1518 2954 1522
rect 2958 1508 2962 1512
rect 2934 1498 2938 1502
rect 2974 1488 2978 1492
rect 2934 1468 2938 1472
rect 2958 1458 2962 1462
rect 2974 1458 2978 1462
rect 2982 1448 2986 1452
rect 2966 1438 2970 1442
rect 2894 1418 2898 1422
rect 2910 1418 2914 1422
rect 2822 1368 2826 1372
rect 2870 1358 2874 1362
rect 2886 1358 2890 1362
rect 2838 1348 2842 1352
rect 2854 1348 2858 1352
rect 2846 1338 2850 1342
rect 2870 1338 2874 1342
rect 2910 1398 2914 1402
rect 2878 1318 2882 1322
rect 2838 1308 2842 1312
rect 2870 1298 2874 1302
rect 2790 1268 2794 1272
rect 2846 1268 2850 1272
rect 2638 1168 2642 1172
rect 2654 1168 2658 1172
rect 2638 1138 2642 1142
rect 2606 1118 2610 1122
rect 2542 998 2546 1002
rect 2566 1048 2570 1052
rect 2566 1038 2570 1042
rect 2558 1018 2562 1022
rect 2550 978 2554 982
rect 2622 1108 2626 1112
rect 2590 1068 2594 1072
rect 2622 1068 2626 1072
rect 2614 1048 2618 1052
rect 2630 1048 2634 1052
rect 2586 1003 2590 1007
rect 2593 1003 2597 1007
rect 2566 958 2570 962
rect 2574 958 2578 962
rect 2750 1248 2754 1252
rect 2710 1238 2714 1242
rect 2766 1208 2770 1212
rect 2726 1168 2730 1172
rect 2694 1158 2698 1162
rect 2702 1148 2706 1152
rect 2678 1138 2682 1142
rect 2702 1128 2706 1132
rect 2686 1118 2690 1122
rect 2662 1108 2666 1112
rect 2806 1258 2810 1262
rect 2838 1238 2842 1242
rect 2798 1198 2802 1202
rect 2782 1158 2786 1162
rect 2846 1158 2850 1162
rect 2774 1148 2778 1152
rect 2862 1148 2866 1152
rect 2766 1138 2770 1142
rect 2654 1088 2658 1092
rect 2702 1088 2706 1092
rect 2750 1118 2754 1122
rect 2782 1138 2786 1142
rect 2774 1078 2778 1082
rect 2662 1068 2666 1072
rect 2670 1068 2674 1072
rect 2718 1068 2722 1072
rect 2686 1058 2690 1062
rect 2782 1058 2786 1062
rect 2694 1048 2698 1052
rect 2678 1028 2682 1032
rect 2678 998 2682 1002
rect 2606 948 2610 952
rect 2654 948 2658 952
rect 2510 918 2514 922
rect 2534 918 2538 922
rect 2502 888 2506 892
rect 2526 888 2530 892
rect 2454 848 2458 852
rect 2574 938 2578 942
rect 2582 898 2586 902
rect 2598 868 2602 872
rect 2566 848 2570 852
rect 2558 838 2562 842
rect 2486 808 2490 812
rect 2478 798 2482 802
rect 2374 788 2378 792
rect 2366 758 2370 762
rect 2270 748 2274 752
rect 2294 748 2298 752
rect 2318 748 2322 752
rect 2414 758 2418 762
rect 2238 738 2242 742
rect 2366 738 2370 742
rect 2134 668 2138 672
rect 2182 668 2186 672
rect 2150 648 2154 652
rect 2166 648 2170 652
rect 2222 648 2226 652
rect 2302 728 2306 732
rect 2390 728 2394 732
rect 2318 718 2322 722
rect 2358 718 2362 722
rect 2262 708 2266 712
rect 2286 678 2290 682
rect 2334 698 2338 702
rect 2374 708 2378 712
rect 2374 688 2378 692
rect 2358 678 2362 682
rect 2294 668 2298 672
rect 2350 668 2354 672
rect 2246 588 2250 592
rect 2190 568 2194 572
rect 2214 568 2218 572
rect 2158 558 2162 562
rect 2206 558 2210 562
rect 2174 548 2178 552
rect 2110 538 2114 542
rect 2118 538 2122 542
rect 2142 538 2146 542
rect 2054 528 2058 532
rect 2074 503 2078 507
rect 2081 503 2085 507
rect 2038 498 2042 502
rect 2062 498 2066 502
rect 2102 498 2106 502
rect 2038 488 2042 492
rect 2022 468 2026 472
rect 2006 458 2010 462
rect 2054 468 2058 472
rect 2070 478 2074 482
rect 2086 428 2090 432
rect 1966 388 1970 392
rect 1910 358 1914 362
rect 1870 348 1874 352
rect 1838 338 1842 342
rect 1846 338 1850 342
rect 1830 318 1834 322
rect 1806 288 1810 292
rect 1798 268 1802 272
rect 1822 268 1826 272
rect 1742 248 1746 252
rect 1718 238 1722 242
rect 1686 228 1690 232
rect 1790 258 1794 262
rect 1774 248 1778 252
rect 1806 248 1810 252
rect 1806 238 1810 242
rect 1758 218 1762 222
rect 1790 198 1794 202
rect 1750 188 1754 192
rect 1710 168 1714 172
rect 1646 158 1650 162
rect 1726 158 1730 162
rect 1742 158 1746 162
rect 1758 158 1762 162
rect 1766 158 1770 162
rect 1710 148 1714 152
rect 1758 148 1762 152
rect 1702 138 1706 142
rect 1742 128 1746 132
rect 1582 108 1586 112
rect 1598 88 1602 92
rect 1614 78 1618 82
rect 1766 118 1770 122
rect 1686 88 1690 92
rect 1710 88 1714 92
rect 1542 68 1546 72
rect 1582 68 1586 72
rect 1854 278 1858 282
rect 1870 278 1874 282
rect 1846 228 1850 232
rect 1846 198 1850 202
rect 1870 248 1874 252
rect 1942 328 1946 332
rect 1958 288 1962 292
rect 1926 278 1930 282
rect 1942 268 1946 272
rect 1974 368 1978 372
rect 2054 408 2058 412
rect 2006 398 2010 402
rect 1990 338 1994 342
rect 1982 258 1986 262
rect 1958 248 1962 252
rect 1990 248 1994 252
rect 1910 238 1914 242
rect 1950 228 1954 232
rect 1942 198 1946 202
rect 1886 178 1890 182
rect 1894 178 1898 182
rect 1910 178 1914 182
rect 1862 158 1866 162
rect 1878 158 1882 162
rect 1958 208 1962 212
rect 1910 148 1914 152
rect 1806 138 1810 142
rect 1854 138 1858 142
rect 1902 138 1906 142
rect 1798 128 1802 132
rect 1822 118 1826 122
rect 1774 98 1778 102
rect 1782 98 1786 102
rect 1798 98 1802 102
rect 1814 78 1818 82
rect 1542 58 1546 62
rect 1574 58 1578 62
rect 1638 59 1642 63
rect 1910 78 1914 82
rect 2030 378 2034 382
rect 2054 378 2058 382
rect 2062 358 2066 362
rect 2022 338 2026 342
rect 2038 338 2042 342
rect 2014 328 2018 332
rect 2014 308 2018 312
rect 2022 248 2026 252
rect 2014 218 2018 222
rect 2030 188 2034 192
rect 1974 158 1978 162
rect 1998 108 2002 112
rect 2030 108 2034 112
rect 1990 98 1994 102
rect 1934 68 1938 72
rect 2014 78 2018 82
rect 2022 68 2026 72
rect 1782 58 1786 62
rect 1830 58 1834 62
rect 1894 58 1898 62
rect 2054 208 2058 212
rect 2054 148 2058 152
rect 2038 88 2042 92
rect 2046 78 2050 82
rect 2094 378 2098 382
rect 2074 303 2078 307
rect 2081 303 2085 307
rect 2126 478 2130 482
rect 2118 468 2122 472
rect 2110 418 2114 422
rect 2126 378 2130 382
rect 2586 803 2590 807
rect 2593 803 2597 807
rect 2550 788 2554 792
rect 2542 768 2546 772
rect 2446 748 2450 752
rect 2414 738 2418 742
rect 2430 738 2434 742
rect 2398 718 2402 722
rect 2406 718 2410 722
rect 2382 658 2386 662
rect 2334 648 2338 652
rect 2350 648 2354 652
rect 2366 648 2370 652
rect 2334 598 2338 602
rect 2318 588 2322 592
rect 2310 558 2314 562
rect 2366 558 2370 562
rect 2382 558 2386 562
rect 2262 548 2266 552
rect 2278 548 2282 552
rect 2302 548 2306 552
rect 2326 548 2330 552
rect 2302 538 2306 542
rect 2174 488 2178 492
rect 2150 468 2154 472
rect 2254 478 2258 482
rect 2262 468 2266 472
rect 2262 458 2266 462
rect 2190 398 2194 402
rect 2174 388 2178 392
rect 2158 368 2162 372
rect 2134 338 2138 342
rect 2142 338 2146 342
rect 2174 338 2178 342
rect 2126 328 2130 332
rect 2094 298 2098 302
rect 2070 258 2074 262
rect 2166 318 2170 322
rect 2214 318 2218 322
rect 2134 308 2138 312
rect 2206 298 2210 302
rect 2190 278 2194 282
rect 2182 268 2186 272
rect 2174 258 2178 262
rect 2174 218 2178 222
rect 2102 158 2106 162
rect 2158 158 2162 162
rect 2126 148 2130 152
rect 2142 148 2146 152
rect 2214 288 2218 292
rect 2206 178 2210 182
rect 2310 528 2314 532
rect 2318 518 2322 522
rect 2326 518 2330 522
rect 2310 508 2314 512
rect 2310 448 2314 452
rect 2270 438 2274 442
rect 2238 318 2242 322
rect 2230 288 2234 292
rect 2342 508 2346 512
rect 2334 478 2338 482
rect 2318 398 2322 402
rect 2302 388 2306 392
rect 2278 368 2282 372
rect 2286 368 2290 372
rect 2318 358 2322 362
rect 2326 358 2330 362
rect 2318 328 2322 332
rect 2278 308 2282 312
rect 2270 288 2274 292
rect 2254 258 2258 262
rect 2230 248 2234 252
rect 2262 248 2266 252
rect 2230 238 2234 242
rect 2254 228 2258 232
rect 2238 218 2242 222
rect 2222 158 2226 162
rect 2246 188 2250 192
rect 2214 148 2218 152
rect 2118 138 2122 142
rect 2190 138 2194 142
rect 2198 138 2202 142
rect 2102 108 2106 112
rect 2174 108 2178 112
rect 2074 103 2078 107
rect 2081 103 2085 107
rect 2070 88 2074 92
rect 2382 538 2386 542
rect 2422 628 2426 632
rect 2414 598 2418 602
rect 2398 578 2402 582
rect 2398 528 2402 532
rect 2470 728 2474 732
rect 2478 688 2482 692
rect 2462 678 2466 682
rect 2446 668 2450 672
rect 2454 658 2458 662
rect 2590 728 2594 732
rect 2598 698 2602 702
rect 2566 688 2570 692
rect 2622 938 2626 942
rect 2646 938 2650 942
rect 2630 908 2634 912
rect 2622 888 2626 892
rect 2646 888 2650 892
rect 2646 868 2650 872
rect 2622 858 2626 862
rect 2614 848 2618 852
rect 2614 758 2618 762
rect 2662 848 2666 852
rect 2670 828 2674 832
rect 2638 798 2642 802
rect 2694 888 2698 892
rect 2686 878 2690 882
rect 2694 868 2698 872
rect 2686 848 2690 852
rect 2694 828 2698 832
rect 2662 788 2666 792
rect 2678 788 2682 792
rect 2654 768 2658 772
rect 2622 748 2626 752
rect 2614 738 2618 742
rect 2646 718 2650 722
rect 2630 698 2634 702
rect 2510 668 2514 672
rect 2614 668 2618 672
rect 2454 648 2458 652
rect 2470 648 2474 652
rect 2606 648 2610 652
rect 2622 648 2626 652
rect 2462 628 2466 632
rect 2566 628 2570 632
rect 2598 628 2602 632
rect 2446 598 2450 602
rect 2430 518 2434 522
rect 2478 568 2482 572
rect 2470 548 2474 552
rect 2518 547 2522 551
rect 2494 528 2498 532
rect 2574 618 2578 622
rect 2586 603 2590 607
rect 2593 603 2597 607
rect 2646 678 2650 682
rect 2654 678 2658 682
rect 2750 1028 2754 1032
rect 2766 1028 2770 1032
rect 2838 1138 2842 1142
rect 2806 1128 2810 1132
rect 2862 1088 2866 1092
rect 2830 1078 2834 1082
rect 2862 1068 2866 1072
rect 2854 1058 2858 1062
rect 2838 1048 2842 1052
rect 2798 998 2802 1002
rect 2830 998 2834 1002
rect 3022 1528 3026 1532
rect 2998 1518 3002 1522
rect 3070 1518 3074 1522
rect 3006 1508 3010 1512
rect 3030 1508 3034 1512
rect 3006 1488 3010 1492
rect 3046 1488 3050 1492
rect 3014 1468 3018 1472
rect 3046 1468 3050 1472
rect 3030 1438 3034 1442
rect 2990 1428 2994 1432
rect 2926 1388 2930 1392
rect 2934 1388 2938 1392
rect 2958 1378 2962 1382
rect 2942 1348 2946 1352
rect 2910 1328 2914 1332
rect 2926 1328 2930 1332
rect 2902 1278 2906 1282
rect 2878 1268 2882 1272
rect 2878 1258 2882 1262
rect 2894 1258 2898 1262
rect 2950 1308 2954 1312
rect 3006 1358 3010 1362
rect 2998 1298 3002 1302
rect 2926 1278 2930 1282
rect 2950 1268 2954 1272
rect 2982 1268 2986 1272
rect 2926 1258 2930 1262
rect 2982 1258 2986 1262
rect 2910 1208 2914 1212
rect 2894 1168 2898 1172
rect 2902 1158 2906 1162
rect 2958 1248 2962 1252
rect 2990 1248 2994 1252
rect 2942 1148 2946 1152
rect 2918 1138 2922 1142
rect 2878 1108 2882 1112
rect 2870 968 2874 972
rect 2822 958 2826 962
rect 2798 928 2802 932
rect 2758 838 2762 842
rect 2782 828 2786 832
rect 2710 778 2714 782
rect 2726 758 2730 762
rect 2670 748 2674 752
rect 2710 728 2714 732
rect 2686 688 2690 692
rect 3022 1248 3026 1252
rect 3078 1468 3082 1472
rect 3070 1408 3074 1412
rect 3062 1378 3066 1382
rect 3062 1358 3066 1362
rect 3078 1358 3082 1362
rect 3054 1228 3058 1232
rect 2998 1158 3002 1162
rect 3022 1147 3026 1151
rect 2958 1138 2962 1142
rect 2966 1138 2970 1142
rect 2982 1138 2986 1142
rect 3046 1138 3050 1142
rect 2942 1128 2946 1132
rect 2982 1118 2986 1122
rect 2934 1098 2938 1102
rect 2934 1078 2938 1082
rect 2926 1068 2930 1072
rect 2934 1058 2938 1062
rect 2926 1048 2930 1052
rect 2942 1048 2946 1052
rect 2998 1088 3002 1092
rect 3070 1078 3074 1082
rect 3006 1068 3010 1072
rect 3038 1068 3042 1072
rect 3038 1058 3042 1062
rect 3078 1048 3082 1052
rect 3022 1008 3026 1012
rect 2966 978 2970 982
rect 2926 958 2930 962
rect 2958 958 2962 962
rect 3054 988 3058 992
rect 3022 958 3026 962
rect 2870 948 2874 952
rect 2918 948 2922 952
rect 2854 938 2858 942
rect 2894 938 2898 942
rect 2878 918 2882 922
rect 2854 898 2858 902
rect 2830 878 2834 882
rect 2846 828 2850 832
rect 2894 888 2898 892
rect 2910 878 2914 882
rect 2886 868 2890 872
rect 2894 858 2898 862
rect 2862 808 2866 812
rect 2798 758 2802 762
rect 2894 798 2898 802
rect 2974 928 2978 932
rect 2982 928 2986 932
rect 2950 898 2954 902
rect 2926 878 2930 882
rect 2966 878 2970 882
rect 2958 868 2962 872
rect 3030 948 3034 952
rect 3078 948 3082 952
rect 3014 938 3018 942
rect 3014 918 3018 922
rect 2918 848 2922 852
rect 2902 748 2906 752
rect 2806 738 2810 742
rect 2790 728 2794 732
rect 2822 678 2826 682
rect 2646 658 2650 662
rect 2614 628 2618 632
rect 2630 618 2634 622
rect 2638 558 2642 562
rect 2502 508 2506 512
rect 2566 508 2570 512
rect 2462 498 2466 502
rect 2510 478 2514 482
rect 2382 468 2386 472
rect 2406 468 2410 472
rect 2430 468 2434 472
rect 2494 468 2498 472
rect 2542 468 2546 472
rect 2350 448 2354 452
rect 2430 458 2434 462
rect 2374 438 2378 442
rect 2382 438 2386 442
rect 2342 418 2346 422
rect 2350 408 2354 412
rect 2366 388 2370 392
rect 2414 438 2418 442
rect 2406 418 2410 422
rect 2374 368 2378 372
rect 2358 338 2362 342
rect 2390 368 2394 372
rect 2334 318 2338 322
rect 2342 318 2346 322
rect 2374 318 2378 322
rect 2398 318 2402 322
rect 2326 308 2330 312
rect 2374 308 2378 312
rect 2382 308 2386 312
rect 2286 298 2290 302
rect 2318 298 2322 302
rect 2286 288 2290 292
rect 2302 278 2306 282
rect 2390 288 2394 292
rect 2382 268 2386 272
rect 2446 448 2450 452
rect 2438 428 2442 432
rect 2438 398 2442 402
rect 2414 368 2418 372
rect 2406 288 2410 292
rect 2414 288 2418 292
rect 2454 388 2458 392
rect 2446 288 2450 292
rect 2486 458 2490 462
rect 2550 448 2554 452
rect 2494 438 2498 442
rect 2470 408 2474 412
rect 2510 368 2514 372
rect 2446 278 2450 282
rect 2462 278 2466 282
rect 2586 403 2590 407
rect 2593 403 2597 407
rect 2678 648 2682 652
rect 2798 658 2802 662
rect 2790 648 2794 652
rect 2718 628 2722 632
rect 2670 618 2674 622
rect 2694 558 2698 562
rect 2750 548 2754 552
rect 2798 548 2802 552
rect 2742 538 2746 542
rect 2774 538 2778 542
rect 2678 528 2682 532
rect 2758 528 2762 532
rect 2662 488 2666 492
rect 2654 478 2658 482
rect 2670 468 2674 472
rect 2726 518 2730 522
rect 2614 458 2618 462
rect 2630 458 2634 462
rect 2678 458 2682 462
rect 2726 458 2730 462
rect 2694 448 2698 452
rect 2662 438 2666 442
rect 2654 398 2658 402
rect 2622 388 2626 392
rect 2606 368 2610 372
rect 2558 358 2562 362
rect 2742 408 2746 412
rect 2734 388 2738 392
rect 2694 368 2698 372
rect 2710 358 2714 362
rect 2654 348 2658 352
rect 2686 348 2690 352
rect 2710 348 2714 352
rect 2686 328 2690 332
rect 2686 308 2690 312
rect 2638 288 2642 292
rect 2646 288 2650 292
rect 2438 258 2442 262
rect 2438 238 2442 242
rect 2286 218 2290 222
rect 2782 478 2786 482
rect 2846 698 2850 702
rect 2854 678 2858 682
rect 2838 588 2842 592
rect 2870 588 2874 592
rect 2838 558 2842 562
rect 2830 518 2834 522
rect 2910 668 2914 672
rect 2886 648 2890 652
rect 2902 648 2906 652
rect 2886 608 2890 612
rect 2982 838 2986 842
rect 2958 828 2962 832
rect 2942 778 2946 782
rect 2926 768 2930 772
rect 2966 788 2970 792
rect 2942 698 2946 702
rect 2934 678 2938 682
rect 2934 658 2938 662
rect 2934 648 2938 652
rect 2950 648 2954 652
rect 2974 758 2978 762
rect 3038 848 3042 852
rect 3014 828 3018 832
rect 3098 1503 3102 1507
rect 3105 1503 3109 1507
rect 3182 1718 3186 1722
rect 3190 1718 3194 1722
rect 3222 1718 3226 1722
rect 3174 1698 3178 1702
rect 3158 1688 3162 1692
rect 3166 1688 3170 1692
rect 3222 1648 3226 1652
rect 3270 1718 3274 1722
rect 3182 1608 3186 1612
rect 3214 1608 3218 1612
rect 3166 1578 3170 1582
rect 3174 1578 3178 1582
rect 3206 1598 3210 1602
rect 3206 1558 3210 1562
rect 3158 1548 3162 1552
rect 3334 2058 3338 2062
rect 3310 1947 3314 1951
rect 3446 2058 3450 2062
rect 3350 2038 3354 2042
rect 3414 2038 3418 2042
rect 3446 2038 3450 2042
rect 3430 2028 3434 2032
rect 3462 2108 3466 2112
rect 3502 2108 3506 2112
rect 3486 2068 3490 2072
rect 3550 2128 3554 2132
rect 3574 2128 3578 2132
rect 3526 2108 3530 2112
rect 3558 2118 3562 2122
rect 3550 2088 3554 2092
rect 3478 2058 3482 2062
rect 3518 2058 3522 2062
rect 3462 2048 3466 2052
rect 3502 2048 3506 2052
rect 3494 2028 3498 2032
rect 3478 2008 3482 2012
rect 3358 1958 3362 1962
rect 3454 1958 3458 1962
rect 3486 1978 3490 1982
rect 3358 1948 3362 1952
rect 3366 1948 3370 1952
rect 3374 1948 3378 1952
rect 3406 1948 3410 1952
rect 3422 1948 3426 1952
rect 3430 1948 3434 1952
rect 3382 1938 3386 1942
rect 3462 1938 3466 1942
rect 3358 1928 3362 1932
rect 3390 1928 3394 1932
rect 3334 1908 3338 1912
rect 3358 1908 3362 1912
rect 3310 1728 3314 1732
rect 3286 1698 3290 1702
rect 3438 1898 3442 1902
rect 3326 1848 3330 1852
rect 3334 1848 3338 1852
rect 3342 1758 3346 1762
rect 3390 1858 3394 1862
rect 3486 1928 3490 1932
rect 3478 1908 3482 1912
rect 3470 1848 3474 1852
rect 3510 1958 3514 1962
rect 3542 2048 3546 2052
rect 3502 1938 3506 1942
rect 3494 1868 3498 1872
rect 3502 1848 3506 1852
rect 3406 1788 3410 1792
rect 3382 1778 3386 1782
rect 3374 1748 3378 1752
rect 3398 1758 3402 1762
rect 3662 2498 3666 2502
rect 3638 2438 3642 2442
rect 3654 2438 3658 2442
rect 3662 2418 3666 2422
rect 3610 2403 3614 2407
rect 3617 2403 3621 2407
rect 3638 2358 3642 2362
rect 3630 2348 3634 2352
rect 3606 2328 3610 2332
rect 3622 2308 3626 2312
rect 3646 2328 3650 2332
rect 3630 2298 3634 2302
rect 3742 2538 3746 2542
rect 3774 2538 3778 2542
rect 3742 2498 3746 2502
rect 3702 2458 3706 2462
rect 3726 2448 3730 2452
rect 3734 2448 3738 2452
rect 3678 2368 3682 2372
rect 3702 2308 3706 2312
rect 3678 2298 3682 2302
rect 3630 2278 3634 2282
rect 3590 2258 3594 2262
rect 3638 2258 3642 2262
rect 3610 2203 3614 2207
rect 3617 2203 3621 2207
rect 3630 2168 3634 2172
rect 3590 2158 3594 2162
rect 3606 2148 3610 2152
rect 3646 2248 3650 2252
rect 3702 2238 3706 2242
rect 3654 2188 3658 2192
rect 3670 2188 3674 2192
rect 3646 2158 3650 2162
rect 3678 2148 3682 2152
rect 3686 2148 3690 2152
rect 3622 2138 3626 2142
rect 3638 2138 3642 2142
rect 3646 2128 3650 2132
rect 3742 2388 3746 2392
rect 3742 2378 3746 2382
rect 4006 3138 4010 3142
rect 4014 3068 4018 3072
rect 4038 3178 4042 3182
rect 4030 3078 4034 3082
rect 4046 3158 4050 3162
rect 4054 3128 4058 3132
rect 4094 3128 4098 3132
rect 4054 3068 4058 3072
rect 4030 3058 4034 3062
rect 4086 3058 4090 3062
rect 3958 2948 3962 2952
rect 3950 2918 3954 2922
rect 4054 3008 4058 3012
rect 4022 2978 4026 2982
rect 4086 2978 4090 2982
rect 4038 2948 4042 2952
rect 4062 2948 4066 2952
rect 3966 2908 3970 2912
rect 4006 2908 4010 2912
rect 4022 2908 4026 2912
rect 3958 2878 3962 2882
rect 3958 2868 3962 2872
rect 3942 2848 3946 2852
rect 3934 2838 3938 2842
rect 3934 2748 3938 2752
rect 3950 2748 3954 2752
rect 4254 3438 4258 3442
rect 4262 3378 4266 3382
rect 4246 3348 4250 3352
rect 4254 3348 4258 3352
rect 4222 3338 4226 3342
rect 4262 3338 4266 3342
rect 4246 3328 4250 3332
rect 4198 3318 4202 3322
rect 4214 3288 4218 3292
rect 4246 3298 4250 3302
rect 4206 3278 4210 3282
rect 4142 3268 4146 3272
rect 4174 3268 4178 3272
rect 4214 3268 4218 3272
rect 4238 3268 4242 3272
rect 4158 3258 4162 3262
rect 4206 3248 4210 3252
rect 4214 3238 4218 3242
rect 4246 3248 4250 3252
rect 4286 3308 4290 3312
rect 4334 3718 4338 3722
rect 4382 3808 4386 3812
rect 4366 3758 4370 3762
rect 4462 3848 4466 3852
rect 4502 3848 4506 3852
rect 4446 3808 4450 3812
rect 4406 3748 4410 3752
rect 4390 3728 4394 3732
rect 4398 3718 4402 3722
rect 4342 3698 4346 3702
rect 4382 3698 4386 3702
rect 4358 3678 4362 3682
rect 4302 3558 4306 3562
rect 4318 3648 4322 3652
rect 4374 3648 4378 3652
rect 4358 3628 4362 3632
rect 4366 3608 4370 3612
rect 4342 3548 4346 3552
rect 4358 3548 4362 3552
rect 4358 3468 4362 3472
rect 4318 3428 4322 3432
rect 4310 3418 4314 3422
rect 4302 3328 4306 3332
rect 4230 3218 4234 3222
rect 4254 3218 4258 3222
rect 4174 3198 4178 3202
rect 4190 3198 4194 3202
rect 4158 3178 4162 3182
rect 4198 3168 4202 3172
rect 4206 3158 4210 3162
rect 4246 3158 4250 3162
rect 4134 3128 4138 3132
rect 4114 3103 4118 3107
rect 4121 3103 4125 3107
rect 4110 3048 4114 3052
rect 4302 3208 4306 3212
rect 4358 3388 4362 3392
rect 4350 3368 4354 3372
rect 4470 3788 4474 3792
rect 4422 3718 4426 3722
rect 4406 3638 4410 3642
rect 4390 3588 4394 3592
rect 4422 3578 4426 3582
rect 4382 3568 4386 3572
rect 4422 3568 4426 3572
rect 4438 3708 4442 3712
rect 4446 3658 4450 3662
rect 4470 3658 4474 3662
rect 4486 3658 4490 3662
rect 4454 3648 4458 3652
rect 4494 3638 4498 3642
rect 4446 3568 4450 3572
rect 4510 3568 4514 3572
rect 4390 3548 4394 3552
rect 4390 3528 4394 3532
rect 4398 3518 4402 3522
rect 4366 3338 4370 3342
rect 4422 3488 4426 3492
rect 4438 3478 4442 3482
rect 4470 3558 4474 3562
rect 4582 3968 4586 3972
rect 4598 3968 4602 3972
rect 4542 3948 4546 3952
rect 4558 3948 4562 3952
rect 4590 3938 4594 3942
rect 4526 3928 4530 3932
rect 4590 3918 4594 3922
rect 4534 3898 4538 3902
rect 4542 3898 4546 3902
rect 4550 3878 4554 3882
rect 4598 3878 4602 3882
rect 4614 4048 4618 4052
rect 4654 4048 4658 4052
rect 4634 4003 4638 4007
rect 4641 4003 4645 4007
rect 4622 3948 4626 3952
rect 4638 3938 4642 3942
rect 4614 3928 4618 3932
rect 4622 3918 4626 3922
rect 4582 3868 4586 3872
rect 4542 3848 4546 3852
rect 4582 3818 4586 3822
rect 4574 3748 4578 3752
rect 4558 3738 4562 3742
rect 4590 3758 4594 3762
rect 4598 3738 4602 3742
rect 4606 3728 4610 3732
rect 4654 3908 4658 3912
rect 4710 4178 4714 4182
rect 4678 4158 4682 4162
rect 4694 4148 4698 4152
rect 4718 4138 4722 4142
rect 4702 4088 4706 4092
rect 4718 4038 4722 4042
rect 4678 3978 4682 3982
rect 4702 3958 4706 3962
rect 4686 3948 4690 3952
rect 4678 3938 4682 3942
rect 4702 3938 4706 3942
rect 4662 3898 4666 3902
rect 4630 3868 4634 3872
rect 4662 3868 4666 3872
rect 4702 3888 4706 3892
rect 4878 4228 4882 4232
rect 4870 4188 4874 4192
rect 4886 4188 4890 4192
rect 4766 4148 4770 4152
rect 4798 4148 4802 4152
rect 4822 4148 4826 4152
rect 4750 4128 4754 4132
rect 4742 4098 4746 4102
rect 4918 4338 4922 4342
rect 4918 4308 4922 4312
rect 4918 4278 4922 4282
rect 4902 4268 4906 4272
rect 4894 4158 4898 4162
rect 4870 4138 4874 4142
rect 4814 4108 4818 4112
rect 4734 4078 4738 4082
rect 4766 4068 4770 4072
rect 4790 4068 4794 4072
rect 4774 4058 4778 4062
rect 4734 3978 4738 3982
rect 4750 3978 4754 3982
rect 4758 3968 4762 3972
rect 4734 3958 4738 3962
rect 4766 3948 4770 3952
rect 4782 3948 4786 3952
rect 4878 4098 4882 4102
rect 4958 4288 4962 4292
rect 4974 4358 4978 4362
rect 5046 4458 5050 4462
rect 5038 4438 5042 4442
rect 5054 4438 5058 4442
rect 5014 4378 5018 4382
rect 5078 4368 5082 4372
rect 5110 4448 5114 4452
rect 5190 4508 5194 4512
rect 5174 4498 5178 4502
rect 5174 4478 5178 4482
rect 5022 4358 5026 4362
rect 5046 4358 5050 4362
rect 5030 4348 5034 4352
rect 5070 4338 5074 4342
rect 5118 4338 5122 4342
rect 5030 4328 5034 4332
rect 5014 4318 5018 4322
rect 5086 4318 5090 4322
rect 5182 4358 5186 4362
rect 5126 4268 5130 4272
rect 5150 4268 5154 4272
rect 4998 4258 5002 4262
rect 4974 4248 4978 4252
rect 5006 4228 5010 4232
rect 4942 4158 4946 4162
rect 5006 4158 5010 4162
rect 4950 4148 4954 4152
rect 4910 4128 4914 4132
rect 4870 4088 4874 4092
rect 4886 4088 4890 4092
rect 4854 4058 4858 4062
rect 4886 4078 4890 4082
rect 4926 4018 4930 4022
rect 4870 3978 4874 3982
rect 4822 3958 4826 3962
rect 4830 3948 4834 3952
rect 4766 3928 4770 3932
rect 4814 3878 4818 3882
rect 4766 3868 4770 3872
rect 4830 3868 4834 3872
rect 4854 3868 4858 3872
rect 4878 3958 4882 3962
rect 4886 3948 4890 3952
rect 4878 3888 4882 3892
rect 4926 3978 4930 3982
rect 4918 3958 4922 3962
rect 4918 3928 4922 3932
rect 4902 3918 4906 3922
rect 4910 3918 4914 3922
rect 4950 4128 4954 4132
rect 4982 4058 4986 4062
rect 4998 4058 5002 4062
rect 4958 4018 4962 4022
rect 4942 3948 4946 3952
rect 4934 3888 4938 3892
rect 4950 3888 4954 3892
rect 4990 3888 4994 3892
rect 4934 3868 4938 3872
rect 4758 3858 4762 3862
rect 4822 3858 4826 3862
rect 4886 3858 4890 3862
rect 4894 3858 4898 3862
rect 4634 3803 4638 3807
rect 4641 3803 4645 3807
rect 4806 3848 4810 3852
rect 4870 3848 4874 3852
rect 4750 3838 4754 3842
rect 4726 3828 4730 3832
rect 4694 3788 4698 3792
rect 4710 3778 4714 3782
rect 4766 3778 4770 3782
rect 4710 3758 4714 3762
rect 4734 3758 4738 3762
rect 4710 3748 4714 3752
rect 4726 3748 4730 3752
rect 4646 3738 4650 3742
rect 4686 3728 4690 3732
rect 4606 3678 4610 3682
rect 4582 3648 4586 3652
rect 4542 3568 4546 3572
rect 4582 3568 4586 3572
rect 4494 3548 4498 3552
rect 4518 3548 4522 3552
rect 4534 3548 4538 3552
rect 4510 3538 4514 3542
rect 4518 3538 4522 3542
rect 4470 3488 4474 3492
rect 4462 3468 4466 3472
rect 4430 3458 4434 3462
rect 4470 3458 4474 3462
rect 4406 3448 4410 3452
rect 4446 3448 4450 3452
rect 4390 3398 4394 3402
rect 4438 3408 4442 3412
rect 4430 3368 4434 3372
rect 4398 3358 4402 3362
rect 4406 3358 4410 3362
rect 4502 3358 4506 3362
rect 4382 3348 4386 3352
rect 4438 3348 4442 3352
rect 4534 3528 4538 3532
rect 4526 3518 4530 3522
rect 4542 3518 4546 3522
rect 4574 3538 4578 3542
rect 4566 3518 4570 3522
rect 4382 3328 4386 3332
rect 4398 3328 4402 3332
rect 4366 3318 4370 3322
rect 4310 3178 4314 3182
rect 4262 3138 4266 3142
rect 4166 3108 4170 3112
rect 4214 3108 4218 3112
rect 4214 3098 4218 3102
rect 4230 3098 4234 3102
rect 4222 3078 4226 3082
rect 4294 3138 4298 3142
rect 4286 3128 4290 3132
rect 4270 3088 4274 3092
rect 4286 3088 4290 3092
rect 4238 3058 4242 3062
rect 4246 3058 4250 3062
rect 4238 3038 4242 3042
rect 4238 3018 4242 3022
rect 4190 2968 4194 2972
rect 4102 2958 4106 2962
rect 4142 2948 4146 2952
rect 4118 2938 4122 2942
rect 4086 2928 4090 2932
rect 4118 2928 4122 2932
rect 4078 2898 4082 2902
rect 4038 2888 4042 2892
rect 4134 2908 4138 2912
rect 4114 2903 4118 2907
rect 4121 2903 4125 2907
rect 4006 2858 4010 2862
rect 4054 2858 4058 2862
rect 4102 2858 4106 2862
rect 4142 2898 4146 2902
rect 4174 2938 4178 2942
rect 4166 2928 4170 2932
rect 4150 2888 4154 2892
rect 4182 2898 4186 2902
rect 4206 2928 4210 2932
rect 4158 2878 4162 2882
rect 4166 2878 4170 2882
rect 4150 2858 4154 2862
rect 4022 2848 4026 2852
rect 3998 2818 4002 2822
rect 3974 2798 3978 2802
rect 3998 2758 4002 2762
rect 3974 2748 3978 2752
rect 4014 2748 4018 2752
rect 3958 2738 3962 2742
rect 3982 2738 3986 2742
rect 3950 2728 3954 2732
rect 3910 2718 3914 2722
rect 3926 2718 3930 2722
rect 3910 2698 3914 2702
rect 3926 2698 3930 2702
rect 3998 2698 4002 2702
rect 3910 2688 3914 2692
rect 3942 2688 3946 2692
rect 3934 2678 3938 2682
rect 4038 2838 4042 2842
rect 4214 2908 4218 2912
rect 4246 2908 4250 2912
rect 4222 2898 4226 2902
rect 4446 3308 4450 3312
rect 4622 3658 4626 3662
rect 4750 3738 4754 3742
rect 4846 3838 4850 3842
rect 4878 3838 4882 3842
rect 4878 3788 4882 3792
rect 4734 3728 4738 3732
rect 4694 3718 4698 3722
rect 4662 3688 4666 3692
rect 4606 3598 4610 3602
rect 4598 3588 4602 3592
rect 4598 3578 4602 3582
rect 4638 3628 4642 3632
rect 4686 3698 4690 3702
rect 4710 3688 4714 3692
rect 4678 3678 4682 3682
rect 4710 3658 4714 3662
rect 4694 3648 4698 3652
rect 4734 3698 4738 3702
rect 4686 3638 4690 3642
rect 4702 3638 4706 3642
rect 4726 3638 4730 3642
rect 4726 3628 4730 3632
rect 4670 3618 4674 3622
rect 4654 3608 4658 3612
rect 4634 3603 4638 3607
rect 4641 3603 4645 3607
rect 4702 3598 4706 3602
rect 4614 3558 4618 3562
rect 4622 3558 4626 3562
rect 4630 3558 4634 3562
rect 4670 3558 4674 3562
rect 4710 3568 4714 3572
rect 4726 3568 4730 3572
rect 4598 3518 4602 3522
rect 4606 3518 4610 3522
rect 4590 3498 4594 3502
rect 4606 3488 4610 3492
rect 4622 3428 4626 3432
rect 4614 3388 4618 3392
rect 4558 3368 4562 3372
rect 4566 3358 4570 3362
rect 4598 3348 4602 3352
rect 4566 3328 4570 3332
rect 4398 3298 4402 3302
rect 4438 3298 4442 3302
rect 4486 3298 4490 3302
rect 4542 3298 4546 3302
rect 4454 3288 4458 3292
rect 4398 3278 4402 3282
rect 4382 3268 4386 3272
rect 4414 3258 4418 3262
rect 4430 3258 4434 3262
rect 4438 3258 4442 3262
rect 4470 3228 4474 3232
rect 4446 3218 4450 3222
rect 4318 3068 4322 3072
rect 4334 3068 4338 3072
rect 4310 3058 4314 3062
rect 4342 3058 4346 3062
rect 4350 3058 4354 3062
rect 4278 3048 4282 3052
rect 4302 3048 4306 3052
rect 4318 3038 4322 3042
rect 4270 3028 4274 3032
rect 4278 3018 4282 3022
rect 4326 2998 4330 3002
rect 4294 2978 4298 2982
rect 4342 2978 4346 2982
rect 4310 2958 4314 2962
rect 4334 2948 4338 2952
rect 4326 2938 4330 2942
rect 4342 2938 4346 2942
rect 4262 2928 4266 2932
rect 4254 2888 4258 2892
rect 4286 2888 4290 2892
rect 4294 2888 4298 2892
rect 4310 2888 4314 2892
rect 4230 2878 4234 2882
rect 4262 2868 4266 2872
rect 4286 2868 4290 2872
rect 4206 2858 4210 2862
rect 4254 2858 4258 2862
rect 4094 2848 4098 2852
rect 4166 2848 4170 2852
rect 4086 2798 4090 2802
rect 4166 2798 4170 2802
rect 4070 2748 4074 2752
rect 4118 2748 4122 2752
rect 4142 2748 4146 2752
rect 4062 2738 4066 2742
rect 4022 2728 4026 2732
rect 4030 2728 4034 2732
rect 4070 2728 4074 2732
rect 4006 2688 4010 2692
rect 4078 2708 4082 2712
rect 4062 2678 4066 2682
rect 3934 2658 3938 2662
rect 4006 2658 4010 2662
rect 3902 2648 3906 2652
rect 3950 2628 3954 2632
rect 3862 2578 3866 2582
rect 3918 2578 3922 2582
rect 3814 2548 3818 2552
rect 3838 2538 3842 2542
rect 3830 2528 3834 2532
rect 3902 2548 3906 2552
rect 3974 2608 3978 2612
rect 4054 2648 4058 2652
rect 4046 2608 4050 2612
rect 4038 2598 4042 2602
rect 4014 2578 4018 2582
rect 4022 2578 4026 2582
rect 3950 2568 3954 2572
rect 3918 2508 3922 2512
rect 3766 2488 3770 2492
rect 3798 2488 3802 2492
rect 3758 2458 3762 2462
rect 3782 2458 3786 2462
rect 3766 2448 3770 2452
rect 3782 2408 3786 2412
rect 3846 2468 3850 2472
rect 3854 2468 3858 2472
rect 3910 2468 3914 2472
rect 3934 2468 3938 2472
rect 3814 2448 3818 2452
rect 3822 2438 3826 2442
rect 3886 2418 3890 2422
rect 3846 2398 3850 2402
rect 3758 2388 3762 2392
rect 3790 2388 3794 2392
rect 3798 2388 3802 2392
rect 3750 2358 3754 2362
rect 3782 2368 3786 2372
rect 3878 2378 3882 2382
rect 3902 2448 3906 2452
rect 3910 2448 3914 2452
rect 3926 2448 3930 2452
rect 3934 2438 3938 2442
rect 4022 2528 4026 2532
rect 4070 2608 4074 2612
rect 4062 2598 4066 2602
rect 4006 2508 4010 2512
rect 4054 2508 4058 2512
rect 3958 2498 3962 2502
rect 3974 2468 3978 2472
rect 3990 2468 3994 2472
rect 3958 2448 3962 2452
rect 3870 2368 3874 2372
rect 3894 2368 3898 2372
rect 3814 2358 3818 2362
rect 3910 2358 3914 2362
rect 3846 2348 3850 2352
rect 3862 2348 3866 2352
rect 3822 2338 3826 2342
rect 3766 2328 3770 2332
rect 3838 2328 3842 2332
rect 3910 2308 3914 2312
rect 3814 2298 3818 2302
rect 3878 2298 3882 2302
rect 3902 2298 3906 2302
rect 3782 2288 3786 2292
rect 3798 2288 3802 2292
rect 3806 2288 3810 2292
rect 3830 2288 3834 2292
rect 3862 2288 3866 2292
rect 3886 2288 3890 2292
rect 3742 2258 3746 2262
rect 3838 2258 3842 2262
rect 3926 2278 3930 2282
rect 3758 2248 3762 2252
rect 3806 2248 3810 2252
rect 3846 2248 3850 2252
rect 3918 2248 3922 2252
rect 3726 2238 3730 2242
rect 3766 2238 3770 2242
rect 3822 2238 3826 2242
rect 3862 2238 3866 2242
rect 3894 2238 3898 2242
rect 3870 2228 3874 2232
rect 3878 2228 3882 2232
rect 3766 2218 3770 2222
rect 3726 2178 3730 2182
rect 3734 2178 3738 2182
rect 3742 2178 3746 2182
rect 3702 2108 3706 2112
rect 3686 2078 3690 2082
rect 3670 2068 3674 2072
rect 3654 2058 3658 2062
rect 3582 2048 3586 2052
rect 3646 2048 3650 2052
rect 3558 2018 3562 2022
rect 3610 2003 3614 2007
rect 3617 2003 3621 2007
rect 3582 1998 3586 2002
rect 3654 2008 3658 2012
rect 3774 2198 3778 2202
rect 3838 2188 3842 2192
rect 3806 2168 3810 2172
rect 3766 2158 3770 2162
rect 3782 2158 3786 2162
rect 3750 2148 3754 2152
rect 3790 2148 3794 2152
rect 3830 2158 3834 2162
rect 3734 2138 3738 2142
rect 3758 2138 3762 2142
rect 3774 2128 3778 2132
rect 3862 2148 3866 2152
rect 3862 2138 3866 2142
rect 3854 2128 3858 2132
rect 3822 2118 3826 2122
rect 3814 2108 3818 2112
rect 3782 2078 3786 2082
rect 3718 2068 3722 2072
rect 3846 2068 3850 2072
rect 3726 2058 3730 2062
rect 3798 2018 3802 2022
rect 3806 2018 3810 2022
rect 3590 1978 3594 1982
rect 3710 1978 3714 1982
rect 3790 1978 3794 1982
rect 3622 1958 3626 1962
rect 3718 1958 3722 1962
rect 3766 1958 3770 1962
rect 3790 1958 3794 1962
rect 3574 1938 3578 1942
rect 3590 1938 3594 1942
rect 3534 1928 3538 1932
rect 3542 1928 3546 1932
rect 3558 1928 3562 1932
rect 3574 1908 3578 1912
rect 3542 1898 3546 1902
rect 3846 1988 3850 1992
rect 3822 1958 3826 1962
rect 3870 2078 3874 2082
rect 3862 2068 3866 2072
rect 3902 2158 3906 2162
rect 3918 2158 3922 2162
rect 3894 2148 3898 2152
rect 3886 2108 3890 2112
rect 3910 2098 3914 2102
rect 3902 2078 3906 2082
rect 3998 2438 4002 2442
rect 3982 2418 3986 2422
rect 3966 2408 3970 2412
rect 3998 2358 4002 2362
rect 4030 2468 4034 2472
rect 4114 2703 4118 2707
rect 4121 2703 4125 2707
rect 4134 2698 4138 2702
rect 4086 2678 4090 2682
rect 4158 2708 4162 2712
rect 4142 2668 4146 2672
rect 4142 2658 4146 2662
rect 4214 2828 4218 2832
rect 4198 2818 4202 2822
rect 4182 2808 4186 2812
rect 4174 2758 4178 2762
rect 4206 2798 4210 2802
rect 4230 2798 4234 2802
rect 4246 2798 4250 2802
rect 4190 2658 4194 2662
rect 4206 2658 4210 2662
rect 4094 2618 4098 2622
rect 4158 2618 4162 2622
rect 4094 2588 4098 2592
rect 4110 2568 4114 2572
rect 4158 2558 4162 2562
rect 4166 2558 4170 2562
rect 4134 2548 4138 2552
rect 4102 2538 4106 2542
rect 4142 2538 4146 2542
rect 4086 2528 4090 2532
rect 4114 2503 4118 2507
rect 4121 2503 4125 2507
rect 4078 2498 4082 2502
rect 4134 2498 4138 2502
rect 4102 2488 4106 2492
rect 4094 2468 4098 2472
rect 4014 2458 4018 2462
rect 4046 2458 4050 2462
rect 4110 2458 4114 2462
rect 4038 2438 4042 2442
rect 4030 2418 4034 2422
rect 4014 2378 4018 2382
rect 4030 2358 4034 2362
rect 4022 2348 4026 2352
rect 3982 2338 3986 2342
rect 4022 2328 4026 2332
rect 3974 2308 3978 2312
rect 3998 2298 4002 2302
rect 3974 2248 3978 2252
rect 3974 2158 3978 2162
rect 4062 2448 4066 2452
rect 4086 2448 4090 2452
rect 4094 2448 4098 2452
rect 4070 2408 4074 2412
rect 4038 2348 4042 2352
rect 4054 2348 4058 2352
rect 4118 2408 4122 2412
rect 4174 2508 4178 2512
rect 4166 2478 4170 2482
rect 4158 2448 4162 2452
rect 4150 2438 4154 2442
rect 4158 2418 4162 2422
rect 4126 2348 4130 2352
rect 4054 2338 4058 2342
rect 4046 2328 4050 2332
rect 4078 2328 4082 2332
rect 4078 2298 4082 2302
rect 4030 2258 4034 2262
rect 4046 2248 4050 2252
rect 4070 2248 4074 2252
rect 4062 2238 4066 2242
rect 4022 2188 4026 2192
rect 4114 2303 4118 2307
rect 4121 2303 4125 2307
rect 4134 2208 4138 2212
rect 4078 2188 4082 2192
rect 4054 2168 4058 2172
rect 4110 2158 4114 2162
rect 4030 2148 4034 2152
rect 4038 2138 4042 2142
rect 3958 2118 3962 2122
rect 3966 2098 3970 2102
rect 3926 2068 3930 2072
rect 3942 2068 3946 2072
rect 4014 2128 4018 2132
rect 4046 2128 4050 2132
rect 4006 2118 4010 2122
rect 3910 2058 3914 2062
rect 3934 2058 3938 2062
rect 3654 1948 3658 1952
rect 3758 1948 3762 1952
rect 3670 1938 3674 1942
rect 3678 1928 3682 1932
rect 3758 1928 3762 1932
rect 3798 1928 3802 1932
rect 3630 1908 3634 1912
rect 3534 1878 3538 1882
rect 3550 1878 3554 1882
rect 3598 1878 3602 1882
rect 3638 1878 3642 1882
rect 3550 1868 3554 1872
rect 3558 1868 3562 1872
rect 3574 1868 3578 1872
rect 3590 1868 3594 1872
rect 3582 1828 3586 1832
rect 3590 1828 3594 1832
rect 3558 1798 3562 1802
rect 3422 1778 3426 1782
rect 3518 1778 3522 1782
rect 3574 1778 3578 1782
rect 3398 1728 3402 1732
rect 3390 1718 3394 1722
rect 3526 1758 3530 1762
rect 3558 1758 3562 1762
rect 3454 1748 3458 1752
rect 3502 1748 3506 1752
rect 3510 1748 3514 1752
rect 3430 1728 3434 1732
rect 3422 1718 3426 1722
rect 3414 1688 3418 1692
rect 3326 1668 3330 1672
rect 3382 1668 3386 1672
rect 3302 1648 3306 1652
rect 3270 1638 3274 1642
rect 3310 1638 3314 1642
rect 3254 1558 3258 1562
rect 3158 1538 3162 1542
rect 3190 1538 3194 1542
rect 3246 1538 3250 1542
rect 3142 1508 3146 1512
rect 3118 1498 3122 1502
rect 3190 1508 3194 1512
rect 3310 1598 3314 1602
rect 3382 1598 3386 1602
rect 3326 1578 3330 1582
rect 3342 1578 3346 1582
rect 3454 1728 3458 1732
rect 3518 1708 3522 1712
rect 3526 1708 3530 1712
rect 3486 1688 3490 1692
rect 3446 1658 3450 1662
rect 3438 1648 3442 1652
rect 3414 1608 3418 1612
rect 3406 1588 3410 1592
rect 3406 1578 3410 1582
rect 3366 1558 3370 1562
rect 3318 1548 3322 1552
rect 3366 1548 3370 1552
rect 3310 1528 3314 1532
rect 3342 1528 3346 1532
rect 3350 1528 3354 1532
rect 3278 1518 3282 1522
rect 3094 1488 3098 1492
rect 3102 1488 3106 1492
rect 3158 1488 3162 1492
rect 3198 1488 3202 1492
rect 3222 1488 3226 1492
rect 3270 1488 3274 1492
rect 3126 1468 3130 1472
rect 3158 1468 3162 1472
rect 3182 1468 3186 1472
rect 3118 1418 3122 1422
rect 3110 1408 3114 1412
rect 3094 1398 3098 1402
rect 3094 1358 3098 1362
rect 3110 1328 3114 1332
rect 3098 1303 3102 1307
rect 3105 1303 3109 1307
rect 3094 1268 3098 1272
rect 3102 1198 3106 1202
rect 3098 1103 3102 1107
rect 3105 1103 3109 1107
rect 3206 1468 3210 1472
rect 3150 1458 3154 1462
rect 3230 1458 3234 1462
rect 3254 1458 3258 1462
rect 3150 1418 3154 1422
rect 3134 1338 3138 1342
rect 3198 1428 3202 1432
rect 3182 1408 3186 1412
rect 3190 1388 3194 1392
rect 3262 1408 3266 1412
rect 3190 1368 3194 1372
rect 3214 1368 3218 1372
rect 3198 1338 3202 1342
rect 3222 1338 3226 1342
rect 3142 1328 3146 1332
rect 3190 1328 3194 1332
rect 3150 1298 3154 1302
rect 3126 1288 3130 1292
rect 3150 1268 3154 1272
rect 3222 1318 3226 1322
rect 3254 1318 3258 1322
rect 3158 1248 3162 1252
rect 3166 1238 3170 1242
rect 3150 1188 3154 1192
rect 3198 1308 3202 1312
rect 3238 1308 3242 1312
rect 3182 1248 3186 1252
rect 3214 1298 3218 1302
rect 3230 1288 3234 1292
rect 3246 1298 3250 1302
rect 3286 1358 3290 1362
rect 3286 1318 3290 1322
rect 3262 1278 3266 1282
rect 3254 1268 3258 1272
rect 3206 1248 3210 1252
rect 3230 1248 3234 1252
rect 3238 1248 3242 1252
rect 3174 1158 3178 1162
rect 3126 1108 3130 1112
rect 3118 1058 3122 1062
rect 3142 1058 3146 1062
rect 3110 1028 3114 1032
rect 3094 998 3098 1002
rect 3094 938 3098 942
rect 3214 1138 3218 1142
rect 3206 1128 3210 1132
rect 3230 1128 3234 1132
rect 3174 1118 3178 1122
rect 3222 1118 3226 1122
rect 3238 1098 3242 1102
rect 3182 1068 3186 1072
rect 3190 1038 3194 1042
rect 3166 978 3170 982
rect 3126 968 3130 972
rect 3118 948 3122 952
rect 3110 928 3114 932
rect 3098 903 3102 907
rect 3105 903 3109 907
rect 3118 898 3122 902
rect 3102 888 3106 892
rect 3174 958 3178 962
rect 3174 948 3178 952
rect 3206 948 3210 952
rect 3134 928 3138 932
rect 3158 928 3162 932
rect 3150 888 3154 892
rect 3126 858 3130 862
rect 3174 878 3178 882
rect 3190 868 3194 872
rect 3134 848 3138 852
rect 3158 848 3162 852
rect 3118 838 3122 842
rect 3110 818 3114 822
rect 3054 778 3058 782
rect 3038 768 3042 772
rect 3022 758 3026 762
rect 3046 758 3050 762
rect 3006 748 3010 752
rect 3006 728 3010 732
rect 3102 758 3106 762
rect 3126 818 3130 822
rect 3166 818 3170 822
rect 3070 748 3074 752
rect 2958 608 2962 612
rect 2966 578 2970 582
rect 2926 568 2930 572
rect 2918 538 2922 542
rect 2878 498 2882 502
rect 2862 488 2866 492
rect 2814 478 2818 482
rect 2862 478 2866 482
rect 2798 468 2802 472
rect 2822 468 2826 472
rect 2774 448 2778 452
rect 2774 408 2778 412
rect 2774 378 2778 382
rect 2806 458 2810 462
rect 2830 458 2834 462
rect 2846 458 2850 462
rect 2814 448 2818 452
rect 2830 448 2834 452
rect 2790 398 2794 402
rect 2814 388 2818 392
rect 2846 388 2850 392
rect 2806 368 2810 372
rect 2798 358 2802 362
rect 2782 348 2786 352
rect 2814 348 2818 352
rect 2718 338 2722 342
rect 2774 338 2778 342
rect 2734 298 2738 302
rect 2606 258 2610 262
rect 2702 258 2706 262
rect 2510 248 2514 252
rect 2494 228 2498 232
rect 2446 208 2450 212
rect 2294 178 2298 182
rect 2326 178 2330 182
rect 2278 158 2282 162
rect 2310 168 2314 172
rect 2326 158 2330 162
rect 2342 158 2346 162
rect 2286 148 2290 152
rect 2318 148 2322 152
rect 2430 168 2434 172
rect 2222 138 2226 142
rect 2246 138 2250 142
rect 2270 138 2274 142
rect 2374 138 2378 142
rect 2254 128 2258 132
rect 2278 128 2282 132
rect 2318 128 2322 132
rect 2430 128 2434 132
rect 2334 118 2338 122
rect 2446 88 2450 92
rect 2206 78 2210 82
rect 2238 78 2242 82
rect 2350 78 2354 82
rect 2478 78 2482 82
rect 2526 218 2530 222
rect 2510 158 2514 162
rect 2586 203 2590 207
rect 2593 203 2597 207
rect 2678 238 2682 242
rect 2694 238 2698 242
rect 2686 198 2690 202
rect 2742 258 2746 262
rect 2702 188 2706 192
rect 2718 188 2722 192
rect 2654 178 2658 182
rect 2726 178 2730 182
rect 2638 168 2642 172
rect 2686 168 2690 172
rect 2678 158 2682 162
rect 2718 168 2722 172
rect 2606 148 2610 152
rect 2662 148 2666 152
rect 2702 138 2706 142
rect 2678 128 2682 132
rect 2686 118 2690 122
rect 2734 168 2738 172
rect 2862 418 2866 422
rect 2918 498 2922 502
rect 2902 488 2906 492
rect 2886 418 2890 422
rect 2878 378 2882 382
rect 2854 348 2858 352
rect 2870 348 2874 352
rect 2798 318 2802 322
rect 2758 308 2762 312
rect 2830 288 2834 292
rect 2774 278 2778 282
rect 2790 278 2794 282
rect 2806 278 2810 282
rect 2750 198 2754 202
rect 2878 308 2882 312
rect 2862 288 2866 292
rect 2790 228 2794 232
rect 2854 228 2858 232
rect 2766 198 2770 202
rect 2758 168 2762 172
rect 2782 188 2786 192
rect 2798 168 2802 172
rect 2822 168 2826 172
rect 2830 168 2834 172
rect 2854 168 2858 172
rect 2870 158 2874 162
rect 2782 148 2786 152
rect 2806 148 2810 152
rect 2822 148 2826 152
rect 2734 128 2738 132
rect 2614 98 2618 102
rect 2542 88 2546 92
rect 2678 78 2682 82
rect 2102 58 2106 62
rect 2166 58 2170 62
rect 2254 58 2258 62
rect 2286 58 2290 62
rect 2382 58 2386 62
rect 2446 58 2450 62
rect 2478 58 2482 62
rect 2702 68 2706 72
rect 494 48 498 52
rect 654 48 658 52
rect 782 48 786 52
rect 942 48 946 52
rect 958 48 962 52
rect 1390 48 1394 52
rect 1526 48 1530 52
rect 1798 48 1802 52
rect 2630 58 2634 62
rect 2670 58 2674 62
rect 2782 138 2786 142
rect 2862 138 2866 142
rect 2846 118 2850 122
rect 2790 88 2794 92
rect 2750 78 2754 82
rect 2766 68 2770 72
rect 2822 68 2826 72
rect 2742 58 2746 62
rect 2654 48 2658 52
rect 2686 48 2690 52
rect 2734 48 2738 52
rect 950 38 954 42
rect 2598 38 2602 42
rect 2862 108 2866 112
rect 2838 98 2842 102
rect 2846 68 2850 72
rect 2830 58 2834 62
rect 2902 318 2906 322
rect 3118 728 3122 732
rect 3078 718 3082 722
rect 3098 703 3102 707
rect 3105 703 3109 707
rect 3062 688 3066 692
rect 3110 668 3114 672
rect 3182 838 3186 842
rect 3174 778 3178 782
rect 3134 768 3138 772
rect 3150 758 3154 762
rect 3174 758 3178 762
rect 3214 928 3218 932
rect 3206 898 3210 902
rect 3214 748 3218 752
rect 3182 738 3186 742
rect 3150 728 3154 732
rect 3174 728 3178 732
rect 3142 688 3146 692
rect 3014 658 3018 662
rect 3054 658 3058 662
rect 3078 658 3082 662
rect 3118 658 3122 662
rect 3022 648 3026 652
rect 3054 638 3058 642
rect 3006 628 3010 632
rect 2998 608 3002 612
rect 3014 588 3018 592
rect 3046 588 3050 592
rect 3022 578 3026 582
rect 2990 568 2994 572
rect 2958 548 2962 552
rect 2950 538 2954 542
rect 2958 528 2962 532
rect 2950 518 2954 522
rect 2934 438 2938 442
rect 2966 478 2970 482
rect 2982 458 2986 462
rect 2958 408 2962 412
rect 2974 408 2978 412
rect 2990 438 2994 442
rect 2990 418 2994 422
rect 2974 358 2978 362
rect 2982 358 2986 362
rect 2966 348 2970 352
rect 2982 348 2986 352
rect 3038 498 3042 502
rect 3038 478 3042 482
rect 3166 678 3170 682
rect 3350 1488 3354 1492
rect 3318 1468 3322 1472
rect 3430 1558 3434 1562
rect 3414 1528 3418 1532
rect 3510 1668 3514 1672
rect 3494 1578 3498 1582
rect 3470 1558 3474 1562
rect 3526 1558 3530 1562
rect 3638 1838 3642 1842
rect 3614 1818 3618 1822
rect 3610 1803 3614 1807
rect 3617 1803 3621 1807
rect 3838 1938 3842 1942
rect 3830 1928 3834 1932
rect 3678 1878 3682 1882
rect 3806 1878 3810 1882
rect 3814 1878 3818 1882
rect 3654 1858 3658 1862
rect 3734 1858 3738 1862
rect 3670 1848 3674 1852
rect 3718 1838 3722 1842
rect 3646 1788 3650 1792
rect 3606 1778 3610 1782
rect 3662 1778 3666 1782
rect 3630 1758 3634 1762
rect 3646 1748 3650 1752
rect 3662 1748 3666 1752
rect 3702 1748 3706 1752
rect 3606 1688 3610 1692
rect 3646 1688 3650 1692
rect 3542 1648 3546 1652
rect 3646 1678 3650 1682
rect 3790 1798 3794 1802
rect 3750 1788 3754 1792
rect 3838 1898 3842 1902
rect 3830 1848 3834 1852
rect 3782 1778 3786 1782
rect 3806 1778 3810 1782
rect 3830 1768 3834 1772
rect 3854 1948 3858 1952
rect 3870 1948 3874 1952
rect 3862 1928 3866 1932
rect 3870 1898 3874 1902
rect 3870 1878 3874 1882
rect 3854 1848 3858 1852
rect 3918 1968 3922 1972
rect 3902 1958 3906 1962
rect 3950 1958 3954 1962
rect 3910 1948 3914 1952
rect 3998 2028 4002 2032
rect 3982 1978 3986 1982
rect 3998 1958 4002 1962
rect 3894 1928 3898 1932
rect 3958 1928 3962 1932
rect 3934 1908 3938 1912
rect 3886 1898 3890 1902
rect 3878 1868 3882 1872
rect 3774 1748 3778 1752
rect 3806 1748 3810 1752
rect 3838 1748 3842 1752
rect 3662 1728 3666 1732
rect 3686 1728 3690 1732
rect 3750 1728 3754 1732
rect 3638 1648 3642 1652
rect 3582 1638 3586 1642
rect 3630 1638 3634 1642
rect 3610 1603 3614 1607
rect 3617 1603 3621 1607
rect 3566 1578 3570 1582
rect 3582 1578 3586 1582
rect 3622 1578 3626 1582
rect 3614 1558 3618 1562
rect 3534 1548 3538 1552
rect 3542 1538 3546 1542
rect 3566 1538 3570 1542
rect 3590 1538 3594 1542
rect 3478 1528 3482 1532
rect 3390 1488 3394 1492
rect 3398 1488 3402 1492
rect 3406 1468 3410 1472
rect 3446 1468 3450 1472
rect 3454 1468 3458 1472
rect 3374 1458 3378 1462
rect 3398 1458 3402 1462
rect 3358 1448 3362 1452
rect 3422 1448 3426 1452
rect 3334 1428 3338 1432
rect 3334 1378 3338 1382
rect 3318 1348 3322 1352
rect 3294 1248 3298 1252
rect 3302 1238 3306 1242
rect 3286 1198 3290 1202
rect 3294 1188 3298 1192
rect 3286 1178 3290 1182
rect 3270 1148 3274 1152
rect 3254 1118 3258 1122
rect 3262 1098 3266 1102
rect 3262 1078 3266 1082
rect 3262 1058 3266 1062
rect 3254 958 3258 962
rect 3278 1048 3282 1052
rect 3270 948 3274 952
rect 3270 938 3274 942
rect 3310 1168 3314 1172
rect 3302 1138 3306 1142
rect 3310 1138 3314 1142
rect 3294 1078 3298 1082
rect 3302 958 3306 962
rect 3334 1268 3338 1272
rect 3358 1268 3362 1272
rect 3358 1228 3362 1232
rect 3382 1428 3386 1432
rect 3374 1358 3378 1362
rect 3470 1448 3474 1452
rect 3534 1518 3538 1522
rect 3510 1488 3514 1492
rect 3542 1488 3546 1492
rect 3526 1468 3530 1472
rect 3582 1488 3586 1492
rect 3646 1548 3650 1552
rect 3686 1698 3690 1702
rect 3726 1688 3730 1692
rect 3702 1668 3706 1672
rect 3798 1728 3802 1732
rect 3758 1718 3762 1722
rect 3790 1708 3794 1712
rect 3758 1678 3762 1682
rect 3766 1668 3770 1672
rect 3670 1638 3674 1642
rect 3662 1528 3666 1532
rect 3654 1488 3658 1492
rect 3670 1508 3674 1512
rect 3670 1498 3674 1502
rect 3518 1458 3522 1462
rect 3550 1458 3554 1462
rect 3574 1458 3578 1462
rect 3606 1458 3610 1462
rect 3478 1428 3482 1432
rect 3454 1398 3458 1402
rect 3430 1368 3434 1372
rect 3414 1358 3418 1362
rect 3438 1358 3442 1362
rect 3494 1398 3498 1402
rect 3382 1338 3386 1342
rect 3502 1338 3506 1342
rect 3414 1328 3418 1332
rect 3390 1298 3394 1302
rect 3382 1288 3386 1292
rect 3374 1238 3378 1242
rect 3350 1218 3354 1222
rect 3366 1218 3370 1222
rect 3326 1208 3330 1212
rect 3326 1178 3330 1182
rect 3334 1148 3338 1152
rect 3374 1148 3378 1152
rect 3326 1118 3330 1122
rect 3358 1108 3362 1112
rect 3366 1088 3370 1092
rect 3382 1078 3386 1082
rect 3350 1068 3354 1072
rect 3374 1038 3378 1042
rect 3350 968 3354 972
rect 3326 958 3330 962
rect 3318 948 3322 952
rect 3254 928 3258 932
rect 3286 928 3290 932
rect 3246 898 3250 902
rect 3238 878 3242 882
rect 3278 918 3282 922
rect 3254 868 3258 872
rect 3246 858 3250 862
rect 3230 818 3234 822
rect 3262 858 3266 862
rect 3358 958 3362 962
rect 3318 898 3322 902
rect 3310 888 3314 892
rect 3286 858 3290 862
rect 3262 828 3266 832
rect 3294 818 3298 822
rect 3286 798 3290 802
rect 3254 778 3258 782
rect 3270 748 3274 752
rect 3198 728 3202 732
rect 3190 678 3194 682
rect 3150 668 3154 672
rect 3166 668 3170 672
rect 3206 668 3210 672
rect 3118 588 3122 592
rect 3094 578 3098 582
rect 3086 558 3090 562
rect 3070 538 3074 542
rect 3142 548 3146 552
rect 3134 538 3138 542
rect 3150 528 3154 532
rect 3098 503 3102 507
rect 3105 503 3109 507
rect 3110 468 3114 472
rect 3134 468 3138 472
rect 3038 458 3042 462
rect 3014 428 3018 432
rect 3014 388 3018 392
rect 2998 368 3002 372
rect 2998 358 3002 362
rect 2974 338 2978 342
rect 3006 318 3010 322
rect 2998 288 3002 292
rect 2974 278 2978 282
rect 3054 448 3058 452
rect 3182 638 3186 642
rect 3174 628 3178 632
rect 3166 618 3170 622
rect 3222 718 3226 722
rect 3438 1328 3442 1332
rect 3646 1448 3650 1452
rect 3550 1428 3554 1432
rect 3534 1398 3538 1402
rect 3526 1358 3530 1362
rect 3610 1403 3614 1407
rect 3617 1403 3621 1407
rect 3638 1388 3642 1392
rect 3646 1388 3650 1392
rect 3574 1348 3578 1352
rect 3422 1298 3426 1302
rect 3518 1298 3522 1302
rect 3550 1298 3554 1302
rect 3430 1288 3434 1292
rect 3446 1288 3450 1292
rect 3406 1268 3410 1272
rect 3470 1278 3474 1282
rect 3414 1258 3418 1262
rect 3398 1218 3402 1222
rect 3446 1258 3450 1262
rect 3478 1248 3482 1252
rect 3438 1198 3442 1202
rect 3526 1218 3530 1222
rect 3494 1198 3498 1202
rect 3462 1178 3466 1182
rect 3502 1168 3506 1172
rect 3462 1158 3466 1162
rect 3510 1148 3514 1152
rect 3398 1108 3402 1112
rect 3422 1108 3426 1112
rect 3462 1098 3466 1102
rect 3494 1128 3498 1132
rect 3478 1088 3482 1092
rect 3502 1088 3506 1092
rect 3526 1088 3530 1092
rect 3454 1078 3458 1082
rect 3414 1068 3418 1072
rect 3430 1068 3434 1072
rect 3438 1048 3442 1052
rect 3398 1038 3402 1042
rect 3390 1008 3394 1012
rect 3422 978 3426 982
rect 3398 958 3402 962
rect 3414 958 3418 962
rect 3350 868 3354 872
rect 3382 868 3386 872
rect 3374 858 3378 862
rect 3342 838 3346 842
rect 3326 828 3330 832
rect 3310 798 3314 802
rect 3294 788 3298 792
rect 3302 758 3306 762
rect 3326 748 3330 752
rect 3374 778 3378 782
rect 3358 768 3362 772
rect 3334 738 3338 742
rect 3358 738 3362 742
rect 3390 738 3394 742
rect 3350 728 3354 732
rect 3238 688 3242 692
rect 3262 688 3266 692
rect 3310 688 3314 692
rect 3310 678 3314 682
rect 3286 668 3290 672
rect 3214 608 3218 612
rect 3222 608 3226 612
rect 3214 568 3218 572
rect 3198 558 3202 562
rect 3174 548 3178 552
rect 3262 548 3266 552
rect 3182 538 3186 542
rect 3174 508 3178 512
rect 3174 478 3178 482
rect 3254 498 3258 502
rect 3190 468 3194 472
rect 3214 468 3218 472
rect 3126 458 3130 462
rect 3310 598 3314 602
rect 3342 588 3346 592
rect 3318 548 3322 552
rect 3334 548 3338 552
rect 3326 538 3330 542
rect 3406 938 3410 942
rect 3414 878 3418 882
rect 3414 858 3418 862
rect 3406 838 3410 842
rect 3422 828 3426 832
rect 3422 788 3426 792
rect 3406 768 3410 772
rect 3406 758 3410 762
rect 3478 1068 3482 1072
rect 3542 1158 3546 1162
rect 3614 1298 3618 1302
rect 3654 1368 3658 1372
rect 3798 1678 3802 1682
rect 3814 1718 3818 1722
rect 3830 1718 3834 1722
rect 3814 1678 3818 1682
rect 3806 1668 3810 1672
rect 3774 1648 3778 1652
rect 3790 1648 3794 1652
rect 3806 1648 3810 1652
rect 3782 1628 3786 1632
rect 3750 1578 3754 1582
rect 3974 1868 3978 1872
rect 3998 1868 4002 1872
rect 3966 1848 3970 1852
rect 3902 1838 3906 1842
rect 3958 1818 3962 1822
rect 3910 1728 3914 1732
rect 3918 1708 3922 1712
rect 3926 1688 3930 1692
rect 3854 1668 3858 1672
rect 3870 1668 3874 1672
rect 3910 1659 3914 1663
rect 3846 1638 3850 1642
rect 3838 1628 3842 1632
rect 3814 1618 3818 1622
rect 3790 1608 3794 1612
rect 3822 1608 3826 1612
rect 3798 1558 3802 1562
rect 3726 1528 3730 1532
rect 3758 1528 3762 1532
rect 3710 1518 3714 1522
rect 3766 1518 3770 1522
rect 3734 1508 3738 1512
rect 3862 1608 3866 1612
rect 3910 1608 3914 1612
rect 3878 1578 3882 1582
rect 3854 1558 3858 1562
rect 3950 1618 3954 1622
rect 3862 1538 3866 1542
rect 3918 1538 3922 1542
rect 3806 1518 3810 1522
rect 3846 1518 3850 1522
rect 3854 1518 3858 1522
rect 3686 1488 3690 1492
rect 3782 1488 3786 1492
rect 3718 1468 3722 1472
rect 3870 1468 3874 1472
rect 3678 1458 3682 1462
rect 3710 1458 3714 1462
rect 3686 1448 3690 1452
rect 3734 1448 3738 1452
rect 3662 1358 3666 1362
rect 3678 1348 3682 1352
rect 3686 1348 3690 1352
rect 3662 1338 3666 1342
rect 3646 1328 3650 1332
rect 3822 1398 3826 1402
rect 3822 1388 3826 1392
rect 3718 1368 3722 1372
rect 3798 1368 3802 1372
rect 3902 1468 3906 1472
rect 3934 1488 3938 1492
rect 3974 1798 3978 1802
rect 3982 1788 3986 1792
rect 3982 1768 3986 1772
rect 3990 1748 3994 1752
rect 4086 2078 4090 2082
rect 4046 2068 4050 2072
rect 4070 2068 4074 2072
rect 4014 2058 4018 2062
rect 4030 1988 4034 1992
rect 4022 1948 4026 1952
rect 4014 1788 4018 1792
rect 4022 1778 4026 1782
rect 4014 1758 4018 1762
rect 4038 1958 4042 1962
rect 4078 2048 4082 2052
rect 4110 2118 4114 2122
rect 4114 2103 4118 2107
rect 4121 2103 4125 2107
rect 4110 2078 4114 2082
rect 4118 2078 4122 2082
rect 4110 2068 4114 2072
rect 4062 2018 4066 2022
rect 4078 2008 4082 2012
rect 4094 2008 4098 2012
rect 4102 1978 4106 1982
rect 4166 2408 4170 2412
rect 4230 2738 4234 2742
rect 4230 2668 4234 2672
rect 4270 2758 4274 2762
rect 4254 2728 4258 2732
rect 4254 2718 4258 2722
rect 4294 2688 4298 2692
rect 4326 2718 4330 2722
rect 4318 2688 4322 2692
rect 4502 3268 4506 3272
rect 4510 3258 4514 3262
rect 4526 3258 4530 3262
rect 4486 3208 4490 3212
rect 4502 3148 4506 3152
rect 4518 3148 4522 3152
rect 4374 3068 4378 3072
rect 4406 3068 4410 3072
rect 4374 3038 4378 3042
rect 4494 3128 4498 3132
rect 4422 3098 4426 3102
rect 4462 3098 4466 3102
rect 4510 3098 4514 3102
rect 4430 3068 4434 3072
rect 4454 3058 4458 3062
rect 4398 2948 4402 2952
rect 4414 2948 4418 2952
rect 4406 2938 4410 2942
rect 4366 2888 4370 2892
rect 4470 3048 4474 3052
rect 4446 3038 4450 3042
rect 4494 3058 4498 3062
rect 4634 3403 4638 3407
rect 4641 3403 4645 3407
rect 4638 3378 4642 3382
rect 4630 3368 4634 3372
rect 4582 3318 4586 3322
rect 4590 3318 4594 3322
rect 4598 3308 4602 3312
rect 4638 3308 4642 3312
rect 4582 3278 4586 3282
rect 4606 3278 4610 3282
rect 4574 3268 4578 3272
rect 4566 3228 4570 3232
rect 4550 3218 4554 3222
rect 4534 3188 4538 3192
rect 4534 3148 4538 3152
rect 4518 3058 4522 3062
rect 4494 3048 4498 3052
rect 4518 3028 4522 3032
rect 4478 3008 4482 3012
rect 4486 3008 4490 3012
rect 4454 2998 4458 3002
rect 4446 2938 4450 2942
rect 4438 2868 4442 2872
rect 4566 3138 4570 3142
rect 4558 3078 4562 3082
rect 4582 3078 4586 3082
rect 4550 3068 4554 3072
rect 4566 3048 4570 3052
rect 4542 3038 4546 3042
rect 4534 2998 4538 3002
rect 4526 2978 4530 2982
rect 4526 2958 4530 2962
rect 4478 2948 4482 2952
rect 4622 3258 4626 3262
rect 4638 3258 4642 3262
rect 4606 3228 4610 3232
rect 4634 3203 4638 3207
rect 4641 3203 4645 3207
rect 4694 3498 4698 3502
rect 4670 3478 4674 3482
rect 4710 3518 4714 3522
rect 4694 3468 4698 3472
rect 4670 3458 4674 3462
rect 4662 3438 4666 3442
rect 4686 3348 4690 3352
rect 4718 3458 4722 3462
rect 4774 3688 4778 3692
rect 4830 3688 4834 3692
rect 4966 3818 4970 3822
rect 4982 3788 4986 3792
rect 4990 3778 4994 3782
rect 4998 3758 5002 3762
rect 4982 3748 4986 3752
rect 4902 3728 4906 3732
rect 4918 3708 4922 3712
rect 4774 3678 4778 3682
rect 4750 3668 4754 3672
rect 4822 3668 4826 3672
rect 4774 3608 4778 3612
rect 4878 3678 4882 3682
rect 4894 3668 4898 3672
rect 4958 3688 4962 3692
rect 4926 3678 4930 3682
rect 4846 3658 4850 3662
rect 4878 3658 4882 3662
rect 4910 3658 4914 3662
rect 4822 3648 4826 3652
rect 4806 3638 4810 3642
rect 4838 3638 4842 3642
rect 4798 3588 4802 3592
rect 4758 3568 4762 3572
rect 4734 3528 4738 3532
rect 4750 3548 4754 3552
rect 4750 3508 4754 3512
rect 4750 3458 4754 3462
rect 4774 3508 4778 3512
rect 4782 3478 4786 3482
rect 4798 3478 4802 3482
rect 4766 3458 4770 3462
rect 4742 3448 4746 3452
rect 4758 3448 4762 3452
rect 4758 3428 4762 3432
rect 4758 3358 4762 3362
rect 4718 3348 4722 3352
rect 4734 3348 4738 3352
rect 4702 3338 4706 3342
rect 4750 3338 4754 3342
rect 4662 3318 4666 3322
rect 4662 3278 4666 3282
rect 4686 3198 4690 3202
rect 4694 3188 4698 3192
rect 4654 3158 4658 3162
rect 4670 3138 4674 3142
rect 4686 3138 4690 3142
rect 4590 3048 4594 3052
rect 4606 3048 4610 3052
rect 4654 3108 4658 3112
rect 4678 3098 4682 3102
rect 4654 3068 4658 3072
rect 4638 3058 4642 3062
rect 4630 3048 4634 3052
rect 4622 3038 4626 3042
rect 4766 3308 4770 3312
rect 4742 3278 4746 3282
rect 4766 3278 4770 3282
rect 4710 3258 4714 3262
rect 4798 3438 4802 3442
rect 4782 3358 4786 3362
rect 4846 3558 4850 3562
rect 4870 3588 4874 3592
rect 4894 3578 4898 3582
rect 4886 3548 4890 3552
rect 4854 3538 4858 3542
rect 4902 3548 4906 3552
rect 4942 3588 4946 3592
rect 4926 3568 4930 3572
rect 4926 3548 4930 3552
rect 4934 3528 4938 3532
rect 4974 3718 4978 3722
rect 4990 3698 4994 3702
rect 4982 3668 4986 3672
rect 4966 3518 4970 3522
rect 4926 3498 4930 3502
rect 4982 3498 4986 3502
rect 4846 3458 4850 3462
rect 4902 3458 4906 3462
rect 4910 3458 4914 3462
rect 4918 3458 4922 3462
rect 4846 3368 4850 3372
rect 4822 3348 4826 3352
rect 4846 3348 4850 3352
rect 4886 3348 4890 3352
rect 4806 3278 4810 3282
rect 4822 3338 4826 3342
rect 4894 3338 4898 3342
rect 4822 3328 4826 3332
rect 4790 3258 4794 3262
rect 4806 3258 4810 3262
rect 4814 3228 4818 3232
rect 4774 3208 4778 3212
rect 4702 3178 4706 3182
rect 4726 3168 4730 3172
rect 4702 3158 4706 3162
rect 4734 3158 4738 3162
rect 4782 3158 4786 3162
rect 4798 3158 4802 3162
rect 4750 3138 4754 3142
rect 4782 3138 4786 3142
rect 4718 3128 4722 3132
rect 4718 3098 4722 3102
rect 4798 3078 4802 3082
rect 4830 3238 4834 3242
rect 4870 3298 4874 3302
rect 4862 3288 4866 3292
rect 4886 3278 4890 3282
rect 4838 3198 4842 3202
rect 4846 3178 4850 3182
rect 4822 3148 4826 3152
rect 4838 3088 4842 3092
rect 4694 3068 4698 3072
rect 4702 3058 4706 3062
rect 4726 3038 4730 3042
rect 4614 3028 4618 3032
rect 4574 3018 4578 3022
rect 4598 3018 4602 3022
rect 4606 3018 4610 3022
rect 4622 3018 4626 3022
rect 4654 3018 4658 3022
rect 4550 2968 4554 2972
rect 4582 2958 4586 2962
rect 4606 2958 4610 2962
rect 4558 2948 4562 2952
rect 4606 2928 4610 2932
rect 4574 2918 4578 2922
rect 4598 2918 4602 2922
rect 4462 2908 4466 2912
rect 4558 2908 4562 2912
rect 4470 2868 4474 2872
rect 4518 2868 4522 2872
rect 4350 2858 4354 2862
rect 4430 2858 4434 2862
rect 4446 2858 4450 2862
rect 4454 2858 4458 2862
rect 4550 2858 4554 2862
rect 4462 2848 4466 2852
rect 4382 2808 4386 2812
rect 4510 2828 4514 2832
rect 4494 2808 4498 2812
rect 4478 2778 4482 2782
rect 4494 2768 4498 2772
rect 4334 2668 4338 2672
rect 4350 2668 4354 2672
rect 4374 2668 4378 2672
rect 4246 2648 4250 2652
rect 4238 2628 4242 2632
rect 4214 2618 4218 2622
rect 4206 2588 4210 2592
rect 4198 2568 4202 2572
rect 4190 2548 4194 2552
rect 4198 2508 4202 2512
rect 4246 2558 4250 2562
rect 4422 2728 4426 2732
rect 4398 2698 4402 2702
rect 4422 2678 4426 2682
rect 4534 2798 4538 2802
rect 4526 2748 4530 2752
rect 4590 2888 4594 2892
rect 4614 2878 4618 2882
rect 4598 2868 4602 2872
rect 4566 2828 4570 2832
rect 4614 2858 4618 2862
rect 4606 2818 4610 2822
rect 4574 2758 4578 2762
rect 4582 2748 4586 2752
rect 4606 2738 4610 2742
rect 4558 2728 4562 2732
rect 4582 2728 4586 2732
rect 4590 2728 4594 2732
rect 4542 2708 4546 2712
rect 4606 2728 4610 2732
rect 4598 2718 4602 2722
rect 4634 3003 4638 3007
rect 4641 3003 4645 3007
rect 4654 2998 4658 3002
rect 4654 2988 4658 2992
rect 4774 3028 4778 3032
rect 4686 3018 4690 3022
rect 4702 3008 4706 3012
rect 4814 2998 4818 3002
rect 4766 2988 4770 2992
rect 4790 2988 4794 2992
rect 4798 2988 4802 2992
rect 4726 2978 4730 2982
rect 4718 2968 4722 2972
rect 4686 2958 4690 2962
rect 4718 2958 4722 2962
rect 4678 2938 4682 2942
rect 4694 2938 4698 2942
rect 4686 2918 4690 2922
rect 4662 2908 4666 2912
rect 4678 2898 4682 2902
rect 4694 2898 4698 2902
rect 4670 2878 4674 2882
rect 4638 2868 4642 2872
rect 4662 2868 4666 2872
rect 4670 2858 4674 2862
rect 4630 2848 4634 2852
rect 4654 2828 4658 2832
rect 4634 2803 4638 2807
rect 4641 2803 4645 2807
rect 4646 2778 4650 2782
rect 4670 2808 4674 2812
rect 4662 2758 4666 2762
rect 4678 2738 4682 2742
rect 4686 2738 4690 2742
rect 4678 2728 4682 2732
rect 4590 2688 4594 2692
rect 4622 2688 4626 2692
rect 4662 2688 4666 2692
rect 4446 2668 4450 2672
rect 4486 2668 4490 2672
rect 4518 2668 4522 2672
rect 4358 2658 4362 2662
rect 4382 2658 4386 2662
rect 4398 2648 4402 2652
rect 4310 2588 4314 2592
rect 4382 2578 4386 2582
rect 4294 2568 4298 2572
rect 4214 2528 4218 2532
rect 4246 2518 4250 2522
rect 4214 2498 4218 2502
rect 4198 2458 4202 2462
rect 4230 2368 4234 2372
rect 4198 2358 4202 2362
rect 4214 2358 4218 2362
rect 4190 2348 4194 2352
rect 4206 2348 4210 2352
rect 4174 2318 4178 2322
rect 4262 2488 4266 2492
rect 4278 2368 4282 2372
rect 4238 2348 4242 2352
rect 4262 2328 4266 2332
rect 4198 2318 4202 2322
rect 4190 2308 4194 2312
rect 4174 2298 4178 2302
rect 4198 2288 4202 2292
rect 4190 2258 4194 2262
rect 4174 2208 4178 2212
rect 4222 2318 4226 2322
rect 4238 2318 4242 2322
rect 4286 2288 4290 2292
rect 4438 2638 4442 2642
rect 4454 2638 4458 2642
rect 4478 2638 4482 2642
rect 4446 2618 4450 2622
rect 4350 2548 4354 2552
rect 4406 2548 4410 2552
rect 4326 2538 4330 2542
rect 4310 2528 4314 2532
rect 4310 2458 4314 2462
rect 4390 2538 4394 2542
rect 4342 2498 4346 2502
rect 4350 2468 4354 2472
rect 4326 2458 4330 2462
rect 4342 2458 4346 2462
rect 4334 2438 4338 2442
rect 4342 2358 4346 2362
rect 4374 2468 4378 2472
rect 4366 2458 4370 2462
rect 4374 2438 4378 2442
rect 4366 2408 4370 2412
rect 4382 2398 4386 2402
rect 4382 2378 4386 2382
rect 4366 2348 4370 2352
rect 4318 2308 4322 2312
rect 4342 2298 4346 2302
rect 4334 2288 4338 2292
rect 4246 2258 4250 2262
rect 4286 2258 4290 2262
rect 4294 2258 4298 2262
rect 4214 2248 4218 2252
rect 4214 2238 4218 2242
rect 4326 2248 4330 2252
rect 4262 2238 4266 2242
rect 4294 2238 4298 2242
rect 4254 2228 4258 2232
rect 4366 2318 4370 2322
rect 4366 2298 4370 2302
rect 4374 2268 4378 2272
rect 4398 2468 4402 2472
rect 4470 2578 4474 2582
rect 4430 2558 4434 2562
rect 4462 2558 4466 2562
rect 4446 2538 4450 2542
rect 4422 2488 4426 2492
rect 4446 2468 4450 2472
rect 4614 2678 4618 2682
rect 4590 2668 4594 2672
rect 4510 2658 4514 2662
rect 4582 2658 4586 2662
rect 4494 2528 4498 2532
rect 4486 2498 4490 2502
rect 4478 2488 4482 2492
rect 4470 2478 4474 2482
rect 4478 2478 4482 2482
rect 4518 2648 4522 2652
rect 4566 2648 4570 2652
rect 4574 2608 4578 2612
rect 4574 2578 4578 2582
rect 4550 2568 4554 2572
rect 4582 2568 4586 2572
rect 4582 2558 4586 2562
rect 4526 2538 4530 2542
rect 4542 2528 4546 2532
rect 4678 2668 4682 2672
rect 4646 2648 4650 2652
rect 4634 2603 4638 2607
rect 4641 2603 4645 2607
rect 4622 2598 4626 2602
rect 4638 2568 4642 2572
rect 4622 2548 4626 2552
rect 4590 2538 4594 2542
rect 4598 2538 4602 2542
rect 4614 2538 4618 2542
rect 4582 2518 4586 2522
rect 4558 2498 4562 2502
rect 4510 2458 4514 2462
rect 4534 2458 4538 2462
rect 4462 2448 4466 2452
rect 4470 2418 4474 2422
rect 4446 2388 4450 2392
rect 4470 2388 4474 2392
rect 4478 2358 4482 2362
rect 4494 2448 4498 2452
rect 4542 2448 4546 2452
rect 4630 2488 4634 2492
rect 4646 2488 4650 2492
rect 4638 2478 4642 2482
rect 4670 2648 4674 2652
rect 4686 2618 4690 2622
rect 4662 2468 4666 2472
rect 4598 2458 4602 2462
rect 4686 2458 4690 2462
rect 4678 2448 4682 2452
rect 4574 2438 4578 2442
rect 4510 2428 4514 2432
rect 4550 2428 4554 2432
rect 4518 2398 4522 2402
rect 4518 2368 4522 2372
rect 4510 2358 4514 2362
rect 4526 2358 4530 2362
rect 4542 2358 4546 2362
rect 4414 2338 4418 2342
rect 4462 2338 4466 2342
rect 4398 2328 4402 2332
rect 4414 2328 4418 2332
rect 4430 2318 4434 2322
rect 4422 2308 4426 2312
rect 4414 2228 4418 2232
rect 4390 2218 4394 2222
rect 4278 2198 4282 2202
rect 4350 2198 4354 2202
rect 4334 2188 4338 2192
rect 4150 2168 4154 2172
rect 4286 2168 4290 2172
rect 4158 2158 4162 2162
rect 4190 2158 4194 2162
rect 4222 2158 4226 2162
rect 4254 2158 4258 2162
rect 4182 2148 4186 2152
rect 4142 2138 4146 2142
rect 4166 2138 4170 2142
rect 4166 2128 4170 2132
rect 4174 2098 4178 2102
rect 4166 2078 4170 2082
rect 4126 2058 4130 2062
rect 4134 2008 4138 2012
rect 4110 1958 4114 1962
rect 4046 1948 4050 1952
rect 4078 1948 4082 1952
rect 4102 1928 4106 1932
rect 4126 1928 4130 1932
rect 4054 1908 4058 1912
rect 4114 1903 4118 1907
rect 4121 1903 4125 1907
rect 4070 1898 4074 1902
rect 4102 1898 4106 1902
rect 4062 1888 4066 1892
rect 4078 1888 4082 1892
rect 4046 1818 4050 1822
rect 4094 1868 4098 1872
rect 4054 1788 4058 1792
rect 4038 1758 4042 1762
rect 4030 1748 4034 1752
rect 4094 1848 4098 1852
rect 4094 1798 4098 1802
rect 4062 1778 4066 1782
rect 4086 1778 4090 1782
rect 3998 1708 4002 1712
rect 3982 1698 3986 1702
rect 4022 1688 4026 1692
rect 3990 1678 3994 1682
rect 3998 1678 4002 1682
rect 3966 1658 3970 1662
rect 3990 1658 3994 1662
rect 3974 1638 3978 1642
rect 4070 1698 4074 1702
rect 4118 1838 4122 1842
rect 4102 1748 4106 1752
rect 4118 1728 4122 1732
rect 4102 1718 4106 1722
rect 4114 1703 4118 1707
rect 4121 1703 4125 1707
rect 4110 1688 4114 1692
rect 4086 1678 4090 1682
rect 4054 1658 4058 1662
rect 4014 1638 4018 1642
rect 4062 1628 4066 1632
rect 4022 1598 4026 1602
rect 4054 1588 4058 1592
rect 3974 1548 3978 1552
rect 4054 1548 4058 1552
rect 3958 1538 3962 1542
rect 3990 1538 3994 1542
rect 3966 1508 3970 1512
rect 3958 1478 3962 1482
rect 3990 1488 3994 1492
rect 3998 1488 4002 1492
rect 3974 1468 3978 1472
rect 3862 1458 3866 1462
rect 3886 1458 3890 1462
rect 3910 1458 3914 1462
rect 3934 1458 3938 1462
rect 3862 1448 3866 1452
rect 3854 1428 3858 1432
rect 3854 1408 3858 1412
rect 3838 1368 3842 1372
rect 3830 1358 3834 1362
rect 3750 1348 3754 1352
rect 3766 1338 3770 1342
rect 3838 1338 3842 1342
rect 3734 1328 3738 1332
rect 3686 1298 3690 1302
rect 3702 1298 3706 1302
rect 3798 1288 3802 1292
rect 3806 1288 3810 1292
rect 3694 1268 3698 1272
rect 3742 1268 3746 1272
rect 3598 1258 3602 1262
rect 3638 1258 3642 1262
rect 3646 1248 3650 1252
rect 3558 1238 3562 1242
rect 3582 1238 3586 1242
rect 3590 1238 3594 1242
rect 3606 1238 3610 1242
rect 3646 1238 3650 1242
rect 3654 1238 3658 1242
rect 3574 1228 3578 1232
rect 3558 1198 3562 1202
rect 3610 1203 3614 1207
rect 3617 1203 3621 1207
rect 3574 1148 3578 1152
rect 3598 1148 3602 1152
rect 3638 1148 3642 1152
rect 3590 1098 3594 1102
rect 3550 1078 3554 1082
rect 3590 1058 3594 1062
rect 3462 948 3466 952
rect 3446 878 3450 882
rect 3446 868 3450 872
rect 3438 828 3442 832
rect 3502 1008 3506 1012
rect 3478 988 3482 992
rect 3494 958 3498 962
rect 3470 938 3474 942
rect 3470 888 3474 892
rect 3502 888 3506 892
rect 3462 878 3466 882
rect 3486 878 3490 882
rect 3502 868 3506 872
rect 3462 828 3466 832
rect 3486 858 3490 862
rect 3478 788 3482 792
rect 3430 768 3434 772
rect 3414 708 3418 712
rect 3382 688 3386 692
rect 3430 728 3434 732
rect 3470 758 3474 762
rect 3446 688 3450 692
rect 3382 598 3386 602
rect 3398 598 3402 602
rect 3366 568 3370 572
rect 3406 588 3410 592
rect 3430 588 3434 592
rect 3454 598 3458 602
rect 3438 578 3442 582
rect 3390 568 3394 572
rect 3438 568 3442 572
rect 3374 558 3378 562
rect 3358 548 3362 552
rect 3398 558 3402 562
rect 3454 558 3458 562
rect 3406 548 3410 552
rect 3430 548 3434 552
rect 3446 548 3450 552
rect 3334 528 3338 532
rect 3342 528 3346 532
rect 3334 518 3338 522
rect 3278 498 3282 502
rect 3270 478 3274 482
rect 3294 468 3298 472
rect 3254 458 3258 462
rect 3102 438 3106 442
rect 3102 418 3106 422
rect 3174 428 3178 432
rect 3038 398 3042 402
rect 3150 398 3154 402
rect 3150 388 3154 392
rect 3046 378 3050 382
rect 3206 368 3210 372
rect 3278 368 3282 372
rect 3310 368 3314 372
rect 3054 358 3058 362
rect 3030 338 3034 342
rect 3022 308 3026 312
rect 3190 348 3194 352
rect 3094 338 3098 342
rect 3126 338 3130 342
rect 3014 288 3018 292
rect 2958 268 2962 272
rect 2982 268 2986 272
rect 3030 278 3034 282
rect 3006 258 3010 262
rect 3022 238 3026 242
rect 2894 188 2898 192
rect 2974 228 2978 232
rect 2886 148 2890 152
rect 2894 88 2898 92
rect 2934 148 2938 152
rect 2918 128 2922 132
rect 2902 78 2906 82
rect 3038 228 3042 232
rect 3022 128 3026 132
rect 2982 78 2986 82
rect 3022 78 3026 82
rect 2934 68 2938 72
rect 2942 68 2946 72
rect 2998 58 3002 62
rect 3062 288 3066 292
rect 3158 328 3162 332
rect 3150 318 3154 322
rect 3098 303 3102 307
rect 3105 303 3109 307
rect 3126 298 3130 302
rect 3126 278 3130 282
rect 3070 259 3074 263
rect 3070 238 3074 242
rect 3054 68 3058 72
rect 3166 298 3170 302
rect 3198 288 3202 292
rect 3222 348 3226 352
rect 3278 348 3282 352
rect 3294 348 3298 352
rect 3270 338 3274 342
rect 3366 528 3370 532
rect 3374 518 3378 522
rect 3454 538 3458 542
rect 3414 528 3418 532
rect 3422 508 3426 512
rect 3470 708 3474 712
rect 3478 698 3482 702
rect 3470 638 3474 642
rect 3502 688 3506 692
rect 3494 658 3498 662
rect 3494 648 3498 652
rect 3486 628 3490 632
rect 3478 618 3482 622
rect 3470 568 3474 572
rect 3590 1038 3594 1042
rect 3614 1088 3618 1092
rect 3614 1078 3618 1082
rect 3614 1058 3618 1062
rect 3646 1058 3650 1062
rect 3606 1048 3610 1052
rect 3598 1008 3602 1012
rect 3610 1003 3614 1007
rect 3617 1003 3621 1007
rect 3614 988 3618 992
rect 3550 958 3554 962
rect 3686 1248 3690 1252
rect 3726 1248 3730 1252
rect 3686 1228 3690 1232
rect 3726 1228 3730 1232
rect 3670 1218 3674 1222
rect 3710 1208 3714 1212
rect 3702 1178 3706 1182
rect 3670 1118 3674 1122
rect 3686 1108 3690 1112
rect 3694 1108 3698 1112
rect 3670 1088 3674 1092
rect 3662 1078 3666 1082
rect 3862 1318 3866 1322
rect 3886 1428 3890 1432
rect 3918 1448 3922 1452
rect 3910 1428 3914 1432
rect 3926 1398 3930 1402
rect 3902 1388 3906 1392
rect 3878 1308 3882 1312
rect 3838 1288 3842 1292
rect 3822 1278 3826 1282
rect 3846 1278 3850 1282
rect 3878 1278 3882 1282
rect 3822 1268 3826 1272
rect 3894 1368 3898 1372
rect 3966 1448 3970 1452
rect 3990 1448 3994 1452
rect 3934 1388 3938 1392
rect 3902 1348 3906 1352
rect 3926 1348 3930 1352
rect 3902 1338 3906 1342
rect 3894 1278 3898 1282
rect 3918 1298 3922 1302
rect 3902 1268 3906 1272
rect 3798 1248 3802 1252
rect 3822 1248 3826 1252
rect 3846 1248 3850 1252
rect 3750 1238 3754 1242
rect 3774 1238 3778 1242
rect 3718 1198 3722 1202
rect 3734 1198 3738 1202
rect 3870 1238 3874 1242
rect 3758 1168 3762 1172
rect 3902 1168 3906 1172
rect 3742 1158 3746 1162
rect 3710 1118 3714 1122
rect 3710 1108 3714 1112
rect 3766 1158 3770 1162
rect 3822 1158 3826 1162
rect 3862 1158 3866 1162
rect 3870 1158 3874 1162
rect 3742 1148 3746 1152
rect 3782 1148 3786 1152
rect 3830 1148 3834 1152
rect 3782 1128 3786 1132
rect 3750 1118 3754 1122
rect 3702 1058 3706 1062
rect 3662 1038 3666 1042
rect 3694 1038 3698 1042
rect 3670 1008 3674 1012
rect 3654 988 3658 992
rect 3638 948 3642 952
rect 3550 938 3554 942
rect 3662 938 3666 942
rect 3518 748 3522 752
rect 3638 928 3642 932
rect 3582 878 3586 882
rect 3670 868 3674 872
rect 3734 1088 3738 1092
rect 3774 1088 3778 1092
rect 3742 1078 3746 1082
rect 3734 1058 3738 1062
rect 3742 1038 3746 1042
rect 3726 1018 3730 1022
rect 3734 998 3738 1002
rect 3726 928 3730 932
rect 3686 878 3690 882
rect 3734 868 3738 872
rect 3566 858 3570 862
rect 3614 858 3618 862
rect 3678 858 3682 862
rect 3558 838 3562 842
rect 3678 838 3682 842
rect 3574 818 3578 822
rect 3526 688 3530 692
rect 3526 678 3530 682
rect 3510 618 3514 622
rect 3502 608 3506 612
rect 3478 548 3482 552
rect 3470 508 3474 512
rect 3462 498 3466 502
rect 3486 498 3490 502
rect 3390 488 3394 492
rect 3446 478 3450 482
rect 3462 478 3466 482
rect 3406 468 3410 472
rect 3438 468 3442 472
rect 3454 468 3458 472
rect 3478 438 3482 442
rect 3398 428 3402 432
rect 3374 408 3378 412
rect 3446 398 3450 402
rect 3494 468 3498 472
rect 3526 648 3530 652
rect 3534 638 3538 642
rect 3518 598 3522 602
rect 3566 598 3570 602
rect 3610 803 3614 807
rect 3617 803 3621 807
rect 3702 858 3706 862
rect 3694 798 3698 802
rect 3686 768 3690 772
rect 3710 848 3714 852
rect 3734 818 3738 822
rect 3782 1038 3786 1042
rect 3758 1008 3762 1012
rect 3750 948 3754 952
rect 3766 958 3770 962
rect 3862 1128 3866 1132
rect 3814 1118 3818 1122
rect 3838 1108 3842 1112
rect 3918 1198 3922 1202
rect 3918 1158 3922 1162
rect 3966 1358 3970 1362
rect 3950 1328 3954 1332
rect 3974 1328 3978 1332
rect 3942 1298 3946 1302
rect 3998 1318 4002 1322
rect 3974 1288 3978 1292
rect 3990 1218 3994 1222
rect 3942 1198 3946 1202
rect 3982 1158 3986 1162
rect 3894 1148 3898 1152
rect 3934 1148 3938 1152
rect 3878 1128 3882 1132
rect 3902 1128 3906 1132
rect 3934 1128 3938 1132
rect 3886 1118 3890 1122
rect 3870 1088 3874 1092
rect 4022 1408 4026 1412
rect 4118 1678 4122 1682
rect 4078 1558 4082 1562
rect 4158 1998 4162 2002
rect 4206 2028 4210 2032
rect 4166 1968 4170 1972
rect 4190 1958 4194 1962
rect 4230 2128 4234 2132
rect 4358 2148 4362 2152
rect 4302 2138 4306 2142
rect 4366 2138 4370 2142
rect 4342 2108 4346 2112
rect 4366 2128 4370 2132
rect 4262 2098 4266 2102
rect 4358 2098 4362 2102
rect 4254 2078 4258 2082
rect 4238 2058 4242 2062
rect 4214 2008 4218 2012
rect 4286 1978 4290 1982
rect 4254 1968 4258 1972
rect 4222 1958 4226 1962
rect 4246 1958 4250 1962
rect 4198 1948 4202 1952
rect 4182 1928 4186 1932
rect 4270 1948 4274 1952
rect 4310 2058 4314 2062
rect 4350 1958 4354 1962
rect 4318 1928 4322 1932
rect 4350 1928 4354 1932
rect 4390 2088 4394 2092
rect 4382 2078 4386 2082
rect 4382 2048 4386 2052
rect 4374 1988 4378 1992
rect 4390 2028 4394 2032
rect 4382 1928 4386 1932
rect 4294 1918 4298 1922
rect 4278 1898 4282 1902
rect 4270 1878 4274 1882
rect 4166 1868 4170 1872
rect 4206 1868 4210 1872
rect 4142 1848 4146 1852
rect 4174 1848 4178 1852
rect 4150 1838 4154 1842
rect 4166 1838 4170 1842
rect 4142 1758 4146 1762
rect 4214 1848 4218 1852
rect 4222 1788 4226 1792
rect 4246 1788 4250 1792
rect 4206 1778 4210 1782
rect 4206 1758 4210 1762
rect 4214 1758 4218 1762
rect 4230 1748 4234 1752
rect 4342 1918 4346 1922
rect 4366 1898 4370 1902
rect 4326 1868 4330 1872
rect 4366 1868 4370 1872
rect 4310 1848 4314 1852
rect 4278 1828 4282 1832
rect 4318 1808 4322 1812
rect 4366 1798 4370 1802
rect 4326 1788 4330 1792
rect 4334 1788 4338 1792
rect 4286 1758 4290 1762
rect 4302 1758 4306 1762
rect 4294 1728 4298 1732
rect 4206 1688 4210 1692
rect 4190 1678 4194 1682
rect 4222 1708 4226 1712
rect 4230 1688 4234 1692
rect 4286 1718 4290 1722
rect 4286 1708 4290 1712
rect 4310 1708 4314 1712
rect 4294 1698 4298 1702
rect 4270 1668 4274 1672
rect 4318 1688 4322 1692
rect 4142 1648 4146 1652
rect 4150 1648 4154 1652
rect 4166 1638 4170 1642
rect 4182 1598 4186 1602
rect 4166 1588 4170 1592
rect 4126 1548 4130 1552
rect 4142 1548 4146 1552
rect 4086 1538 4090 1542
rect 4102 1528 4106 1532
rect 4094 1518 4098 1522
rect 4070 1498 4074 1502
rect 4094 1498 4098 1502
rect 4114 1503 4118 1507
rect 4121 1503 4125 1507
rect 4150 1528 4154 1532
rect 4174 1518 4178 1522
rect 4134 1498 4138 1502
rect 4102 1478 4106 1482
rect 4054 1468 4058 1472
rect 4062 1468 4066 1472
rect 4038 1408 4042 1412
rect 4158 1468 4162 1472
rect 4126 1448 4130 1452
rect 4134 1438 4138 1442
rect 4126 1388 4130 1392
rect 4046 1358 4050 1362
rect 4118 1358 4122 1362
rect 4054 1348 4058 1352
rect 4030 1338 4034 1342
rect 4038 1338 4042 1342
rect 4014 1318 4018 1322
rect 4006 1288 4010 1292
rect 4086 1338 4090 1342
rect 4054 1328 4058 1332
rect 4070 1328 4074 1332
rect 4046 1298 4050 1302
rect 4086 1288 4090 1292
rect 4070 1278 4074 1282
rect 4114 1303 4118 1307
rect 4121 1303 4125 1307
rect 4150 1418 4154 1422
rect 4166 1328 4170 1332
rect 4166 1288 4170 1292
rect 4142 1278 4146 1282
rect 4110 1238 4114 1242
rect 4094 1228 4098 1232
rect 4126 1228 4130 1232
rect 4038 1208 4042 1212
rect 4022 1158 4026 1162
rect 3838 1068 3842 1072
rect 3926 1068 3930 1072
rect 3854 1058 3858 1062
rect 3958 1058 3962 1062
rect 3790 1028 3794 1032
rect 3822 1018 3826 1022
rect 3798 978 3802 982
rect 3830 958 3834 962
rect 3806 948 3810 952
rect 3798 938 3802 942
rect 3822 938 3826 942
rect 3774 928 3778 932
rect 3782 908 3786 912
rect 3782 898 3786 902
rect 3758 888 3762 892
rect 3750 868 3754 872
rect 3758 858 3762 862
rect 3814 928 3818 932
rect 3806 898 3810 902
rect 3822 888 3826 892
rect 3838 878 3842 882
rect 3758 848 3762 852
rect 3774 848 3778 852
rect 3822 838 3826 842
rect 3798 818 3802 822
rect 3822 818 3826 822
rect 3782 808 3786 812
rect 3846 808 3850 812
rect 3766 778 3770 782
rect 3798 778 3802 782
rect 3830 758 3834 762
rect 3710 748 3714 752
rect 3726 748 3730 752
rect 3782 748 3786 752
rect 3582 658 3586 662
rect 3610 603 3614 607
rect 3617 603 3621 607
rect 3526 588 3530 592
rect 3542 588 3546 592
rect 3518 578 3522 582
rect 3590 578 3594 582
rect 3550 568 3554 572
rect 3526 548 3530 552
rect 3566 558 3570 562
rect 3582 548 3586 552
rect 3510 538 3514 542
rect 3622 568 3626 572
rect 3630 548 3634 552
rect 3574 518 3578 522
rect 3510 478 3514 482
rect 3494 458 3498 462
rect 3502 378 3506 382
rect 3454 368 3458 372
rect 3462 368 3466 372
rect 3486 368 3490 372
rect 3406 348 3410 352
rect 3454 338 3458 342
rect 3326 328 3330 332
rect 3238 318 3242 322
rect 3254 298 3258 302
rect 3326 298 3330 302
rect 3334 298 3338 302
rect 3246 278 3250 282
rect 3174 258 3178 262
rect 3110 248 3114 252
rect 3222 218 3226 222
rect 3166 208 3170 212
rect 3158 178 3162 182
rect 3142 158 3146 162
rect 3086 148 3090 152
rect 3098 103 3102 107
rect 3105 103 3109 107
rect 3110 88 3114 92
rect 3174 168 3178 172
rect 3198 168 3202 172
rect 3214 168 3218 172
rect 3206 158 3210 162
rect 3238 138 3242 142
rect 3198 108 3202 112
rect 3230 98 3234 102
rect 3230 88 3234 92
rect 3310 288 3314 292
rect 3318 278 3322 282
rect 3342 278 3346 282
rect 3310 268 3314 272
rect 3342 248 3346 252
rect 3286 218 3290 222
rect 3366 318 3370 322
rect 3438 318 3442 322
rect 3422 298 3426 302
rect 3358 288 3362 292
rect 3446 308 3450 312
rect 3430 288 3434 292
rect 3358 268 3362 272
rect 3350 158 3354 162
rect 3390 248 3394 252
rect 3478 348 3482 352
rect 3486 338 3490 342
rect 3414 228 3418 232
rect 3382 218 3386 222
rect 3526 418 3530 422
rect 3518 368 3522 372
rect 3550 438 3554 442
rect 3526 348 3530 352
rect 3542 348 3546 352
rect 3566 428 3570 432
rect 3582 508 3586 512
rect 3590 488 3594 492
rect 3622 508 3626 512
rect 3686 738 3690 742
rect 3718 738 3722 742
rect 3726 658 3730 662
rect 3678 648 3682 652
rect 3670 618 3674 622
rect 3654 518 3658 522
rect 3638 478 3642 482
rect 3742 708 3746 712
rect 3822 748 3826 752
rect 3838 748 3842 752
rect 3814 688 3818 692
rect 3798 678 3802 682
rect 3854 678 3858 682
rect 3846 668 3850 672
rect 3750 658 3754 662
rect 3774 658 3778 662
rect 3750 638 3754 642
rect 3742 618 3746 622
rect 3742 608 3746 612
rect 3782 578 3786 582
rect 3734 568 3738 572
rect 3758 568 3762 572
rect 3766 568 3770 572
rect 3790 568 3794 572
rect 3678 538 3682 542
rect 3790 538 3794 542
rect 3806 608 3810 612
rect 3814 588 3818 592
rect 3822 578 3826 582
rect 3830 578 3834 582
rect 3814 568 3818 572
rect 3870 898 3874 902
rect 3870 838 3874 842
rect 3990 1048 3994 1052
rect 3918 1038 3922 1042
rect 3902 998 3906 1002
rect 3918 988 3922 992
rect 3950 1008 3954 1012
rect 3942 988 3946 992
rect 3926 978 3930 982
rect 3990 998 3994 1002
rect 4014 1078 4018 1082
rect 4086 1188 4090 1192
rect 4094 1188 4098 1192
rect 4046 1158 4050 1162
rect 4102 1158 4106 1162
rect 4054 1138 4058 1142
rect 4070 1138 4074 1142
rect 4142 1178 4146 1182
rect 4142 1168 4146 1172
rect 4286 1638 4290 1642
rect 4278 1618 4282 1622
rect 4246 1598 4250 1602
rect 4246 1588 4250 1592
rect 4270 1588 4274 1592
rect 4230 1558 4234 1562
rect 4190 1478 4194 1482
rect 4286 1578 4290 1582
rect 4318 1578 4322 1582
rect 4310 1558 4314 1562
rect 4238 1538 4242 1542
rect 4286 1538 4290 1542
rect 4238 1498 4242 1502
rect 4286 1528 4290 1532
rect 4318 1498 4322 1502
rect 4246 1478 4250 1482
rect 4262 1478 4266 1482
rect 4350 1778 4354 1782
rect 4366 1658 4370 1662
rect 4358 1648 4362 1652
rect 4350 1588 4354 1592
rect 4494 2288 4498 2292
rect 4534 2318 4538 2322
rect 4606 2438 4610 2442
rect 4590 2428 4594 2432
rect 4634 2403 4638 2407
rect 4641 2403 4645 2407
rect 4598 2338 4602 2342
rect 4574 2288 4578 2292
rect 4622 2328 4626 2332
rect 4646 2318 4650 2322
rect 4686 2278 4690 2282
rect 4470 2258 4474 2262
rect 4478 2258 4482 2262
rect 4510 2258 4514 2262
rect 4430 2248 4434 2252
rect 4438 2248 4442 2252
rect 4462 2248 4466 2252
rect 4422 2208 4426 2212
rect 4414 2138 4418 2142
rect 4414 2088 4418 2092
rect 4406 2048 4410 2052
rect 4414 2028 4418 2032
rect 4582 2238 4586 2242
rect 4462 2228 4466 2232
rect 4502 2228 4506 2232
rect 4438 2168 4442 2172
rect 4446 2158 4450 2162
rect 4494 2158 4498 2162
rect 4526 2158 4530 2162
rect 4462 2148 4466 2152
rect 4486 2148 4490 2152
rect 4518 2148 4522 2152
rect 4430 2098 4434 2102
rect 4454 2088 4458 2092
rect 4438 2078 4442 2082
rect 4438 2058 4442 2062
rect 4446 2048 4450 2052
rect 4422 2008 4426 2012
rect 4470 2078 4474 2082
rect 4502 2128 4506 2132
rect 4534 2128 4538 2132
rect 4518 2108 4522 2112
rect 4630 2258 4634 2262
rect 4614 2228 4618 2232
rect 4646 2228 4650 2232
rect 4590 2138 4594 2142
rect 4634 2203 4638 2207
rect 4641 2203 4645 2207
rect 4622 2078 4626 2082
rect 4486 2068 4490 2072
rect 4566 2068 4570 2072
rect 4582 2068 4586 2072
rect 4478 2058 4482 2062
rect 4454 1998 4458 2002
rect 4470 1978 4474 1982
rect 4454 1968 4458 1972
rect 4470 1958 4474 1962
rect 4422 1948 4426 1952
rect 4438 1948 4442 1952
rect 4430 1928 4434 1932
rect 4398 1908 4402 1912
rect 4406 1908 4410 1912
rect 4390 1898 4394 1902
rect 4382 1808 4386 1812
rect 4382 1758 4386 1762
rect 4382 1698 4386 1702
rect 4462 1928 4466 1932
rect 4438 1898 4442 1902
rect 4494 2038 4498 2042
rect 4518 2038 4522 2042
rect 4502 1998 4506 2002
rect 4494 1948 4498 1952
rect 4518 1948 4522 1952
rect 4486 1898 4490 1902
rect 4478 1888 4482 1892
rect 4454 1868 4458 1872
rect 4486 1868 4490 1872
rect 4430 1848 4434 1852
rect 4454 1848 4458 1852
rect 4486 1848 4490 1852
rect 4406 1828 4410 1832
rect 4414 1748 4418 1752
rect 4390 1668 4394 1672
rect 4382 1638 4386 1642
rect 4390 1608 4394 1612
rect 4422 1728 4426 1732
rect 4414 1718 4418 1722
rect 4414 1688 4418 1692
rect 4422 1638 4426 1642
rect 4470 1768 4474 1772
rect 4438 1758 4442 1762
rect 4470 1758 4474 1762
rect 4502 1788 4506 1792
rect 4478 1748 4482 1752
rect 4494 1748 4498 1752
rect 4590 2058 4594 2062
rect 4606 2048 4610 2052
rect 4774 2968 4778 2972
rect 4862 3248 4866 3252
rect 4918 3438 4922 3442
rect 4934 3378 4938 3382
rect 4950 3378 4954 3382
rect 5022 4248 5026 4252
rect 5070 4238 5074 4242
rect 5054 4178 5058 4182
rect 5046 4158 5050 4162
rect 5086 4158 5090 4162
rect 5062 4148 5066 4152
rect 5030 4128 5034 4132
rect 5062 4098 5066 4102
rect 5030 4078 5034 4082
rect 5014 3978 5018 3982
rect 5014 3958 5018 3962
rect 5086 4148 5090 4152
rect 5118 4168 5122 4172
rect 5182 4148 5186 4152
rect 5174 4138 5178 4142
rect 5102 4088 5106 4092
rect 5086 4048 5090 4052
rect 5086 3978 5090 3982
rect 5046 3968 5050 3972
rect 5070 3948 5074 3952
rect 5054 3938 5058 3942
rect 5070 3938 5074 3942
rect 5022 3908 5026 3912
rect 5014 3868 5018 3872
rect 5014 3758 5018 3762
rect 5038 3758 5042 3762
rect 5038 3728 5042 3732
rect 5070 3928 5074 3932
rect 5078 3888 5082 3892
rect 5094 3958 5098 3962
rect 5110 3998 5114 4002
rect 5118 3958 5122 3962
rect 5142 3958 5146 3962
rect 5102 3938 5106 3942
rect 5094 3918 5098 3922
rect 5126 3948 5130 3952
rect 5174 3928 5178 3932
rect 5134 3918 5138 3922
rect 5102 3908 5106 3912
rect 5094 3868 5098 3872
rect 5086 3858 5090 3862
rect 5054 3838 5058 3842
rect 5078 3838 5082 3842
rect 5086 3828 5090 3832
rect 5070 3818 5074 3822
rect 5086 3768 5090 3772
rect 5150 3848 5154 3852
rect 5134 3768 5138 3772
rect 5126 3758 5130 3762
rect 5078 3748 5082 3752
rect 5102 3738 5106 3742
rect 5054 3688 5058 3692
rect 5190 3708 5194 3712
rect 5022 3668 5026 3672
rect 5046 3668 5050 3672
rect 5030 3658 5034 3662
rect 5086 3668 5090 3672
rect 5102 3668 5106 3672
rect 5150 3668 5154 3672
rect 5166 3668 5170 3672
rect 5062 3658 5066 3662
rect 5110 3658 5114 3662
rect 5078 3618 5082 3622
rect 5014 3558 5018 3562
rect 5054 3548 5058 3552
rect 5062 3488 5066 3492
rect 5030 3458 5034 3462
rect 5006 3448 5010 3452
rect 4910 3368 4914 3372
rect 4918 3358 4922 3362
rect 4934 3358 4938 3362
rect 4966 3358 4970 3362
rect 4950 3348 4954 3352
rect 4918 3318 4922 3322
rect 4926 3278 4930 3282
rect 4926 3258 4930 3262
rect 4886 3248 4890 3252
rect 4910 3248 4914 3252
rect 4934 3248 4938 3252
rect 4878 3238 4882 3242
rect 4886 3198 4890 3202
rect 4910 3188 4914 3192
rect 4918 3178 4922 3182
rect 4934 3168 4938 3172
rect 4894 3148 4898 3152
rect 4870 3138 4874 3142
rect 4918 3138 4922 3142
rect 4862 3118 4866 3122
rect 4854 3078 4858 3082
rect 4870 3088 4874 3092
rect 4886 3088 4890 3092
rect 4878 3078 4882 3082
rect 4870 3058 4874 3062
rect 4862 3048 4866 3052
rect 4862 3028 4866 3032
rect 4870 2968 4874 2972
rect 4822 2948 4826 2952
rect 4846 2948 4850 2952
rect 4838 2938 4842 2942
rect 4870 2928 4874 2932
rect 4750 2888 4754 2892
rect 4798 2888 4802 2892
rect 4734 2868 4738 2872
rect 4710 2858 4714 2862
rect 4726 2858 4730 2862
rect 4814 2868 4818 2872
rect 4822 2858 4826 2862
rect 4790 2838 4794 2842
rect 4742 2798 4746 2802
rect 4758 2798 4762 2802
rect 4798 2758 4802 2762
rect 4742 2748 4746 2752
rect 4734 2738 4738 2742
rect 4838 2828 4842 2832
rect 4846 2818 4850 2822
rect 4910 3108 4914 3112
rect 4958 3338 4962 3342
rect 4998 3368 5002 3372
rect 4998 3348 5002 3352
rect 4974 3288 4978 3292
rect 4966 3198 4970 3202
rect 4982 3168 4986 3172
rect 4974 3148 4978 3152
rect 5054 3348 5058 3352
rect 5046 3328 5050 3332
rect 5094 3538 5098 3542
rect 5110 3538 5114 3542
rect 5134 3618 5138 3622
rect 5150 3598 5154 3602
rect 5158 3538 5162 3542
rect 5150 3528 5154 3532
rect 5166 3528 5170 3532
rect 5078 3518 5082 3522
rect 5086 3468 5090 3472
rect 5126 3498 5130 3502
rect 5118 3488 5122 3492
rect 5134 3468 5138 3472
rect 5150 3498 5154 3502
rect 5158 3478 5162 3482
rect 5150 3468 5154 3472
rect 5158 3448 5162 3452
rect 5174 3448 5178 3452
rect 5182 3438 5186 3442
rect 5166 3428 5170 3432
rect 5174 3388 5178 3392
rect 5166 3368 5170 3372
rect 5110 3358 5114 3362
rect 5142 3358 5146 3362
rect 5158 3358 5162 3362
rect 5102 3338 5106 3342
rect 5134 3338 5138 3342
rect 5070 3328 5074 3332
rect 5102 3328 5106 3332
rect 4998 3268 5002 3272
rect 5006 3258 5010 3262
rect 5094 3258 5098 3262
rect 5094 3198 5098 3202
rect 5062 3188 5066 3192
rect 5054 3158 5058 3162
rect 4998 3148 5002 3152
rect 5046 3148 5050 3152
rect 4998 3138 5002 3142
rect 5006 3138 5010 3142
rect 5030 3138 5034 3142
rect 4950 3118 4954 3122
rect 4990 3118 4994 3122
rect 4942 3088 4946 3092
rect 4894 2948 4898 2952
rect 4902 2928 4906 2932
rect 4886 2878 4890 2882
rect 5014 3118 5018 3122
rect 4990 3088 4994 3092
rect 5006 3068 5010 3072
rect 4974 3058 4978 3062
rect 4958 3048 4962 3052
rect 4926 3038 4930 3042
rect 4982 3008 4986 3012
rect 4990 2988 4994 2992
rect 4942 2968 4946 2972
rect 4966 2938 4970 2942
rect 4918 2878 4922 2882
rect 4886 2868 4890 2872
rect 4910 2868 4914 2872
rect 4822 2748 4826 2752
rect 4806 2728 4810 2732
rect 4838 2728 4842 2732
rect 4910 2808 4914 2812
rect 4902 2778 4906 2782
rect 4894 2758 4898 2762
rect 4886 2738 4890 2742
rect 4910 2728 4914 2732
rect 4862 2718 4866 2722
rect 4718 2708 4722 2712
rect 4750 2708 4754 2712
rect 4774 2678 4778 2682
rect 4870 2668 4874 2672
rect 4702 2558 4706 2562
rect 4710 2558 4714 2562
rect 4694 2258 4698 2262
rect 4790 2638 4794 2642
rect 4806 2618 4810 2622
rect 4830 2618 4834 2622
rect 4838 2618 4842 2622
rect 4750 2608 4754 2612
rect 4766 2578 4770 2582
rect 4782 2558 4786 2562
rect 4758 2548 4762 2552
rect 4806 2548 4810 2552
rect 4798 2538 4802 2542
rect 4814 2538 4818 2542
rect 4734 2528 4738 2532
rect 4782 2528 4786 2532
rect 4814 2528 4818 2532
rect 4846 2528 4850 2532
rect 4750 2498 4754 2502
rect 4734 2488 4738 2492
rect 4750 2448 4754 2452
rect 4758 2428 4762 2432
rect 4782 2488 4786 2492
rect 4838 2488 4842 2492
rect 4830 2478 4834 2482
rect 4782 2448 4786 2452
rect 4790 2438 4794 2442
rect 4766 2388 4770 2392
rect 4774 2378 4778 2382
rect 4782 2358 4786 2362
rect 4710 2338 4714 2342
rect 4750 2338 4754 2342
rect 4734 2328 4738 2332
rect 4734 2318 4738 2322
rect 4862 2478 4866 2482
rect 4846 2468 4850 2472
rect 4926 2798 4930 2802
rect 4926 2778 4930 2782
rect 4966 2918 4970 2922
rect 4950 2898 4954 2902
rect 5094 3178 5098 3182
rect 5078 3128 5082 3132
rect 5070 3078 5074 3082
rect 5046 3048 5050 3052
rect 5062 3048 5066 3052
rect 5070 3048 5074 3052
rect 5086 3048 5090 3052
rect 5070 2978 5074 2982
rect 5030 2958 5034 2962
rect 5054 2948 5058 2952
rect 5022 2898 5026 2902
rect 5022 2878 5026 2882
rect 5038 2878 5042 2882
rect 5054 2878 5058 2882
rect 5054 2868 5058 2872
rect 5094 2948 5098 2952
rect 4958 2848 4962 2852
rect 4966 2798 4970 2802
rect 4942 2778 4946 2782
rect 5022 2758 5026 2762
rect 5030 2758 5034 2762
rect 4958 2728 4962 2732
rect 4926 2718 4930 2722
rect 4958 2698 4962 2702
rect 4942 2678 4946 2682
rect 4966 2678 4970 2682
rect 4918 2618 4922 2622
rect 4990 2738 4994 2742
rect 5022 2678 5026 2682
rect 5086 2878 5090 2882
rect 5070 2848 5074 2852
rect 5070 2748 5074 2752
rect 5062 2708 5066 2712
rect 5086 2708 5090 2712
rect 5054 2668 5058 2672
rect 5078 2668 5082 2672
rect 4958 2658 4962 2662
rect 4974 2658 4978 2662
rect 4982 2658 4986 2662
rect 4998 2658 5002 2662
rect 5022 2658 5026 2662
rect 5038 2648 5042 2652
rect 5054 2648 5058 2652
rect 5062 2648 5066 2652
rect 4942 2628 4946 2632
rect 4878 2568 4882 2572
rect 4926 2568 4930 2572
rect 4934 2568 4938 2572
rect 4910 2558 4914 2562
rect 5062 2548 5066 2552
rect 4894 2528 4898 2532
rect 4878 2478 4882 2482
rect 4886 2478 4890 2482
rect 4862 2458 4866 2462
rect 4870 2458 4874 2462
rect 4846 2448 4850 2452
rect 4878 2438 4882 2442
rect 4798 2418 4802 2422
rect 4822 2418 4826 2422
rect 4854 2408 4858 2412
rect 4854 2378 4858 2382
rect 4806 2368 4810 2372
rect 4830 2358 4834 2362
rect 4966 2518 4970 2522
rect 4910 2478 4914 2482
rect 4982 2498 4986 2502
rect 5046 2498 5050 2502
rect 4998 2488 5002 2492
rect 4942 2448 4946 2452
rect 4902 2418 4906 2422
rect 4982 2398 4986 2402
rect 4934 2368 4938 2372
rect 4886 2358 4890 2362
rect 4902 2358 4906 2362
rect 4798 2348 4802 2352
rect 4854 2348 4858 2352
rect 4894 2348 4898 2352
rect 5142 3318 5146 3322
rect 5110 3198 5114 3202
rect 5158 3318 5162 3322
rect 5182 3258 5186 3262
rect 5182 3248 5186 3252
rect 5166 3188 5170 3192
rect 5150 3168 5154 3172
rect 5142 3148 5146 3152
rect 5126 3068 5130 3072
rect 5118 3048 5122 3052
rect 5126 2938 5130 2942
rect 5118 2868 5122 2872
rect 5118 2748 5122 2752
rect 5142 3098 5146 3102
rect 5158 3058 5162 3062
rect 5158 3048 5162 3052
rect 5174 3038 5178 3042
rect 5174 2968 5178 2972
rect 5150 2938 5154 2942
rect 5166 2938 5170 2942
rect 5166 2928 5170 2932
rect 5142 2908 5146 2912
rect 5142 2858 5146 2862
rect 5158 2818 5162 2822
rect 5118 2728 5122 2732
rect 5110 2688 5114 2692
rect 5102 2598 5106 2602
rect 5134 2688 5138 2692
rect 5182 2888 5186 2892
rect 5182 2768 5186 2772
rect 5182 2658 5186 2662
rect 5142 2648 5146 2652
rect 5166 2638 5170 2642
rect 5142 2618 5146 2622
rect 5126 2588 5130 2592
rect 5118 2578 5122 2582
rect 5102 2568 5106 2572
rect 5174 2568 5178 2572
rect 5094 2528 5098 2532
rect 5110 2558 5114 2562
rect 5158 2558 5162 2562
rect 5110 2548 5114 2552
rect 5126 2548 5130 2552
rect 5150 2538 5154 2542
rect 5134 2528 5138 2532
rect 5150 2518 5154 2522
rect 5150 2508 5154 2512
rect 5142 2488 5146 2492
rect 5118 2478 5122 2482
rect 5174 2498 5178 2502
rect 5182 2498 5186 2502
rect 5174 2468 5178 2472
rect 5118 2458 5122 2462
rect 5142 2458 5146 2462
rect 5110 2438 5114 2442
rect 5038 2368 5042 2372
rect 5086 2368 5090 2372
rect 4990 2358 4994 2362
rect 4870 2338 4874 2342
rect 4910 2338 4914 2342
rect 4926 2338 4930 2342
rect 4822 2318 4826 2322
rect 4798 2308 4802 2312
rect 4790 2298 4794 2302
rect 4830 2278 4834 2282
rect 4774 2268 4778 2272
rect 4694 2248 4698 2252
rect 4686 2198 4690 2202
rect 4694 2178 4698 2182
rect 4726 2248 4730 2252
rect 4726 2208 4730 2212
rect 4766 2208 4770 2212
rect 4734 2168 4738 2172
rect 4758 2168 4762 2172
rect 4670 2148 4674 2152
rect 4654 2138 4658 2142
rect 4702 2118 4706 2122
rect 4822 2258 4826 2262
rect 4846 2258 4850 2262
rect 4854 2258 4858 2262
rect 4790 2238 4794 2242
rect 4798 2238 4802 2242
rect 4798 2228 4802 2232
rect 4790 2158 4794 2162
rect 4798 2148 4802 2152
rect 4750 2138 4754 2142
rect 4766 2138 4770 2142
rect 4790 2138 4794 2142
rect 4718 2128 4722 2132
rect 4718 2118 4722 2122
rect 4710 2088 4714 2092
rect 4662 2068 4666 2072
rect 4662 2038 4666 2042
rect 4702 2048 4706 2052
rect 4638 2028 4642 2032
rect 4662 2028 4666 2032
rect 4670 2028 4674 2032
rect 4678 2028 4682 2032
rect 4634 2003 4638 2007
rect 4641 2003 4645 2007
rect 4566 1988 4570 1992
rect 4582 1978 4586 1982
rect 4526 1918 4530 1922
rect 4542 1908 4546 1912
rect 4526 1878 4530 1882
rect 4518 1838 4522 1842
rect 4462 1698 4466 1702
rect 4510 1698 4514 1702
rect 4550 1868 4554 1872
rect 4534 1858 4538 1862
rect 4558 1818 4562 1822
rect 4574 1928 4578 1932
rect 4590 1968 4594 1972
rect 4598 1958 4602 1962
rect 4646 1958 4650 1962
rect 4638 1948 4642 1952
rect 4654 1938 4658 1942
rect 4614 1918 4618 1922
rect 4654 1888 4658 1892
rect 4622 1878 4626 1882
rect 4574 1848 4578 1852
rect 4574 1828 4578 1832
rect 4582 1818 4586 1822
rect 4566 1808 4570 1812
rect 4534 1758 4538 1762
rect 4574 1728 4578 1732
rect 4590 1768 4594 1772
rect 4598 1768 4602 1772
rect 4614 1758 4618 1762
rect 4606 1748 4610 1752
rect 4606 1728 4610 1732
rect 4566 1718 4570 1722
rect 4582 1718 4586 1722
rect 4478 1688 4482 1692
rect 4534 1688 4538 1692
rect 4614 1688 4618 1692
rect 4502 1678 4506 1682
rect 4510 1678 4514 1682
rect 4446 1668 4450 1672
rect 4454 1668 4458 1672
rect 4634 1803 4638 1807
rect 4641 1803 4645 1807
rect 4630 1778 4634 1782
rect 4638 1678 4642 1682
rect 4558 1668 4562 1672
rect 4606 1668 4610 1672
rect 4622 1668 4626 1672
rect 4638 1668 4642 1672
rect 4734 2088 4738 2092
rect 4774 2068 4778 2072
rect 4710 1958 4714 1962
rect 4694 1948 4698 1952
rect 4678 1938 4682 1942
rect 4694 1938 4698 1942
rect 4702 1928 4706 1932
rect 4830 2188 4834 2192
rect 4798 2058 4802 2062
rect 4814 2048 4818 2052
rect 4734 1968 4738 1972
rect 4790 1968 4794 1972
rect 4822 1968 4826 1972
rect 4774 1958 4778 1962
rect 4774 1948 4778 1952
rect 4806 1948 4810 1952
rect 4750 1928 4754 1932
rect 4726 1918 4730 1922
rect 4742 1878 4746 1882
rect 4678 1868 4682 1872
rect 4662 1798 4666 1802
rect 4494 1658 4498 1662
rect 4566 1658 4570 1662
rect 4582 1658 4586 1662
rect 4438 1648 4442 1652
rect 4430 1618 4434 1622
rect 4414 1578 4418 1582
rect 4342 1548 4346 1552
rect 4374 1548 4378 1552
rect 4334 1488 4338 1492
rect 4254 1468 4258 1472
rect 4326 1468 4330 1472
rect 4254 1408 4258 1412
rect 4230 1388 4234 1392
rect 4254 1388 4258 1392
rect 4190 1368 4194 1372
rect 4182 1348 4186 1352
rect 4198 1348 4202 1352
rect 4206 1338 4210 1342
rect 4254 1308 4258 1312
rect 4206 1288 4210 1292
rect 4222 1288 4226 1292
rect 4246 1288 4250 1292
rect 4238 1278 4242 1282
rect 4278 1338 4282 1342
rect 4270 1318 4274 1322
rect 4262 1298 4266 1302
rect 4278 1298 4282 1302
rect 4262 1248 4266 1252
rect 4262 1238 4266 1242
rect 4246 1218 4250 1222
rect 4230 1188 4234 1192
rect 4198 1178 4202 1182
rect 4174 1168 4178 1172
rect 4214 1168 4218 1172
rect 4150 1158 4154 1162
rect 4206 1148 4210 1152
rect 4094 1128 4098 1132
rect 4046 1118 4050 1122
rect 4038 1068 4042 1072
rect 4062 1068 4066 1072
rect 4046 1058 4050 1062
rect 4062 1048 4066 1052
rect 4086 1008 4090 1012
rect 3990 978 3994 982
rect 3886 958 3890 962
rect 3926 948 3930 952
rect 3934 938 3938 942
rect 3934 918 3938 922
rect 3926 888 3930 892
rect 3918 868 3922 872
rect 3878 758 3882 762
rect 3894 798 3898 802
rect 3886 708 3890 712
rect 3910 768 3914 772
rect 3902 688 3906 692
rect 3862 638 3866 642
rect 3934 858 3938 862
rect 3926 848 3930 852
rect 3950 908 3954 912
rect 3950 898 3954 902
rect 3974 958 3978 962
rect 3982 928 3986 932
rect 3966 888 3970 892
rect 3958 868 3962 872
rect 3950 858 3954 862
rect 3982 828 3986 832
rect 3998 968 4002 972
rect 4022 968 4026 972
rect 4006 958 4010 962
rect 4014 948 4018 952
rect 3998 828 4002 832
rect 3982 788 3986 792
rect 3942 768 3946 772
rect 4094 958 4098 962
rect 4038 948 4042 952
rect 4078 948 4082 952
rect 4054 938 4058 942
rect 4070 938 4074 942
rect 4022 928 4026 932
rect 4030 928 4034 932
rect 4086 908 4090 912
rect 4078 888 4082 892
rect 4054 878 4058 882
rect 4022 868 4026 872
rect 4030 858 4034 862
rect 4014 828 4018 832
rect 4006 778 4010 782
rect 4014 758 4018 762
rect 4062 768 4066 772
rect 3926 748 3930 752
rect 3958 748 3962 752
rect 4070 748 4074 752
rect 3934 738 3938 742
rect 3934 728 3938 732
rect 3958 728 3962 732
rect 3998 728 4002 732
rect 3918 668 3922 672
rect 3886 628 3890 632
rect 3862 598 3866 602
rect 3854 588 3858 592
rect 3846 578 3850 582
rect 3878 568 3882 572
rect 3806 538 3810 542
rect 3862 538 3866 542
rect 3782 508 3786 512
rect 3798 508 3802 512
rect 3678 478 3682 482
rect 3742 478 3746 482
rect 3630 458 3634 462
rect 3610 403 3614 407
rect 3617 403 3621 407
rect 3574 378 3578 382
rect 3550 338 3554 342
rect 3558 328 3562 332
rect 3654 468 3658 472
rect 3638 398 3642 402
rect 3654 398 3658 402
rect 3646 358 3650 362
rect 3590 318 3594 322
rect 3510 268 3514 272
rect 3630 288 3634 292
rect 3550 278 3554 282
rect 3598 278 3602 282
rect 3630 278 3634 282
rect 3534 238 3538 242
rect 3502 228 3506 232
rect 3526 218 3530 222
rect 3470 208 3474 212
rect 3374 198 3378 202
rect 3590 248 3594 252
rect 3558 228 3562 232
rect 3590 228 3594 232
rect 3438 188 3442 192
rect 3526 188 3530 192
rect 3414 158 3418 162
rect 3390 138 3394 142
rect 3366 118 3370 122
rect 3470 178 3474 182
rect 3494 178 3498 182
rect 3454 148 3458 152
rect 3518 168 3522 172
rect 3486 148 3490 152
rect 3502 148 3506 152
rect 3406 138 3410 142
rect 3454 138 3458 142
rect 3398 98 3402 102
rect 3262 88 3266 92
rect 3350 88 3354 92
rect 3318 78 3322 82
rect 3086 68 3090 72
rect 3198 68 3202 72
rect 3214 68 3218 72
rect 3246 68 3250 72
rect 3030 58 3034 62
rect 2878 48 2882 52
rect 3014 48 3018 52
rect 3046 48 3050 52
rect 3166 48 3170 52
rect 3038 38 3042 42
rect 3382 68 3386 72
rect 3222 58 3226 62
rect 3494 108 3498 112
rect 3438 98 3442 102
rect 3446 88 3450 92
rect 3478 88 3482 92
rect 3478 68 3482 72
rect 3510 98 3514 102
rect 3470 58 3474 62
rect 3494 58 3498 62
rect 3534 178 3538 182
rect 3630 238 3634 242
rect 3670 468 3674 472
rect 3734 468 3738 472
rect 3694 398 3698 402
rect 3686 368 3690 372
rect 3678 348 3682 352
rect 3726 348 3730 352
rect 3750 408 3754 412
rect 3670 338 3674 342
rect 3678 338 3682 342
rect 3734 338 3738 342
rect 3670 298 3674 302
rect 3710 298 3714 302
rect 3662 268 3666 272
rect 3694 268 3698 272
rect 3726 288 3730 292
rect 3718 278 3722 282
rect 3750 298 3754 302
rect 3742 278 3746 282
rect 3694 238 3698 242
rect 3638 228 3642 232
rect 3610 203 3614 207
rect 3617 203 3621 207
rect 3734 248 3738 252
rect 3726 218 3730 222
rect 3662 188 3666 192
rect 3710 188 3714 192
rect 3638 168 3642 172
rect 3710 178 3714 182
rect 3670 168 3674 172
rect 3598 138 3602 142
rect 3646 138 3650 142
rect 3590 128 3594 132
rect 3670 118 3674 122
rect 3662 108 3666 112
rect 3670 108 3674 112
rect 3638 88 3642 92
rect 3686 88 3690 92
rect 3654 78 3658 82
rect 3662 68 3666 72
rect 3670 68 3674 72
rect 3582 58 3586 62
rect 3814 518 3818 522
rect 3854 518 3858 522
rect 3822 508 3826 512
rect 3886 508 3890 512
rect 3902 578 3906 582
rect 3902 538 3906 542
rect 3878 498 3882 502
rect 3894 498 3898 502
rect 3846 478 3850 482
rect 3782 468 3786 472
rect 3774 458 3778 462
rect 3790 418 3794 422
rect 3790 388 3794 392
rect 3822 458 3826 462
rect 3870 459 3874 463
rect 3830 428 3834 432
rect 3862 428 3866 432
rect 3814 408 3818 412
rect 3806 388 3810 392
rect 3798 338 3802 342
rect 3758 288 3762 292
rect 3782 288 3786 292
rect 3758 258 3762 262
rect 3774 258 3778 262
rect 3758 248 3762 252
rect 3774 248 3778 252
rect 3782 238 3786 242
rect 3814 368 3818 372
rect 3838 368 3842 372
rect 3846 368 3850 372
rect 3886 388 3890 392
rect 3822 358 3826 362
rect 3830 348 3834 352
rect 3854 348 3858 352
rect 3814 338 3818 342
rect 3806 268 3810 272
rect 3790 148 3794 152
rect 3814 148 3818 152
rect 3878 338 3882 342
rect 3854 318 3858 322
rect 3838 308 3842 312
rect 3838 278 3842 282
rect 3846 258 3850 262
rect 3830 218 3834 222
rect 3974 718 3978 722
rect 3966 708 3970 712
rect 3942 688 3946 692
rect 3934 668 3938 672
rect 3950 668 3954 672
rect 3934 648 3938 652
rect 3926 538 3930 542
rect 3926 518 3930 522
rect 3926 498 3930 502
rect 3934 488 3938 492
rect 3918 368 3922 372
rect 3958 598 3962 602
rect 3982 648 3986 652
rect 4070 718 4074 722
rect 4046 698 4050 702
rect 4054 688 4058 692
rect 4078 678 4082 682
rect 4070 638 4074 642
rect 4114 1103 4118 1107
rect 4121 1103 4125 1107
rect 4134 1058 4138 1062
rect 4142 998 4146 1002
rect 4114 903 4118 907
rect 4121 903 4125 907
rect 4126 888 4130 892
rect 4126 858 4130 862
rect 4134 758 4138 762
rect 4102 728 4106 732
rect 4114 703 4118 707
rect 4121 703 4125 707
rect 4086 628 4090 632
rect 4094 628 4098 632
rect 4070 578 4074 582
rect 4102 558 4106 562
rect 4006 548 4010 552
rect 3982 488 3986 492
rect 3950 478 3954 482
rect 3974 478 3978 482
rect 3966 468 3970 472
rect 3982 438 3986 442
rect 3966 358 3970 362
rect 3918 338 3922 342
rect 3894 278 3898 282
rect 4046 548 4050 552
rect 4062 548 4066 552
rect 4086 538 4090 542
rect 4054 518 4058 522
rect 4030 508 4034 512
rect 4094 508 4098 512
rect 4114 503 4118 507
rect 4121 503 4125 507
rect 4046 478 4050 482
rect 4086 478 4090 482
rect 4038 468 4042 472
rect 4030 398 4034 402
rect 4030 348 4034 352
rect 4014 328 4018 332
rect 3950 308 3954 312
rect 3958 308 3962 312
rect 3998 308 4002 312
rect 3934 278 3938 282
rect 3902 268 3906 272
rect 3910 258 3914 262
rect 3950 258 3954 262
rect 3854 178 3858 182
rect 3862 168 3866 172
rect 3838 148 3842 152
rect 3726 138 3730 142
rect 3814 128 3818 132
rect 3774 98 3778 102
rect 3822 98 3826 102
rect 3710 58 3714 62
rect 3406 48 3410 52
rect 3422 48 3426 52
rect 3438 48 3442 52
rect 3486 48 3490 52
rect 3502 48 3506 52
rect 3598 48 3602 52
rect 3718 48 3722 52
rect 3854 58 3858 62
rect 3870 58 3874 62
rect 4166 1138 4170 1142
rect 4174 1078 4178 1082
rect 4206 1068 4210 1072
rect 4214 1058 4218 1062
rect 4190 1038 4194 1042
rect 4214 968 4218 972
rect 4158 948 4162 952
rect 4214 938 4218 942
rect 4190 918 4194 922
rect 4214 918 4218 922
rect 4254 1018 4258 1022
rect 4302 1448 4306 1452
rect 4326 1438 4330 1442
rect 4310 1428 4314 1432
rect 4302 1298 4306 1302
rect 4294 1288 4298 1292
rect 4350 1448 4354 1452
rect 4334 1418 4338 1422
rect 4342 1388 4346 1392
rect 4398 1538 4402 1542
rect 4390 1528 4394 1532
rect 4398 1498 4402 1502
rect 4390 1488 4394 1492
rect 4366 1468 4370 1472
rect 4406 1468 4410 1472
rect 4390 1448 4394 1452
rect 4390 1378 4394 1382
rect 4422 1378 4426 1382
rect 4358 1368 4362 1372
rect 4374 1288 4378 1292
rect 4390 1288 4394 1292
rect 4326 1278 4330 1282
rect 4358 1278 4362 1282
rect 4318 1228 4322 1232
rect 4310 1178 4314 1182
rect 4302 1158 4306 1162
rect 4406 1268 4410 1272
rect 4358 1258 4362 1262
rect 4382 1258 4386 1262
rect 4350 1248 4354 1252
rect 4342 1228 4346 1232
rect 4382 1198 4386 1202
rect 4366 1188 4370 1192
rect 4342 1168 4346 1172
rect 4350 1158 4354 1162
rect 4286 1128 4290 1132
rect 4310 1078 4314 1082
rect 4326 1078 4330 1082
rect 4414 1248 4418 1252
rect 4582 1648 4586 1652
rect 4598 1648 4602 1652
rect 4462 1628 4466 1632
rect 4534 1618 4538 1622
rect 4462 1558 4466 1562
rect 4526 1548 4530 1552
rect 4462 1488 4466 1492
rect 4502 1518 4506 1522
rect 4486 1478 4490 1482
rect 4550 1568 4554 1572
rect 4566 1548 4570 1552
rect 4566 1488 4570 1492
rect 4574 1468 4578 1472
rect 4542 1458 4546 1462
rect 4542 1428 4546 1432
rect 4510 1408 4514 1412
rect 4534 1408 4538 1412
rect 4446 1398 4450 1402
rect 4478 1388 4482 1392
rect 4470 1328 4474 1332
rect 4462 1318 4466 1322
rect 4438 1298 4442 1302
rect 4518 1378 4522 1382
rect 4518 1338 4522 1342
rect 4486 1328 4490 1332
rect 4510 1328 4514 1332
rect 4486 1298 4490 1302
rect 4470 1288 4474 1292
rect 4446 1248 4450 1252
rect 4422 1218 4426 1222
rect 4582 1318 4586 1322
rect 4654 1648 4658 1652
rect 4646 1638 4650 1642
rect 4634 1603 4638 1607
rect 4641 1603 4645 1607
rect 4606 1588 4610 1592
rect 4654 1588 4658 1592
rect 4614 1568 4618 1572
rect 4638 1558 4642 1562
rect 4622 1518 4626 1522
rect 4614 1478 4618 1482
rect 4634 1403 4638 1407
rect 4641 1403 4645 1407
rect 4710 1838 4714 1842
rect 4822 1938 4826 1942
rect 4782 1908 4786 1912
rect 4798 1898 4802 1902
rect 4782 1868 4786 1872
rect 4750 1848 4754 1852
rect 4750 1828 4754 1832
rect 4774 1808 4778 1812
rect 4774 1778 4778 1782
rect 4758 1768 4762 1772
rect 4854 2158 4858 2162
rect 4846 2138 4850 2142
rect 4886 2238 4890 2242
rect 4862 2128 4866 2132
rect 4918 2158 4922 2162
rect 4934 2278 4938 2282
rect 4950 2268 4954 2272
rect 4934 2258 4938 2262
rect 4966 2248 4970 2252
rect 4974 2218 4978 2222
rect 4966 2148 4970 2152
rect 4966 2138 4970 2142
rect 4950 2128 4954 2132
rect 4878 2088 4882 2092
rect 4918 2078 4922 2082
rect 5070 2358 5074 2362
rect 5054 2338 5058 2342
rect 5086 2338 5090 2342
rect 5102 2338 5106 2342
rect 5046 2328 5050 2332
rect 5086 2328 5090 2332
rect 5126 2448 5130 2452
rect 5142 2448 5146 2452
rect 5158 2448 5162 2452
rect 5118 2348 5122 2352
rect 5134 2358 5138 2362
rect 5126 2328 5130 2332
rect 5030 2308 5034 2312
rect 5022 2288 5026 2292
rect 5054 2288 5058 2292
rect 5006 2278 5010 2282
rect 5006 2248 5010 2252
rect 4998 2128 5002 2132
rect 4990 2108 4994 2112
rect 4982 2078 4986 2082
rect 4974 2068 4978 2072
rect 4894 2048 4898 2052
rect 4942 2048 4946 2052
rect 4950 2048 4954 2052
rect 4950 2028 4954 2032
rect 4934 2018 4938 2022
rect 4950 2018 4954 2022
rect 4894 1978 4898 1982
rect 4854 1958 4858 1962
rect 4878 1958 4882 1962
rect 4862 1948 4866 1952
rect 4854 1898 4858 1902
rect 4838 1878 4842 1882
rect 4958 1958 4962 1962
rect 4990 2068 4994 2072
rect 5030 2228 5034 2232
rect 5014 2168 5018 2172
rect 5022 2108 5026 2112
rect 5054 2118 5058 2122
rect 5070 2308 5074 2312
rect 5078 2298 5082 2302
rect 5094 2298 5098 2302
rect 5078 2288 5082 2292
rect 5086 2278 5090 2282
rect 5134 2318 5138 2322
rect 5110 2298 5114 2302
rect 5102 2288 5106 2292
rect 5126 2288 5130 2292
rect 5102 2278 5106 2282
rect 5110 2268 5114 2272
rect 5078 2148 5082 2152
rect 5062 2098 5066 2102
rect 5030 2078 5034 2082
rect 5014 2068 5018 2072
rect 5038 2068 5042 2072
rect 5070 2068 5074 2072
rect 5046 2058 5050 2062
rect 5062 2058 5066 2062
rect 5006 2018 5010 2022
rect 5022 2008 5026 2012
rect 5022 1978 5026 1982
rect 4958 1918 4962 1922
rect 4966 1908 4970 1912
rect 4974 1888 4978 1892
rect 4998 1918 5002 1922
rect 5006 1888 5010 1892
rect 5014 1868 5018 1872
rect 4814 1848 4818 1852
rect 4838 1848 4842 1852
rect 4846 1848 4850 1852
rect 4870 1848 4874 1852
rect 4822 1828 4826 1832
rect 4838 1828 4842 1832
rect 4806 1818 4810 1822
rect 4790 1748 4794 1752
rect 4718 1728 4722 1732
rect 4726 1728 4730 1732
rect 4710 1718 4714 1722
rect 4782 1718 4786 1722
rect 4702 1688 4706 1692
rect 4678 1678 4682 1682
rect 4670 1668 4674 1672
rect 4758 1708 4762 1712
rect 4766 1668 4770 1672
rect 4718 1658 4722 1662
rect 4734 1658 4738 1662
rect 4750 1658 4754 1662
rect 4830 1778 4834 1782
rect 4814 1758 4818 1762
rect 4822 1738 4826 1742
rect 4798 1708 4802 1712
rect 4806 1708 4810 1712
rect 4862 1768 4866 1772
rect 4846 1728 4850 1732
rect 4830 1718 4834 1722
rect 4798 1698 4802 1702
rect 4814 1698 4818 1702
rect 4766 1648 4770 1652
rect 4790 1648 4794 1652
rect 4686 1628 4690 1632
rect 4774 1628 4778 1632
rect 4734 1618 4738 1622
rect 4662 1558 4666 1562
rect 4678 1558 4682 1562
rect 4710 1558 4714 1562
rect 4678 1548 4682 1552
rect 4742 1538 4746 1542
rect 4694 1518 4698 1522
rect 4694 1488 4698 1492
rect 4678 1468 4682 1472
rect 4686 1458 4690 1462
rect 4710 1448 4714 1452
rect 4662 1438 4666 1442
rect 4686 1438 4690 1442
rect 4654 1398 4658 1402
rect 4670 1368 4674 1372
rect 4662 1338 4666 1342
rect 4606 1318 4610 1322
rect 4598 1308 4602 1312
rect 4582 1278 4586 1282
rect 4502 1258 4506 1262
rect 4534 1258 4538 1262
rect 4462 1188 4466 1192
rect 4470 1168 4474 1172
rect 4566 1258 4570 1262
rect 4590 1248 4594 1252
rect 4622 1248 4626 1252
rect 4662 1238 4666 1242
rect 4634 1203 4638 1207
rect 4641 1203 4645 1207
rect 4550 1188 4554 1192
rect 4646 1178 4650 1182
rect 4598 1168 4602 1172
rect 4486 1158 4490 1162
rect 4510 1158 4514 1162
rect 4518 1158 4522 1162
rect 4414 1148 4418 1152
rect 4422 1148 4426 1152
rect 4438 1148 4442 1152
rect 4462 1148 4466 1152
rect 4470 1148 4474 1152
rect 4478 1148 4482 1152
rect 4502 1148 4506 1152
rect 4526 1148 4530 1152
rect 4374 1138 4378 1142
rect 4414 1128 4418 1132
rect 4406 1118 4410 1122
rect 4398 1098 4402 1102
rect 4390 1088 4394 1092
rect 4358 1068 4362 1072
rect 4342 1048 4346 1052
rect 4422 1068 4426 1072
rect 4478 1138 4482 1142
rect 4454 1078 4458 1082
rect 4430 1058 4434 1062
rect 4390 988 4394 992
rect 4398 978 4402 982
rect 4454 978 4458 982
rect 4390 968 4394 972
rect 4326 958 4330 962
rect 4342 958 4346 962
rect 4414 958 4418 962
rect 4550 1128 4554 1132
rect 4518 1108 4522 1112
rect 4630 1158 4634 1162
rect 4766 1508 4770 1512
rect 4742 1498 4746 1502
rect 4726 1488 4730 1492
rect 4750 1478 4754 1482
rect 4734 1448 4738 1452
rect 4758 1448 4762 1452
rect 4766 1408 4770 1412
rect 4782 1548 4786 1552
rect 4806 1678 4810 1682
rect 4950 1848 4954 1852
rect 4910 1838 4914 1842
rect 4958 1828 4962 1832
rect 4886 1788 4890 1792
rect 4918 1778 4922 1782
rect 4950 1768 4954 1772
rect 4894 1758 4898 1762
rect 4926 1758 4930 1762
rect 5014 1748 5018 1752
rect 4910 1738 4914 1742
rect 4934 1738 4938 1742
rect 4966 1738 4970 1742
rect 4974 1728 4978 1732
rect 4918 1718 4922 1722
rect 4958 1718 4962 1722
rect 4950 1688 4954 1692
rect 5022 1708 5026 1712
rect 4958 1668 4962 1672
rect 4838 1658 4842 1662
rect 4846 1648 4850 1652
rect 4838 1638 4842 1642
rect 4806 1618 4810 1622
rect 4870 1598 4874 1602
rect 4894 1598 4898 1602
rect 4854 1588 4858 1592
rect 4814 1528 4818 1532
rect 4878 1578 4882 1582
rect 4926 1638 4930 1642
rect 4910 1608 4914 1612
rect 4902 1588 4906 1592
rect 4830 1548 4834 1552
rect 4846 1548 4850 1552
rect 4854 1548 4858 1552
rect 4894 1548 4898 1552
rect 4822 1518 4826 1522
rect 4846 1498 4850 1502
rect 4886 1508 4890 1512
rect 4862 1488 4866 1492
rect 4878 1488 4882 1492
rect 4942 1648 4946 1652
rect 4934 1558 4938 1562
rect 4982 1548 4986 1552
rect 4998 1548 5002 1552
rect 4974 1538 4978 1542
rect 4934 1508 4938 1512
rect 4926 1478 4930 1482
rect 4934 1478 4938 1482
rect 4942 1478 4946 1482
rect 4830 1468 4834 1472
rect 4862 1468 4866 1472
rect 4902 1468 4906 1472
rect 4782 1418 4786 1422
rect 4814 1448 4818 1452
rect 4846 1448 4850 1452
rect 4822 1438 4826 1442
rect 4814 1428 4818 1432
rect 4830 1428 4834 1432
rect 4798 1408 4802 1412
rect 4758 1398 4762 1402
rect 4734 1358 4738 1362
rect 4702 1338 4706 1342
rect 4702 1318 4706 1322
rect 4734 1308 4738 1312
rect 4710 1298 4714 1302
rect 4702 1278 4706 1282
rect 4750 1278 4754 1282
rect 4822 1348 4826 1352
rect 4806 1338 4810 1342
rect 4790 1318 4794 1322
rect 4718 1268 4722 1272
rect 4686 1258 4690 1262
rect 4702 1248 4706 1252
rect 4750 1248 4754 1252
rect 4790 1248 4794 1252
rect 4726 1228 4730 1232
rect 4670 1158 4674 1162
rect 4742 1188 4746 1192
rect 4710 1158 4714 1162
rect 4582 1148 4586 1152
rect 4630 1148 4634 1152
rect 4662 1148 4666 1152
rect 4702 1148 4706 1152
rect 4598 1138 4602 1142
rect 4694 1138 4698 1142
rect 4566 1078 4570 1082
rect 4590 1078 4594 1082
rect 4630 1078 4634 1082
rect 4662 1078 4666 1082
rect 4526 1068 4530 1072
rect 4510 1058 4514 1062
rect 4486 988 4490 992
rect 4278 947 4282 951
rect 4342 948 4346 952
rect 4350 948 4354 952
rect 4446 948 4450 952
rect 4462 948 4466 952
rect 4358 938 4362 942
rect 4382 938 4386 942
rect 4278 928 4282 932
rect 4318 928 4322 932
rect 4446 928 4450 932
rect 4478 928 4482 932
rect 4302 918 4306 922
rect 4374 918 4378 922
rect 4302 898 4306 902
rect 4230 878 4234 882
rect 4246 878 4250 882
rect 4350 888 4354 892
rect 4310 878 4314 882
rect 4182 858 4186 862
rect 4254 858 4258 862
rect 4310 858 4314 862
rect 4190 848 4194 852
rect 4254 838 4258 842
rect 4214 758 4218 762
rect 4294 818 4298 822
rect 4374 848 4378 852
rect 4374 788 4378 792
rect 4350 778 4354 782
rect 4238 748 4242 752
rect 4254 748 4258 752
rect 4206 728 4210 732
rect 4206 688 4210 692
rect 4270 728 4274 732
rect 4246 698 4250 702
rect 4222 678 4226 682
rect 4246 678 4250 682
rect 4214 658 4218 662
rect 4198 648 4202 652
rect 4206 648 4210 652
rect 4158 638 4162 642
rect 4182 638 4186 642
rect 4190 628 4194 632
rect 4278 628 4282 632
rect 4238 608 4242 612
rect 4270 588 4274 592
rect 4294 758 4298 762
rect 4334 758 4338 762
rect 4302 748 4306 752
rect 4294 708 4298 712
rect 4326 708 4330 712
rect 4318 698 4322 702
rect 4310 688 4314 692
rect 4414 908 4418 912
rect 4438 908 4442 912
rect 4406 868 4410 872
rect 4470 888 4474 892
rect 4446 878 4450 882
rect 4454 868 4458 872
rect 4510 948 4514 952
rect 4574 1058 4578 1062
rect 4598 1058 4602 1062
rect 4630 1058 4634 1062
rect 4574 1018 4578 1022
rect 4542 968 4546 972
rect 4526 918 4530 922
rect 4526 888 4530 892
rect 4494 878 4498 882
rect 4566 888 4570 892
rect 4558 868 4562 872
rect 4582 878 4586 882
rect 4550 858 4554 862
rect 4422 848 4426 852
rect 4470 848 4474 852
rect 4502 808 4506 812
rect 4590 848 4594 852
rect 4590 838 4594 842
rect 4438 778 4442 782
rect 4510 768 4514 772
rect 4398 758 4402 762
rect 4438 758 4442 762
rect 4358 748 4362 752
rect 4390 748 4394 752
rect 4374 728 4378 732
rect 4398 728 4402 732
rect 4350 678 4354 682
rect 4366 678 4370 682
rect 4414 718 4418 722
rect 4518 718 4522 722
rect 4422 708 4426 712
rect 4478 708 4482 712
rect 4502 708 4506 712
rect 4438 688 4442 692
rect 4462 688 4466 692
rect 4422 678 4426 682
rect 4390 668 4394 672
rect 4406 668 4410 672
rect 4190 578 4194 582
rect 4166 568 4170 572
rect 4158 508 4162 512
rect 4190 498 4194 502
rect 4230 548 4234 552
rect 4262 548 4266 552
rect 4214 538 4218 542
rect 4254 508 4258 512
rect 4230 498 4234 502
rect 4254 498 4258 502
rect 4182 478 4186 482
rect 4222 468 4226 472
rect 4166 448 4170 452
rect 4070 408 4074 412
rect 4078 368 4082 372
rect 4070 348 4074 352
rect 4062 338 4066 342
rect 4062 318 4066 322
rect 4238 488 4242 492
rect 4262 478 4266 482
rect 4254 468 4258 472
rect 4486 698 4490 702
rect 4542 688 4546 692
rect 4454 678 4458 682
rect 4430 668 4434 672
rect 4446 668 4450 672
rect 4406 658 4410 662
rect 4414 658 4418 662
rect 4382 638 4386 642
rect 4374 598 4378 602
rect 4470 648 4474 652
rect 4486 648 4490 652
rect 4534 648 4538 652
rect 4462 638 4466 642
rect 4390 568 4394 572
rect 4454 558 4458 562
rect 4390 538 4394 542
rect 4318 498 4322 502
rect 4278 488 4282 492
rect 4310 468 4314 472
rect 4374 488 4378 492
rect 4374 468 4378 472
rect 4230 438 4234 442
rect 4150 408 4154 412
rect 4182 408 4186 412
rect 4134 358 4138 362
rect 4166 368 4170 372
rect 4198 368 4202 372
rect 4206 358 4210 362
rect 4166 348 4170 352
rect 4190 348 4194 352
rect 4214 348 4218 352
rect 4102 318 4106 322
rect 4114 303 4118 307
rect 4121 303 4125 307
rect 4046 288 4050 292
rect 4014 268 4018 272
rect 4030 268 4034 272
rect 4046 268 4050 272
rect 4054 268 4058 272
rect 4126 268 4130 272
rect 3974 248 3978 252
rect 4110 258 4114 262
rect 4054 198 4058 202
rect 4094 198 4098 202
rect 4014 188 4018 192
rect 4062 188 4066 192
rect 3974 148 3978 152
rect 4046 148 4050 152
rect 3910 138 3914 142
rect 3950 138 3954 142
rect 3998 128 4002 132
rect 3982 108 3986 112
rect 3950 88 3954 92
rect 4014 98 4018 102
rect 4022 98 4026 102
rect 4030 98 4034 102
rect 4006 88 4010 92
rect 3982 78 3986 82
rect 3958 68 3962 72
rect 3990 68 3994 72
rect 3910 58 3914 62
rect 4014 68 4018 72
rect 4070 178 4074 182
rect 4142 188 4146 192
rect 4198 338 4202 342
rect 4262 428 4266 432
rect 4238 418 4242 422
rect 4230 318 4234 322
rect 4238 318 4242 322
rect 4182 278 4186 282
rect 4190 268 4194 272
rect 4174 248 4178 252
rect 4238 308 4242 312
rect 4358 438 4362 442
rect 4334 408 4338 412
rect 4270 398 4274 402
rect 4342 358 4346 362
rect 4350 348 4354 352
rect 4286 308 4290 312
rect 4302 308 4306 312
rect 4214 238 4218 242
rect 4238 238 4242 242
rect 4206 228 4210 232
rect 4230 228 4234 232
rect 4214 218 4218 222
rect 4142 168 4146 172
rect 4166 168 4170 172
rect 4198 168 4202 172
rect 4118 148 4122 152
rect 4174 158 4178 162
rect 4198 158 4202 162
rect 4278 258 4282 262
rect 4262 208 4266 212
rect 4254 178 4258 182
rect 4238 168 4242 172
rect 4254 168 4258 172
rect 4254 158 4258 162
rect 4326 158 4330 162
rect 4230 148 4234 152
rect 4110 138 4114 142
rect 4158 138 4162 142
rect 4214 138 4218 142
rect 4246 138 4250 142
rect 4078 128 4082 132
rect 4222 128 4226 132
rect 4230 128 4234 132
rect 4190 118 4194 122
rect 4114 103 4118 107
rect 4121 103 4125 107
rect 4070 98 4074 102
rect 4198 108 4202 112
rect 4062 88 4066 92
rect 4046 68 4050 72
rect 4358 308 4362 312
rect 4358 298 4362 302
rect 4398 518 4402 522
rect 4422 548 4426 552
rect 4414 538 4418 542
rect 4446 538 4450 542
rect 4430 528 4434 532
rect 4438 468 4442 472
rect 4454 468 4458 472
rect 4430 458 4434 462
rect 4446 458 4450 462
rect 4406 448 4410 452
rect 4422 448 4426 452
rect 4382 418 4386 422
rect 4414 438 4418 442
rect 4390 368 4394 372
rect 4406 368 4410 372
rect 4406 348 4410 352
rect 4430 408 4434 412
rect 4422 328 4426 332
rect 4406 308 4410 312
rect 4406 298 4410 302
rect 4350 288 4354 292
rect 4374 288 4378 292
rect 4366 278 4370 282
rect 4382 268 4386 272
rect 4478 548 4482 552
rect 4478 518 4482 522
rect 4470 488 4474 492
rect 4494 528 4498 532
rect 4590 748 4594 752
rect 4726 1108 4730 1112
rect 4718 1048 4722 1052
rect 4614 1038 4618 1042
rect 4654 1038 4658 1042
rect 4694 1038 4698 1042
rect 4710 1038 4714 1042
rect 4622 1008 4626 1012
rect 4614 908 4618 912
rect 4634 1003 4638 1007
rect 4641 1003 4645 1007
rect 4638 988 4642 992
rect 4678 1028 4682 1032
rect 4702 998 4706 1002
rect 4734 988 4738 992
rect 4790 1228 4794 1232
rect 4830 1338 4834 1342
rect 4918 1448 4922 1452
rect 4998 1508 5002 1512
rect 4950 1438 4954 1442
rect 4958 1428 4962 1432
rect 4942 1368 4946 1372
rect 4950 1358 4954 1362
rect 4990 1358 4994 1362
rect 4886 1348 4890 1352
rect 4902 1348 4906 1352
rect 4950 1338 4954 1342
rect 4870 1308 4874 1312
rect 4894 1308 4898 1312
rect 4878 1278 4882 1282
rect 4934 1268 4938 1272
rect 4814 1258 4818 1262
rect 4838 1228 4842 1232
rect 4806 1168 4810 1172
rect 4798 1138 4802 1142
rect 4774 1128 4778 1132
rect 4806 1078 4810 1082
rect 4758 1068 4762 1072
rect 4750 1038 4754 1042
rect 4718 958 4722 962
rect 4678 948 4682 952
rect 4726 948 4730 952
rect 4694 938 4698 942
rect 4718 938 4722 942
rect 4726 888 4730 892
rect 4702 878 4706 882
rect 4774 1028 4778 1032
rect 4814 1068 4818 1072
rect 4854 1218 4858 1222
rect 4982 1308 4986 1312
rect 4974 1278 4978 1282
rect 5046 1988 5050 1992
rect 5094 2078 5098 2082
rect 5086 2058 5090 2062
rect 5110 2078 5114 2082
rect 5118 2078 5122 2082
rect 5110 2058 5114 2062
rect 5150 2428 5154 2432
rect 5166 2418 5170 2422
rect 5150 2288 5154 2292
rect 5142 2248 5146 2252
rect 5134 2228 5138 2232
rect 5158 2178 5162 2182
rect 5134 2128 5138 2132
rect 5150 2118 5154 2122
rect 5166 2098 5170 2102
rect 5150 2068 5154 2072
rect 5086 2018 5090 2022
rect 5102 2018 5106 2022
rect 5078 1958 5082 1962
rect 5078 1908 5082 1912
rect 5126 1988 5130 1992
rect 5102 1878 5106 1882
rect 5054 1868 5058 1872
rect 5150 2038 5154 2042
rect 5150 1988 5154 1992
rect 5190 2258 5194 2262
rect 5182 2208 5186 2212
rect 5174 2088 5178 2092
rect 5182 2068 5186 2072
rect 5174 2048 5178 2052
rect 5182 2038 5186 2042
rect 5182 1978 5186 1982
rect 5166 1938 5170 1942
rect 5174 1928 5178 1932
rect 5142 1888 5146 1892
rect 5174 1908 5178 1912
rect 5118 1858 5122 1862
rect 5166 1858 5170 1862
rect 5102 1848 5106 1852
rect 5062 1808 5066 1812
rect 5078 1798 5082 1802
rect 5078 1758 5082 1762
rect 5102 1758 5106 1762
rect 5110 1738 5114 1742
rect 5134 1738 5138 1742
rect 5150 1738 5154 1742
rect 5110 1728 5114 1732
rect 5030 1698 5034 1702
rect 5054 1678 5058 1682
rect 5078 1678 5082 1682
rect 5070 1658 5074 1662
rect 5054 1648 5058 1652
rect 5062 1558 5066 1562
rect 5070 1558 5074 1562
rect 5070 1548 5074 1552
rect 5062 1538 5066 1542
rect 5086 1538 5090 1542
rect 5046 1528 5050 1532
rect 5070 1528 5074 1532
rect 5038 1518 5042 1522
rect 5022 1488 5026 1492
rect 5046 1488 5050 1492
rect 5054 1468 5058 1472
rect 5190 1968 5194 1972
rect 5182 1748 5186 1752
rect 5150 1708 5154 1712
rect 5150 1638 5154 1642
rect 5142 1548 5146 1552
rect 5134 1508 5138 1512
rect 5086 1488 5090 1492
rect 5062 1458 5066 1462
rect 5086 1458 5090 1462
rect 5134 1458 5138 1462
rect 5094 1448 5098 1452
rect 5022 1438 5026 1442
rect 5126 1438 5130 1442
rect 5086 1428 5090 1432
rect 5030 1378 5034 1382
rect 5006 1358 5010 1362
rect 5062 1358 5066 1362
rect 5038 1348 5042 1352
rect 5134 1348 5138 1352
rect 4998 1338 5002 1342
rect 5022 1338 5026 1342
rect 5054 1338 5058 1342
rect 5014 1328 5018 1332
rect 5038 1328 5042 1332
rect 5014 1298 5018 1302
rect 5030 1268 5034 1272
rect 4990 1258 4994 1262
rect 5006 1258 5010 1262
rect 5014 1258 5018 1262
rect 5038 1258 5042 1262
rect 4950 1218 4954 1222
rect 4854 1148 4858 1152
rect 4878 1148 4882 1152
rect 4886 1148 4890 1152
rect 4918 1148 4922 1152
rect 4934 1148 4938 1152
rect 4966 1148 4970 1152
rect 4998 1148 5002 1152
rect 4886 1138 4890 1142
rect 4902 1138 4906 1142
rect 4926 1138 4930 1142
rect 4982 1138 4986 1142
rect 5006 1138 5010 1142
rect 4870 1118 4874 1122
rect 4894 1118 4898 1122
rect 4918 1118 4922 1122
rect 4830 1098 4834 1102
rect 4862 1088 4866 1092
rect 4878 1088 4882 1092
rect 4862 1078 4866 1082
rect 4902 1068 4906 1072
rect 4790 1008 4794 1012
rect 4798 988 4802 992
rect 4758 968 4762 972
rect 4782 968 4786 972
rect 4766 948 4770 952
rect 4774 938 4778 942
rect 4814 958 4818 962
rect 4798 948 4802 952
rect 4758 888 4762 892
rect 4654 868 4658 872
rect 4606 858 4610 862
rect 4638 858 4642 862
rect 4574 738 4578 742
rect 4598 738 4602 742
rect 4606 738 4610 742
rect 4558 698 4562 702
rect 4566 678 4570 682
rect 4582 668 4586 672
rect 4634 803 4638 807
rect 4641 803 4645 807
rect 4662 838 4666 842
rect 4734 858 4738 862
rect 4686 838 4690 842
rect 4710 838 4714 842
rect 4750 838 4754 842
rect 4758 828 4762 832
rect 4750 768 4754 772
rect 4822 918 4826 922
rect 4854 1058 4858 1062
rect 4878 1048 4882 1052
rect 4926 1048 4930 1052
rect 4870 968 4874 972
rect 4894 958 4898 962
rect 4910 958 4914 962
rect 4894 948 4898 952
rect 4926 948 4930 952
rect 4886 938 4890 942
rect 4870 908 4874 912
rect 4862 878 4866 882
rect 4814 868 4818 872
rect 4814 858 4818 862
rect 4806 828 4810 832
rect 4870 758 4874 762
rect 4766 748 4770 752
rect 4798 748 4802 752
rect 4806 748 4810 752
rect 4678 738 4682 742
rect 4734 738 4738 742
rect 4766 738 4770 742
rect 4862 738 4866 742
rect 4654 678 4658 682
rect 4622 668 4626 672
rect 4590 658 4594 662
rect 4598 658 4602 662
rect 4606 618 4610 622
rect 4646 618 4650 622
rect 4634 603 4638 607
rect 4641 603 4645 607
rect 4598 578 4602 582
rect 4694 708 4698 712
rect 4710 698 4714 702
rect 4758 698 4762 702
rect 4734 678 4738 682
rect 4790 728 4794 732
rect 4774 718 4778 722
rect 4806 718 4810 722
rect 4862 698 4866 702
rect 4782 688 4786 692
rect 4766 668 4770 672
rect 4862 668 4866 672
rect 4734 658 4738 662
rect 4758 658 4762 662
rect 4718 648 4722 652
rect 4726 648 4730 652
rect 4750 648 4754 652
rect 4702 638 4706 642
rect 4654 568 4658 572
rect 4630 558 4634 562
rect 4646 548 4650 552
rect 4606 538 4610 542
rect 4638 538 4642 542
rect 4558 528 4562 532
rect 4582 528 4586 532
rect 4654 528 4658 532
rect 4550 518 4554 522
rect 4510 478 4514 482
rect 4534 478 4538 482
rect 4590 508 4594 512
rect 4598 508 4602 512
rect 4622 508 4626 512
rect 4502 448 4506 452
rect 4494 438 4498 442
rect 4558 418 4562 422
rect 4526 368 4530 372
rect 4478 358 4482 362
rect 4510 358 4514 362
rect 4534 358 4538 362
rect 4718 498 4722 502
rect 4710 478 4714 482
rect 4590 458 4594 462
rect 4582 358 4586 362
rect 4518 348 4522 352
rect 4542 348 4546 352
rect 4470 288 4474 292
rect 4454 278 4458 282
rect 4446 268 4450 272
rect 4390 228 4394 232
rect 4526 338 4530 342
rect 4558 338 4562 342
rect 4566 328 4570 332
rect 4518 318 4522 322
rect 4518 298 4522 302
rect 4574 298 4578 302
rect 4634 403 4638 407
rect 4641 403 4645 407
rect 4622 398 4626 402
rect 4662 468 4666 472
rect 4686 468 4690 472
rect 4590 308 4594 312
rect 4590 298 4594 302
rect 4494 238 4498 242
rect 4462 218 4466 222
rect 4406 198 4410 202
rect 4422 198 4426 202
rect 4374 168 4378 172
rect 4366 158 4370 162
rect 4358 148 4362 152
rect 4382 148 4386 152
rect 4438 138 4442 142
rect 4358 128 4362 132
rect 4342 108 4346 112
rect 4230 98 4234 102
rect 4238 98 4242 102
rect 4198 78 4202 82
rect 4238 88 4242 92
rect 4342 88 4346 92
rect 4094 68 4098 72
rect 4190 68 4194 72
rect 4206 68 4210 72
rect 4222 68 4226 72
rect 3982 58 3986 62
rect 4022 58 4026 62
rect 3886 48 3890 52
rect 3966 48 3970 52
rect 3990 48 3994 52
rect 4014 48 4018 52
rect 4030 48 4034 52
rect 4302 78 4306 82
rect 4366 98 4370 102
rect 4382 98 4386 102
rect 4318 68 4322 72
rect 4366 68 4370 72
rect 4502 188 4506 192
rect 4614 308 4618 312
rect 4622 308 4626 312
rect 4654 288 4658 292
rect 4750 638 4754 642
rect 4798 648 4802 652
rect 4822 628 4826 632
rect 4758 578 4762 582
rect 4742 548 4746 552
rect 4782 538 4786 542
rect 4798 538 4802 542
rect 4814 538 4818 542
rect 4750 528 4754 532
rect 4758 488 4762 492
rect 4766 488 4770 492
rect 4734 468 4738 472
rect 4806 528 4810 532
rect 4910 788 4914 792
rect 4894 728 4898 732
rect 4886 698 4890 702
rect 4950 1128 4954 1132
rect 4942 1088 4946 1092
rect 4966 1078 4970 1082
rect 5014 1128 5018 1132
rect 4942 1068 4946 1072
rect 5062 1328 5066 1332
rect 5086 1288 5090 1292
rect 5174 1288 5178 1292
rect 5102 1278 5106 1282
rect 5166 1278 5170 1282
rect 5182 1278 5186 1282
rect 5062 1268 5066 1272
rect 5078 1258 5082 1262
rect 5054 1238 5058 1242
rect 5062 1238 5066 1242
rect 5118 1248 5122 1252
rect 5078 1148 5082 1152
rect 5054 1088 5058 1092
rect 5046 1068 5050 1072
rect 4990 1058 4994 1062
rect 5006 1058 5010 1062
rect 5030 1058 5034 1062
rect 5126 1028 5130 1032
rect 5174 1028 5178 1032
rect 4998 978 5002 982
rect 5030 958 5034 962
rect 5102 958 5106 962
rect 4942 948 4946 952
rect 4990 948 4994 952
rect 4982 898 4986 902
rect 4990 868 4994 872
rect 5150 948 5154 952
rect 5038 938 5042 942
rect 5134 938 5138 942
rect 5158 938 5162 942
rect 5014 928 5018 932
rect 5142 928 5146 932
rect 5166 928 5170 932
rect 5182 928 5186 932
rect 5126 918 5130 922
rect 5014 868 5018 872
rect 5078 848 5082 852
rect 4990 838 4994 842
rect 5046 788 5050 792
rect 4926 778 4930 782
rect 4950 778 4954 782
rect 4998 778 5002 782
rect 4958 758 4962 762
rect 4974 738 4978 742
rect 4918 708 4922 712
rect 4902 688 4906 692
rect 4910 688 4914 692
rect 5054 768 5058 772
rect 5062 768 5066 772
rect 5022 758 5026 762
rect 4990 668 4994 672
rect 5046 668 5050 672
rect 4926 658 4930 662
rect 4886 568 4890 572
rect 4910 558 4914 562
rect 5134 858 5138 862
rect 5118 798 5122 802
rect 5094 748 5098 752
rect 5070 738 5074 742
rect 5094 728 5098 732
rect 4998 658 5002 662
rect 5014 658 5018 662
rect 5086 668 5090 672
rect 5062 648 5066 652
rect 5030 588 5034 592
rect 4974 558 4978 562
rect 5062 568 5066 572
rect 5078 568 5082 572
rect 4846 548 4850 552
rect 4862 548 4866 552
rect 4878 548 4882 552
rect 4934 548 4938 552
rect 5046 548 5050 552
rect 4870 538 4874 542
rect 5046 538 5050 542
rect 4894 528 4898 532
rect 4918 528 4922 532
rect 4782 458 4786 462
rect 4790 458 4794 462
rect 4678 358 4682 362
rect 4670 308 4674 312
rect 4606 258 4610 262
rect 4662 258 4666 262
rect 4526 248 4530 252
rect 4590 248 4594 252
rect 4542 238 4546 242
rect 4550 238 4554 242
rect 4526 208 4530 212
rect 4510 148 4514 152
rect 4510 98 4514 102
rect 4518 98 4522 102
rect 4462 88 4466 92
rect 4510 88 4514 92
rect 4390 78 4394 82
rect 4406 78 4410 82
rect 4566 128 4570 132
rect 4518 68 4522 72
rect 4542 68 4546 72
rect 4414 58 4418 62
rect 4634 203 4638 207
rect 4641 203 4645 207
rect 4670 198 4674 202
rect 4646 168 4650 172
rect 4686 298 4690 302
rect 4742 358 4746 362
rect 4774 358 4778 362
rect 4822 498 4826 502
rect 4846 498 4850 502
rect 4950 488 4954 492
rect 5038 488 5042 492
rect 4878 468 4882 472
rect 5006 468 5010 472
rect 4830 458 4834 462
rect 4854 458 4858 462
rect 4894 458 4898 462
rect 4814 448 4818 452
rect 4806 428 4810 432
rect 4854 388 4858 392
rect 4862 378 4866 382
rect 4798 368 4802 372
rect 4942 448 4946 452
rect 4966 358 4970 362
rect 5006 358 5010 362
rect 4782 348 4786 352
rect 4790 348 4794 352
rect 4790 338 4794 342
rect 4750 328 4754 332
rect 4758 328 4762 332
rect 4734 318 4738 322
rect 4766 318 4770 322
rect 4702 288 4706 292
rect 4726 288 4730 292
rect 4718 268 4722 272
rect 4710 258 4714 262
rect 4774 268 4778 272
rect 4798 318 4802 322
rect 4806 298 4810 302
rect 4782 258 4786 262
rect 4774 248 4778 252
rect 4734 198 4738 202
rect 4726 178 4730 182
rect 4702 158 4706 162
rect 4606 148 4610 152
rect 4758 208 4762 212
rect 4750 188 4754 192
rect 4750 158 4754 162
rect 4750 148 4754 152
rect 4606 138 4610 142
rect 4598 108 4602 112
rect 4574 78 4578 82
rect 4582 68 4586 72
rect 4054 48 4058 52
rect 4110 48 4114 52
rect 4126 48 4130 52
rect 4230 48 4234 52
rect 4446 48 4450 52
rect 4558 48 4562 52
rect 3958 38 3962 42
rect 4062 38 4066 42
rect 4238 38 4242 42
rect 4366 38 4370 42
rect 4390 38 4394 42
rect 4406 38 4410 42
rect 4622 128 4626 132
rect 4702 108 4706 112
rect 4774 198 4778 202
rect 5014 348 5018 352
rect 4870 328 4874 332
rect 4830 318 4834 322
rect 4886 318 4890 322
rect 5078 538 5082 542
rect 5054 528 5058 532
rect 5182 858 5186 862
rect 5158 788 5162 792
rect 5174 798 5178 802
rect 5174 788 5178 792
rect 5166 768 5170 772
rect 5102 708 5106 712
rect 5126 708 5130 712
rect 5182 718 5186 722
rect 5190 718 5194 722
rect 5142 658 5146 662
rect 5134 548 5138 552
rect 5054 468 5058 472
rect 5070 468 5074 472
rect 5062 458 5066 462
rect 5062 368 5066 372
rect 5086 368 5090 372
rect 5054 348 5058 352
rect 5046 338 5050 342
rect 5062 338 5066 342
rect 5094 338 5098 342
rect 5182 418 5186 422
rect 4910 328 4914 332
rect 4894 288 4898 292
rect 4918 288 4922 292
rect 4942 268 4946 272
rect 4974 268 4978 272
rect 4862 258 4866 262
rect 4894 258 4898 262
rect 5062 298 5066 302
rect 5038 288 5042 292
rect 5126 298 5130 302
rect 5102 288 5106 292
rect 5110 288 5114 292
rect 5182 288 5186 292
rect 5110 278 5114 282
rect 5014 258 5018 262
rect 5046 258 5050 262
rect 5078 258 5082 262
rect 4854 248 4858 252
rect 4870 248 4874 252
rect 4830 218 4834 222
rect 4902 188 4906 192
rect 4790 178 4794 182
rect 4846 178 4850 182
rect 4870 178 4874 182
rect 4766 158 4770 162
rect 4814 168 4818 172
rect 4798 118 4802 122
rect 4806 118 4810 122
rect 4782 98 4786 102
rect 4838 158 4842 162
rect 4894 168 4898 172
rect 5022 218 5026 222
rect 4966 198 4970 202
rect 4998 178 5002 182
rect 4902 148 4906 152
rect 4894 128 4898 132
rect 4854 98 4858 102
rect 5054 158 5058 162
rect 5126 258 5130 262
rect 5110 208 5114 212
rect 5110 188 5114 192
rect 5166 158 5170 162
rect 5054 138 5058 142
rect 4830 88 4834 92
rect 4958 88 4962 92
rect 5014 88 5018 92
rect 4838 78 4842 82
rect 4950 78 4954 82
rect 4686 68 4690 72
rect 4902 68 4906 72
rect 5038 78 5042 82
rect 5126 68 5130 72
rect 5174 108 5178 112
rect 4758 58 4762 62
rect 4822 58 4826 62
rect 5134 58 5138 62
rect 4822 48 4826 52
rect 4854 48 4858 52
rect 2750 28 2754 32
rect 2774 28 2778 32
rect 3214 28 3218 32
rect 3790 28 3794 32
rect 4606 28 4610 32
rect 538 3 542 7
rect 545 3 549 7
rect 1562 3 1566 7
rect 1569 3 1573 7
rect 3254 8 3258 12
rect 2586 3 2590 7
rect 2593 3 2597 7
rect 3610 3 3614 7
rect 3617 3 3621 7
rect 4634 3 4638 7
rect 4641 3 4645 7
<< metal3 >>
rect 1048 4903 1050 4907
rect 1054 4903 1057 4907
rect 1062 4903 1064 4907
rect 2072 4903 2074 4907
rect 2078 4903 2081 4907
rect 2086 4903 2088 4907
rect 3096 4903 3098 4907
rect 3102 4903 3105 4907
rect 3110 4903 3112 4907
rect 4112 4903 4114 4907
rect 4118 4903 4121 4907
rect 4126 4903 4128 4907
rect 850 4888 958 4891
rect 962 4888 966 4891
rect 2314 4888 2398 4891
rect 3626 4888 3830 4891
rect 3994 4888 4078 4891
rect 5010 4888 5166 4891
rect 234 4878 286 4881
rect 290 4878 422 4881
rect 426 4878 454 4881
rect 458 4878 598 4881
rect 842 4878 870 4881
rect 1254 4881 1257 4888
rect 1194 4878 1257 4881
rect 1778 4878 1806 4881
rect 1810 4878 1838 4881
rect 1842 4878 1958 4881
rect 1962 4878 1974 4881
rect 2270 4881 2273 4888
rect 2178 4878 2273 4881
rect 2386 4878 2462 4881
rect 2602 4878 2894 4881
rect 3074 4878 3214 4881
rect 3218 4878 3342 4881
rect 3562 4878 3865 4881
rect 690 4868 710 4871
rect 714 4868 742 4871
rect 754 4868 990 4871
rect 994 4868 1070 4871
rect 1258 4868 1286 4871
rect 1502 4871 1505 4878
rect 3862 4872 3865 4878
rect 1502 4868 1550 4871
rect 1602 4868 1686 4871
rect 1762 4868 1790 4871
rect 1818 4868 1822 4871
rect 2138 4868 2254 4871
rect 2306 4868 2350 4871
rect 2434 4868 2438 4871
rect 2738 4868 3225 4871
rect 3354 4868 3678 4871
rect 3882 4868 4206 4871
rect 4238 4871 4241 4878
rect 4238 4868 4286 4871
rect 4370 4868 4510 4871
rect 4514 4868 4574 4871
rect 4702 4868 4806 4871
rect 4882 4868 4921 4871
rect 5042 4868 5062 4871
rect 182 4861 185 4868
rect 138 4858 185 4861
rect 214 4861 217 4868
rect 246 4861 249 4868
rect 582 4862 585 4868
rect 214 4858 249 4861
rect 258 4858 566 4861
rect 570 4858 574 4861
rect 706 4858 782 4861
rect 818 4858 846 4861
rect 882 4858 913 4861
rect 1050 4858 1150 4861
rect 1234 4858 1238 4861
rect 1338 4859 1358 4861
rect 1482 4859 1534 4861
rect 1338 4858 1361 4859
rect 1478 4858 1534 4859
rect 1554 4858 1678 4861
rect 1682 4858 1814 4861
rect 2094 4861 2097 4868
rect 2010 4858 2097 4861
rect 2122 4858 2190 4861
rect 2194 4858 2246 4861
rect 2250 4858 2342 4861
rect 2362 4859 2366 4861
rect 2358 4858 2366 4859
rect 2478 4861 2481 4868
rect 2686 4862 2689 4868
rect 3222 4862 3225 4868
rect 4702 4862 4705 4868
rect 4918 4862 4921 4868
rect 2442 4858 2481 4861
rect 2506 4858 2654 4861
rect 2714 4858 2782 4861
rect 2818 4858 2838 4861
rect 2962 4858 2982 4861
rect 3018 4858 3086 4861
rect 3194 4858 3198 4861
rect 3226 4858 3230 4861
rect 3290 4858 3358 4861
rect 3402 4858 3478 4861
rect 3794 4858 3854 4861
rect 3858 4858 3870 4861
rect 3878 4858 4182 4861
rect 4218 4858 4246 4861
rect 4250 4858 4254 4861
rect 4610 4858 4614 4861
rect 4774 4858 4822 4861
rect 4866 4858 4870 4861
rect 5034 4858 5046 4861
rect 910 4852 913 4858
rect 3878 4852 3881 4858
rect 4774 4852 4777 4858
rect 4934 4852 4937 4858
rect 5070 4852 5073 4858
rect 5102 4852 5105 4858
rect 194 4848 249 4851
rect 574 4848 582 4851
rect 586 4848 614 4851
rect 642 4848 766 4851
rect 770 4848 878 4851
rect 882 4848 894 4851
rect 1298 4848 2550 4851
rect 2686 4848 2705 4851
rect 3194 4848 3254 4851
rect 4050 4848 4606 4851
rect 4850 4848 4894 4851
rect 5222 4851 5226 4852
rect 5154 4848 5226 4851
rect 246 4842 249 4848
rect 2686 4842 2689 4848
rect 2702 4842 2705 4848
rect 698 4838 710 4841
rect 1242 4838 1270 4841
rect 1274 4838 1702 4841
rect 1738 4838 1790 4841
rect 2066 4838 2118 4841
rect 2254 4838 2270 4841
rect 2450 4838 2502 4841
rect 3046 4838 3054 4841
rect 3058 4838 3126 4841
rect 3154 4838 3225 4841
rect 3386 4838 3406 4841
rect 3410 4838 3790 4841
rect 3922 4838 4134 4841
rect 4146 4838 4678 4841
rect 4754 4838 4782 4841
rect 5010 4838 5102 4841
rect 2254 4832 2257 4838
rect 3222 4832 3225 4838
rect 82 4828 374 4831
rect 378 4828 750 4831
rect 834 4828 862 4831
rect 866 4828 1246 4831
rect 1298 4828 1302 4831
rect 1626 4828 1710 4831
rect 2674 4828 2742 4831
rect 3370 4828 3462 4831
rect 3586 4828 3694 4831
rect 3698 4828 3782 4831
rect 3786 4828 3910 4831
rect 4066 4828 4166 4831
rect 4170 4828 4318 4831
rect 4322 4828 4558 4831
rect 4690 4828 4950 4831
rect 162 4818 206 4821
rect 274 4818 382 4821
rect 506 4818 526 4821
rect 530 4818 710 4821
rect 1310 4821 1313 4828
rect 1074 4818 1422 4821
rect 1426 4818 1886 4821
rect 2058 4818 2086 4821
rect 2090 4818 2438 4821
rect 2522 4818 2534 4821
rect 2538 4818 2854 4821
rect 3226 4818 3374 4821
rect 3738 4818 4046 4821
rect 4226 4818 4358 4821
rect 4362 4818 4694 4821
rect 4818 4818 4934 4821
rect 4986 4818 5150 4821
rect 346 4808 366 4811
rect 1330 4808 1414 4811
rect 1658 4808 1670 4811
rect 1698 4808 1750 4811
rect 1770 4808 2078 4811
rect 2082 4808 2302 4811
rect 3770 4808 4166 4811
rect 4202 4808 4366 4811
rect 4906 4808 5014 4811
rect 5042 4808 5094 4811
rect 536 4803 538 4807
rect 542 4803 545 4807
rect 550 4803 552 4807
rect 1560 4803 1562 4807
rect 1566 4803 1569 4807
rect 1574 4803 1576 4807
rect 2584 4803 2586 4807
rect 2590 4803 2593 4807
rect 2598 4803 2600 4807
rect 3608 4803 3610 4807
rect 3614 4803 3617 4807
rect 3622 4803 3624 4807
rect 4632 4803 4634 4807
rect 4638 4803 4641 4807
rect 4646 4803 4648 4807
rect 578 4798 678 4801
rect 682 4798 782 4801
rect 2898 4798 3246 4801
rect 3338 4798 3446 4801
rect 3978 4798 4446 4801
rect 5022 4792 5025 4798
rect 370 4788 990 4791
rect 1530 4788 1814 4791
rect 2218 4788 2230 4791
rect 3098 4788 3406 4791
rect 3434 4788 3806 4791
rect 3834 4788 4206 4791
rect 4626 4788 4774 4791
rect 682 4778 726 4781
rect 1546 4778 1566 4781
rect 1954 4778 2086 4781
rect 2122 4778 2270 4781
rect 3210 4778 3414 4781
rect 3674 4778 4110 4781
rect 4138 4778 4190 4781
rect 4626 4778 4750 4781
rect 4754 4778 4902 4781
rect 106 4768 137 4771
rect 134 4762 137 4768
rect 822 4768 910 4771
rect 1506 4768 1518 4771
rect 1562 4768 1609 4771
rect 1730 4768 1950 4771
rect 1954 4768 2174 4771
rect 2198 4768 2206 4771
rect 2210 4768 2286 4771
rect 2290 4768 2318 4771
rect 2358 4768 2366 4771
rect 2370 4768 2430 4771
rect 2434 4768 2478 4771
rect 2502 4768 2694 4771
rect 2698 4768 2702 4771
rect 2718 4768 2750 4771
rect 3430 4771 3433 4778
rect 3242 4768 3433 4771
rect 3826 4768 4158 4771
rect 4258 4768 4830 4771
rect 4834 4768 4854 4771
rect 178 4758 310 4761
rect 686 4761 689 4768
rect 618 4758 689 4761
rect 806 4761 809 4768
rect 802 4758 809 4761
rect 822 4762 825 4768
rect 1606 4762 1609 4768
rect 1018 4758 1174 4761
rect 1178 4758 1182 4761
rect 1426 4758 1574 4761
rect 2042 4758 2102 4761
rect 2182 4761 2185 4768
rect 2502 4762 2505 4768
rect 2718 4762 2721 4768
rect 2182 4758 2198 4761
rect 2222 4758 2230 4761
rect 2234 4758 2278 4761
rect 2354 4758 2502 4761
rect 2522 4758 2566 4761
rect 2742 4758 2750 4761
rect 2754 4758 2814 4761
rect 3066 4758 3382 4761
rect 3582 4761 3585 4768
rect 3514 4758 3585 4761
rect 3810 4758 3846 4761
rect 3850 4758 3894 4761
rect 3978 4758 4070 4761
rect 4074 4758 4278 4761
rect 4282 4758 4446 4761
rect 4530 4758 4862 4761
rect 4866 4758 4918 4761
rect 5002 4758 5014 4761
rect 50 4748 121 4751
rect 162 4748 190 4751
rect 314 4748 678 4751
rect 706 4748 726 4751
rect 770 4748 793 4751
rect 854 4751 857 4758
rect 1358 4752 1361 4758
rect 802 4748 857 4751
rect 1186 4748 1190 4751
rect 1290 4748 1318 4751
rect 1322 4748 1350 4751
rect 1506 4748 1510 4751
rect 1602 4748 1622 4751
rect 1634 4748 1638 4751
rect 1682 4748 1686 4751
rect 1818 4748 1846 4751
rect 1890 4748 1998 4751
rect 2002 4748 2046 4751
rect 2154 4748 2246 4751
rect 2374 4748 2433 4751
rect 2450 4748 2510 4751
rect 2554 4748 2630 4751
rect 118 4742 121 4748
rect 758 4742 761 4748
rect 170 4738 182 4741
rect 250 4738 342 4741
rect 470 4738 486 4741
rect 650 4738 718 4741
rect 770 4738 774 4741
rect 790 4741 793 4748
rect 790 4738 822 4741
rect 1154 4738 1182 4741
rect 1274 4738 1286 4741
rect 1374 4741 1377 4748
rect 1622 4742 1625 4748
rect 1702 4742 1705 4748
rect 2374 4742 2377 4748
rect 2430 4742 2433 4748
rect 2758 4748 3238 4751
rect 3258 4748 3334 4751
rect 3410 4748 3438 4751
rect 3442 4748 3470 4751
rect 3474 4748 3606 4751
rect 3778 4748 3790 4751
rect 3866 4748 3942 4751
rect 4194 4748 4350 4751
rect 4546 4748 4622 4751
rect 4690 4748 4710 4751
rect 4842 4748 4918 4751
rect 4986 4748 5038 4751
rect 2758 4742 2761 4748
rect 1290 4738 1377 4741
rect 1402 4738 1606 4741
rect 1642 4738 1694 4741
rect 1706 4738 1734 4741
rect 1738 4738 1806 4741
rect 1882 4738 2054 4741
rect 2266 4738 2326 4741
rect 2330 4738 2334 4741
rect 2546 4738 2558 4741
rect 2562 4738 2654 4741
rect 2722 4738 2758 4741
rect 2842 4738 2977 4741
rect 3018 4738 3174 4741
rect 3178 4738 3206 4741
rect 3242 4738 3262 4741
rect 3418 4738 3446 4741
rect 3450 4738 3470 4741
rect 3714 4738 3766 4741
rect 3842 4738 3926 4741
rect 4106 4738 4113 4741
rect 4298 4738 4318 4741
rect 4538 4738 4574 4741
rect 470 4732 473 4738
rect 1206 4732 1209 4738
rect 138 4728 158 4731
rect 386 4728 470 4731
rect 530 4728 798 4731
rect 1090 4728 1126 4731
rect 1522 4728 1662 4731
rect 1666 4728 1766 4731
rect 1870 4731 1873 4738
rect 2230 4732 2233 4738
rect 2974 4732 2977 4738
rect 4110 4732 4113 4738
rect 1794 4728 1873 4731
rect 2026 4728 2158 4731
rect 2162 4728 2166 4731
rect 2530 4728 2686 4731
rect 2978 4728 3038 4731
rect 3042 4728 3110 4731
rect 3194 4728 3294 4731
rect 3370 4728 3486 4731
rect 3578 4728 3886 4731
rect 3890 4728 4110 4731
rect 4114 4728 4190 4731
rect 4466 4728 4510 4731
rect 4602 4728 4817 4731
rect 114 4718 262 4721
rect 298 4718 310 4721
rect 314 4718 350 4721
rect 358 4718 550 4721
rect 554 4718 758 4721
rect 1194 4718 1318 4721
rect 1330 4718 1598 4721
rect 1602 4718 1726 4721
rect 1858 4718 1902 4721
rect 2014 4721 2017 4728
rect 4814 4722 4817 4728
rect 2014 4718 2030 4721
rect 2106 4718 2134 4721
rect 2498 4718 2694 4721
rect 3002 4718 3118 4721
rect 3178 4718 3222 4721
rect 3554 4718 3558 4721
rect 3562 4718 3622 4721
rect 3658 4718 3750 4721
rect 3874 4718 3878 4721
rect 4002 4718 4030 4721
rect 4098 4718 4510 4721
rect 4514 4718 4582 4721
rect 4818 4718 4862 4721
rect 4954 4718 5030 4721
rect 5034 4718 5126 4721
rect 58 4708 102 4711
rect 178 4708 262 4711
rect 358 4711 361 4718
rect 314 4708 361 4711
rect 434 4708 566 4711
rect 578 4708 678 4711
rect 682 4708 686 4711
rect 714 4708 718 4711
rect 802 4708 846 4711
rect 1074 4708 1262 4711
rect 1546 4708 1862 4711
rect 1866 4708 1886 4711
rect 2002 4708 2022 4711
rect 2178 4708 2366 4711
rect 2494 4711 2497 4718
rect 2370 4708 2497 4711
rect 2906 4708 3030 4711
rect 3186 4708 3198 4711
rect 3642 4708 3838 4711
rect 4146 4708 4534 4711
rect 4618 4708 4638 4711
rect 1048 4703 1050 4707
rect 1054 4703 1057 4707
rect 1062 4703 1064 4707
rect 2072 4703 2074 4707
rect 2078 4703 2081 4707
rect 2086 4703 2088 4707
rect 3096 4703 3098 4707
rect 3102 4703 3105 4707
rect 3110 4703 3112 4707
rect 4112 4703 4114 4707
rect 4118 4703 4121 4707
rect 4126 4703 4128 4707
rect 210 4698 470 4701
rect 562 4698 750 4701
rect 1130 4698 1278 4701
rect 1306 4698 1318 4701
rect 1458 4698 1638 4701
rect 1818 4698 1974 4701
rect 2218 4698 2414 4701
rect 2418 4698 2726 4701
rect 2730 4698 2742 4701
rect 3146 4698 3182 4701
rect 3218 4698 3334 4701
rect 3386 4698 3390 4701
rect 3514 4698 3822 4701
rect 3834 4698 4006 4701
rect 4154 4698 4302 4701
rect 4306 4698 4374 4701
rect 4378 4698 4446 4701
rect 4554 4698 4686 4701
rect 4690 4698 4870 4701
rect 4874 4698 4966 4701
rect 94 4691 97 4698
rect 94 4688 134 4691
rect 186 4688 310 4691
rect 330 4688 478 4691
rect 482 4688 582 4691
rect 738 4688 798 4691
rect 970 4688 1161 4691
rect 1170 4688 1198 4691
rect 1250 4688 1433 4691
rect 1946 4688 2062 4691
rect 2354 4688 2390 4691
rect 2698 4688 2742 4691
rect 2866 4688 3014 4691
rect 3026 4688 3078 4691
rect 3082 4688 3150 4691
rect 3474 4688 3574 4691
rect 4082 4688 4158 4691
rect 4166 4688 4174 4691
rect 4178 4688 4246 4691
rect 4282 4688 4358 4691
rect 4370 4688 4422 4691
rect 4426 4688 4654 4691
rect 106 4678 318 4681
rect 346 4678 678 4681
rect 754 4678 806 4681
rect 810 4678 854 4681
rect 886 4681 889 4688
rect 858 4678 889 4681
rect 1158 4682 1161 4688
rect 1186 4678 1230 4681
rect 1238 4681 1241 4688
rect 1430 4682 1433 4688
rect 1238 4678 1302 4681
rect 1578 4678 1646 4681
rect 1714 4678 1894 4681
rect 1914 4678 2134 4681
rect 2238 4681 2241 4688
rect 2162 4678 2241 4681
rect 2298 4678 2422 4681
rect 2426 4678 3070 4681
rect 3230 4681 3233 4688
rect 3162 4678 3233 4681
rect 3250 4678 3366 4681
rect 3370 4678 3414 4681
rect 3426 4678 3534 4681
rect 3574 4681 3577 4688
rect 3574 4678 3614 4681
rect 3618 4678 3646 4681
rect 3650 4678 3830 4681
rect 3878 4681 3881 4688
rect 3878 4678 3910 4681
rect 4010 4678 4110 4681
rect 4114 4678 4134 4681
rect 4162 4678 4214 4681
rect 4218 4678 4318 4681
rect 4322 4678 4382 4681
rect 4418 4678 4526 4681
rect 4854 4678 4862 4681
rect 4866 4678 4942 4681
rect 1334 4672 1337 4678
rect 42 4668 126 4671
rect 194 4668 302 4671
rect 306 4668 334 4671
rect 338 4668 366 4671
rect 370 4668 430 4671
rect 450 4668 462 4671
rect 546 4668 566 4671
rect 590 4668 710 4671
rect 778 4668 878 4671
rect 1010 4668 1134 4671
rect 1138 4668 1150 4671
rect 1162 4668 1190 4671
rect 1194 4668 1254 4671
rect 1470 4671 1473 4678
rect 1378 4668 1473 4671
rect 1770 4668 1774 4671
rect 1898 4668 1958 4671
rect 2042 4668 2054 4671
rect 2242 4668 2262 4671
rect 2322 4668 2342 4671
rect 2346 4668 2374 4671
rect 2378 4668 2534 4671
rect 2562 4668 2630 4671
rect 2658 4668 2881 4671
rect 3154 4668 3174 4671
rect 3218 4668 3230 4671
rect 3242 4668 3374 4671
rect 3378 4668 3406 4671
rect 3578 4668 3582 4671
rect 3682 4668 3686 4671
rect 3802 4668 3894 4671
rect 3898 4668 3958 4671
rect 3978 4668 4169 4671
rect 4194 4668 4254 4671
rect 4266 4668 4326 4671
rect 4354 4668 4358 4671
rect 4374 4668 4406 4671
rect 4410 4668 4486 4671
rect 4578 4668 4630 4671
rect 4634 4668 4678 4671
rect 4682 4668 4702 4671
rect 4706 4668 4814 4671
rect 4990 4671 4993 4678
rect 4818 4668 4993 4671
rect 5050 4668 5054 4671
rect 5122 4668 5134 4671
rect 114 4658 142 4661
rect 146 4658 150 4661
rect 250 4658 286 4661
rect 290 4658 342 4661
rect 394 4658 422 4661
rect 426 4658 430 4661
rect 498 4658 502 4661
rect 590 4661 593 4668
rect 522 4658 593 4661
rect 602 4658 670 4661
rect 766 4661 769 4668
rect 746 4658 769 4661
rect 802 4658 814 4661
rect 934 4661 937 4668
rect 2782 4662 2785 4668
rect 2878 4662 2881 4668
rect 842 4658 937 4661
rect 1090 4658 1206 4661
rect 1218 4658 1222 4661
rect 1258 4658 1302 4661
rect 1314 4658 1318 4661
rect 1386 4658 1390 4661
rect 1438 4658 1454 4661
rect 1506 4658 1590 4661
rect 1714 4658 1782 4661
rect 1810 4658 1950 4661
rect 1954 4658 1998 4661
rect 2034 4658 2078 4661
rect 2082 4658 2230 4661
rect 2266 4658 2294 4661
rect 2298 4658 2326 4661
rect 2402 4658 2478 4661
rect 2554 4658 2694 4661
rect 2730 4658 2742 4661
rect 2986 4658 2990 4661
rect 3034 4658 3062 4661
rect 3170 4658 3190 4661
rect 3322 4658 3366 4661
rect 3402 4658 3473 4661
rect 3554 4658 3558 4661
rect 3726 4661 3729 4668
rect 4166 4662 4169 4668
rect 3674 4658 3729 4661
rect 3878 4658 3942 4661
rect 3986 4658 4006 4661
rect 4114 4658 4150 4661
rect 4170 4658 4174 4661
rect 4178 4658 4350 4661
rect 4374 4661 4377 4668
rect 4354 4658 4377 4661
rect 4386 4658 4438 4661
rect 4450 4658 4510 4661
rect 4514 4658 4550 4661
rect 4602 4658 4742 4661
rect 4746 4658 4790 4661
rect 4850 4658 4854 4661
rect 4874 4658 4886 4661
rect 4890 4658 5022 4661
rect 5074 4658 5126 4661
rect 106 4648 254 4651
rect 450 4648 510 4651
rect 850 4648 857 4651
rect 262 4641 265 4648
rect 854 4642 857 4648
rect 1014 4651 1017 4658
rect 882 4648 1017 4651
rect 1438 4651 1441 4658
rect 1622 4652 1625 4658
rect 3470 4652 3473 4658
rect 3646 4652 3649 4658
rect 3878 4652 3881 4658
rect 4054 4652 4057 4658
rect 1146 4648 1441 4651
rect 1450 4648 1582 4651
rect 1586 4648 1590 4651
rect 1802 4648 1817 4651
rect 194 4638 265 4641
rect 378 4638 526 4641
rect 658 4638 702 4641
rect 870 4641 873 4648
rect 870 4638 990 4641
rect 1134 4641 1137 4648
rect 1606 4642 1609 4648
rect 1814 4642 1817 4648
rect 1942 4648 1950 4651
rect 2122 4648 2718 4651
rect 2742 4648 2798 4651
rect 2986 4648 2998 4651
rect 3058 4648 3062 4651
rect 3086 4648 3110 4651
rect 3554 4648 3582 4651
rect 3674 4648 3798 4651
rect 3930 4648 3982 4651
rect 4058 4648 4494 4651
rect 4498 4648 4590 4651
rect 4642 4648 4678 4651
rect 4714 4648 4750 4651
rect 4770 4648 4774 4651
rect 4882 4648 4990 4651
rect 4994 4648 5030 4651
rect 5058 4648 5070 4651
rect 1134 4638 1230 4641
rect 1322 4638 1422 4641
rect 1434 4638 1446 4641
rect 1926 4641 1929 4648
rect 1842 4638 1929 4641
rect 1942 4642 1945 4648
rect 2742 4642 2745 4648
rect 3086 4642 3089 4648
rect 3190 4642 3193 4648
rect 4862 4642 4865 4648
rect 1978 4638 2214 4641
rect 2390 4638 2398 4641
rect 2402 4638 2422 4641
rect 2570 4638 2574 4641
rect 2770 4638 2854 4641
rect 2906 4638 2993 4641
rect 3298 4638 3302 4641
rect 3666 4638 3782 4641
rect 3818 4638 3862 4641
rect 3926 4638 3942 4641
rect 4050 4638 4086 4641
rect 4150 4638 4166 4641
rect 4210 4638 4286 4641
rect 4310 4638 4326 4641
rect 4346 4638 4358 4641
rect 4374 4638 4390 4641
rect 4586 4638 4590 4641
rect 4594 4638 4598 4641
rect 4610 4638 4654 4641
rect 4682 4638 4814 4641
rect 4866 4638 4886 4641
rect 2990 4632 2993 4638
rect 3926 4632 3929 4638
rect 4150 4632 4153 4638
rect 4310 4632 4313 4638
rect 4374 4632 4377 4638
rect 266 4628 486 4631
rect 522 4628 862 4631
rect 874 4628 1022 4631
rect 1026 4628 1310 4631
rect 1562 4628 1622 4631
rect 1778 4628 1918 4631
rect 1922 4628 1982 4631
rect 2018 4628 2262 4631
rect 2386 4628 2534 4631
rect 2538 4628 2582 4631
rect 2586 4628 2718 4631
rect 2722 4628 2758 4631
rect 3090 4628 3198 4631
rect 3202 4628 3222 4631
rect 3226 4628 3318 4631
rect 3354 4628 3870 4631
rect 4082 4628 4134 4631
rect 4426 4628 4518 4631
rect 4522 4628 4550 4631
rect 4562 4628 5046 4631
rect 5050 4628 5078 4631
rect 586 4618 654 4621
rect 658 4618 822 4621
rect 906 4618 942 4621
rect 1186 4618 1246 4621
rect 1250 4618 1502 4621
rect 1506 4618 1510 4621
rect 1514 4618 1558 4621
rect 1570 4618 1582 4621
rect 1770 4618 1798 4621
rect 2418 4618 2526 4621
rect 2530 4618 2542 4621
rect 2554 4618 3014 4621
rect 3018 4618 3486 4621
rect 3606 4618 3614 4621
rect 3618 4618 3646 4621
rect 3754 4618 3806 4621
rect 3810 4618 3910 4621
rect 3938 4618 4158 4621
rect 4210 4618 4246 4621
rect 4250 4618 4294 4621
rect 4586 4618 4598 4621
rect 4610 4618 4713 4621
rect 4786 4618 4998 4621
rect 5002 4618 5014 4621
rect 5082 4618 5142 4621
rect 4710 4612 4713 4618
rect 562 4608 662 4611
rect 666 4608 1142 4611
rect 1186 4608 1198 4611
rect 1586 4608 1694 4611
rect 1698 4608 1822 4611
rect 1826 4608 2102 4611
rect 2250 4608 2270 4611
rect 3978 4608 4526 4611
rect 4530 4608 4622 4611
rect 536 4603 538 4607
rect 542 4603 545 4607
rect 550 4603 552 4607
rect 1560 4603 1562 4607
rect 1566 4603 1569 4607
rect 1574 4603 1576 4607
rect 2584 4603 2586 4607
rect 2590 4603 2593 4607
rect 2598 4603 2600 4607
rect 3608 4603 3610 4607
rect 3614 4603 3617 4607
rect 3622 4603 3624 4607
rect 4632 4603 4634 4607
rect 4638 4603 4641 4607
rect 4646 4603 4648 4607
rect 642 4598 758 4601
rect 762 4598 1382 4601
rect 2042 4598 2542 4601
rect 2962 4598 3054 4601
rect 3874 4598 4094 4601
rect 4154 4598 4414 4601
rect 4818 4598 4838 4601
rect 2038 4592 2041 4598
rect 10 4588 46 4591
rect 50 4588 1230 4591
rect 1530 4588 1550 4591
rect 1554 4588 1590 4591
rect 1634 4588 1670 4591
rect 1674 4588 1790 4591
rect 1794 4588 2038 4591
rect 2162 4588 2726 4591
rect 2802 4588 3238 4591
rect 3690 4588 3734 4591
rect 3738 4588 3878 4591
rect 3882 4588 4110 4591
rect 4114 4588 4190 4591
rect 4194 4588 4246 4591
rect 4250 4588 4830 4591
rect 4834 4588 4862 4591
rect 290 4578 382 4581
rect 386 4578 558 4581
rect 658 4578 766 4581
rect 810 4578 1222 4581
rect 1418 4578 1950 4581
rect 2530 4578 2534 4581
rect 2698 4578 2702 4581
rect 2714 4578 3078 4581
rect 4066 4578 4102 4581
rect 4106 4578 4142 4581
rect 4282 4578 4326 4581
rect 4418 4578 4550 4581
rect 4570 4578 4678 4581
rect 278 4571 281 4578
rect 194 4568 281 4571
rect 322 4568 430 4571
rect 642 4568 662 4571
rect 714 4568 718 4571
rect 730 4568 766 4571
rect 794 4568 822 4571
rect 830 4568 838 4571
rect 842 4568 950 4571
rect 994 4568 1198 4571
rect 1218 4568 1246 4571
rect 1978 4568 2190 4571
rect 2226 4568 2254 4571
rect 2258 4568 2286 4571
rect 2390 4568 2590 4571
rect 2874 4568 3022 4571
rect 3054 4568 3062 4571
rect 3066 4568 3086 4571
rect 3410 4568 3814 4571
rect 4018 4568 4126 4571
rect 4282 4568 4382 4571
rect 4410 4568 4446 4571
rect 4618 4568 4630 4571
rect 4730 4568 4894 4571
rect 4898 4568 4926 4571
rect 274 4558 374 4561
rect 466 4558 686 4561
rect 690 4558 902 4561
rect 922 4558 958 4561
rect 1162 4558 1286 4561
rect 1802 4558 1814 4561
rect 1926 4561 1929 4568
rect 2390 4562 2393 4568
rect 1890 4558 1929 4561
rect 2090 4558 2142 4561
rect 2146 4558 2169 4561
rect 2282 4558 2318 4561
rect 2426 4558 2470 4561
rect 2702 4561 2705 4568
rect 2718 4561 2721 4568
rect 2702 4558 2721 4561
rect 2866 4558 2942 4561
rect 2978 4558 2982 4561
rect 3018 4558 3022 4561
rect 3034 4558 3134 4561
rect 3350 4561 3353 4568
rect 3350 4558 3406 4561
rect 3510 4558 3534 4561
rect 3570 4558 3686 4561
rect 4010 4558 4078 4561
rect 4518 4561 4521 4568
rect 4106 4558 4521 4561
rect 4546 4558 4566 4561
rect 4618 4558 4742 4561
rect 4746 4558 4798 4561
rect 4890 4558 5046 4561
rect 5050 4558 5094 4561
rect 5162 4558 5166 4561
rect 94 4551 97 4558
rect 94 4548 118 4551
rect 282 4548 302 4551
rect 314 4548 326 4551
rect 366 4548 417 4551
rect 490 4548 494 4551
rect 682 4548 702 4551
rect 710 4548 774 4551
rect 794 4548 846 4551
rect 970 4548 990 4551
rect 1242 4548 1246 4551
rect 1282 4548 1342 4551
rect 1362 4548 1374 4551
rect 1450 4548 1454 4551
rect 1498 4548 1502 4551
rect 1538 4548 1598 4551
rect 1798 4551 1801 4558
rect 2166 4552 2169 4558
rect 1730 4548 1801 4551
rect 1818 4548 1830 4551
rect 2050 4548 2126 4551
rect 2130 4548 2150 4551
rect 2390 4551 2393 4558
rect 3510 4552 3513 4558
rect 2274 4548 2393 4551
rect 2466 4548 2486 4551
rect 2522 4548 2526 4551
rect 2578 4548 2614 4551
rect 70 4541 73 4548
rect 166 4541 169 4548
rect 366 4542 369 4548
rect 414 4542 417 4548
rect 18 4538 169 4541
rect 426 4538 502 4541
rect 506 4538 518 4541
rect 710 4541 713 4548
rect 1638 4542 1641 4548
rect 2534 4542 2537 4548
rect 2698 4548 2790 4551
rect 2914 4548 2990 4551
rect 3002 4548 3022 4551
rect 3058 4548 3102 4551
rect 3154 4548 3230 4551
rect 3338 4548 3350 4551
rect 3490 4548 3494 4551
rect 3566 4551 3569 4558
rect 3522 4548 3569 4551
rect 3594 4548 3630 4551
rect 3722 4548 3758 4551
rect 3926 4551 3929 4558
rect 3818 4548 3905 4551
rect 3926 4548 3982 4551
rect 4010 4548 4030 4551
rect 4098 4548 4182 4551
rect 4218 4548 4310 4551
rect 4482 4548 4486 4551
rect 3902 4542 3905 4548
rect 4430 4542 4433 4548
rect 4494 4542 4497 4548
rect 4510 4542 4513 4548
rect 4802 4548 4846 4551
rect 4906 4548 4982 4551
rect 594 4538 713 4541
rect 754 4538 758 4541
rect 762 4538 806 4541
rect 842 4538 894 4541
rect 1298 4538 1366 4541
rect 1386 4538 1398 4541
rect 1450 4538 1614 4541
rect 1714 4538 1782 4541
rect 1978 4538 1982 4541
rect 2034 4538 2094 4541
rect 2186 4538 2190 4541
rect 2238 4538 2254 4541
rect 2362 4538 2374 4541
rect 2378 4538 2454 4541
rect 2674 4538 2678 4541
rect 2802 4538 2862 4541
rect 2986 4538 2990 4541
rect 3082 4538 3086 4541
rect 3146 4538 3158 4541
rect 3442 4538 3470 4541
rect 3530 4538 3534 4541
rect 3594 4538 3662 4541
rect 3670 4538 3678 4541
rect 4274 4538 4278 4541
rect 4298 4538 4398 4541
rect 4530 4538 4534 4541
rect 4546 4538 4558 4541
rect 4730 4538 4750 4541
rect 4822 4538 4966 4541
rect 5162 4538 5174 4541
rect 318 4532 321 4538
rect 734 4532 737 4538
rect 982 4532 985 4538
rect 1614 4532 1617 4538
rect 2238 4532 2241 4538
rect 2502 4532 2505 4538
rect 2966 4532 2969 4538
rect 3670 4532 3673 4538
rect 4062 4532 4065 4538
rect 4398 4532 4401 4538
rect 4822 4532 4825 4538
rect 338 4528 398 4531
rect 530 4528 646 4531
rect 650 4528 678 4531
rect 754 4528 790 4531
rect 858 4528 862 4531
rect 1242 4528 1574 4531
rect 1602 4528 1606 4531
rect 1714 4528 1718 4531
rect 1914 4528 1918 4531
rect 1970 4528 1982 4531
rect 2122 4528 2150 4531
rect 2210 4528 2214 4531
rect 2346 4528 2358 4531
rect 2530 4528 2686 4531
rect 2986 4528 3318 4531
rect 3322 4528 3534 4531
rect 3898 4528 3918 4531
rect 3922 4528 3982 4531
rect 4098 4528 4366 4531
rect 4458 4528 4558 4531
rect 4866 4528 4870 4531
rect 4930 4528 4942 4531
rect 4946 4528 4974 4531
rect 1926 4522 1929 4528
rect 3886 4522 3889 4528
rect 354 4518 470 4521
rect 474 4518 582 4521
rect 690 4518 750 4521
rect 762 4518 814 4521
rect 990 4518 998 4521
rect 1130 4518 1193 4521
rect 1218 4518 1230 4521
rect 1234 4518 1614 4521
rect 1618 4518 1622 4521
rect 1754 4518 1769 4521
rect 2234 4518 2454 4521
rect 2578 4518 2662 4521
rect 2914 4518 3374 4521
rect 3378 4518 3462 4521
rect 4018 4518 4214 4521
rect 4354 4518 4398 4521
rect 4410 4518 4486 4521
rect 4690 4518 4710 4521
rect 4862 4521 4865 4528
rect 4738 4518 4865 4521
rect 990 4512 993 4518
rect 1190 4512 1193 4518
rect 1766 4512 1769 4518
rect 826 4508 982 4511
rect 1346 4508 1398 4511
rect 1402 4508 1521 4511
rect 1554 4508 1630 4511
rect 1634 4508 1654 4511
rect 1770 4508 1774 4511
rect 1906 4508 2022 4511
rect 2194 4508 2270 4511
rect 2282 4508 2430 4511
rect 2450 4508 2566 4511
rect 2698 4508 2718 4511
rect 2826 4508 2942 4511
rect 3018 4508 3022 4511
rect 3026 4508 3086 4511
rect 3130 4508 3182 4511
rect 3386 4508 3398 4511
rect 3530 4508 3534 4511
rect 3546 4508 3550 4511
rect 3770 4508 3790 4511
rect 3826 4508 3934 4511
rect 3970 4508 4102 4511
rect 4162 4508 4590 4511
rect 4714 4508 5086 4511
rect 5090 4508 5190 4511
rect 1048 4503 1050 4507
rect 1054 4503 1057 4507
rect 1062 4503 1064 4507
rect 26 4498 94 4501
rect 770 4498 942 4501
rect 1314 4498 1438 4501
rect 1518 4501 1521 4508
rect 2072 4503 2074 4507
rect 2078 4503 2081 4507
rect 2086 4503 2088 4507
rect 3096 4503 3098 4507
rect 3102 4503 3105 4507
rect 3110 4503 3112 4507
rect 4112 4503 4114 4507
rect 4118 4503 4121 4507
rect 4126 4503 4128 4507
rect 1518 4498 1758 4501
rect 2250 4498 2254 4501
rect 2262 4498 2350 4501
rect 2402 4498 2462 4501
rect 2466 4498 2814 4501
rect 3458 4498 3606 4501
rect 3970 4498 3974 4501
rect 4202 4498 4462 4501
rect 4466 4498 4854 4501
rect 4866 4498 4878 4501
rect 5178 4498 5182 4501
rect 298 4488 318 4491
rect 322 4488 382 4491
rect 802 4488 1070 4491
rect 1074 4488 1158 4491
rect 1162 4488 1625 4491
rect 1650 4488 1758 4491
rect 1770 4488 2014 4491
rect 2262 4491 2265 4498
rect 2178 4488 2265 4491
rect 2482 4488 2518 4491
rect 2538 4488 2670 4491
rect 2730 4488 2742 4491
rect 2754 4488 2790 4491
rect 2794 4488 2838 4491
rect 2882 4488 3126 4491
rect 3298 4488 3518 4491
rect 3538 4488 3542 4491
rect 3770 4488 3782 4491
rect 3882 4488 3902 4491
rect 3954 4488 4065 4491
rect 4146 4488 4254 4491
rect 4262 4488 4454 4491
rect 4514 4488 4678 4491
rect 4682 4488 4694 4491
rect 4698 4488 4801 4491
rect 4858 4488 4918 4491
rect 4922 4488 5062 4491
rect 5066 4488 5078 4491
rect 1622 4482 1625 4488
rect 4062 4482 4065 4488
rect 106 4478 110 4481
rect 402 4478 422 4481
rect 642 4478 702 4481
rect 706 4478 758 4481
rect 786 4478 878 4481
rect 882 4478 894 4481
rect 1242 4478 1310 4481
rect 1314 4478 1342 4481
rect 1426 4478 1510 4481
rect 1626 4478 1878 4481
rect 1890 4478 2038 4481
rect 2138 4478 2310 4481
rect 2314 4478 2678 4481
rect 2738 4478 3150 4481
rect 3266 4478 3334 4481
rect 3410 4478 3486 4481
rect 3490 4478 4030 4481
rect 4262 4481 4265 4488
rect 4798 4482 4801 4488
rect 4122 4478 4265 4481
rect 4298 4478 4574 4481
rect 5042 4478 5062 4481
rect 5082 4478 5174 4481
rect 218 4468 326 4471
rect 354 4468 414 4471
rect 522 4468 614 4471
rect 782 4471 785 4478
rect 682 4468 785 4471
rect 810 4468 934 4471
rect 938 4468 1022 4471
rect 1102 4471 1105 4478
rect 1422 4472 1425 4478
rect 1026 4468 1105 4471
rect 1154 4468 1174 4471
rect 1338 4468 1358 4471
rect 1498 4468 1558 4471
rect 1594 4468 1598 4471
rect 1850 4468 1854 4471
rect 1922 4468 1926 4471
rect 2010 4468 2022 4471
rect 2242 4468 2246 4471
rect 2274 4468 2278 4471
rect 2306 4468 2414 4471
rect 2426 4468 2486 4471
rect 2490 4468 2534 4471
rect 2698 4468 2702 4471
rect 2722 4468 2742 4471
rect 2810 4468 2886 4471
rect 2978 4468 2982 4471
rect 3202 4468 3206 4471
rect 3250 4468 3278 4471
rect 3370 4468 3590 4471
rect 3802 4468 3806 4471
rect 3954 4468 3998 4471
rect 4294 4471 4297 4478
rect 4018 4468 4297 4471
rect 4442 4468 4446 4471
rect 4486 4468 4494 4471
rect 4498 4468 4582 4471
rect 4666 4468 4678 4471
rect 4682 4468 4814 4471
rect 4922 4468 4926 4471
rect 5022 4471 5025 4478
rect 5022 4468 5094 4471
rect 1190 4462 1193 4468
rect 114 4458 126 4461
rect 130 4458 166 4461
rect 250 4458 254 4461
rect 258 4458 278 4461
rect 282 4458 438 4461
rect 490 4458 702 4461
rect 714 4458 718 4461
rect 730 4458 734 4461
rect 738 4458 1094 4461
rect 1098 4458 1158 4461
rect 1222 4461 1225 4468
rect 1222 4458 1273 4461
rect 194 4448 265 4451
rect 446 4451 449 4458
rect 1270 4452 1273 4458
rect 1430 4458 1454 4461
rect 1506 4458 1510 4461
rect 1594 4458 1622 4461
rect 1678 4461 1681 4468
rect 1650 4458 1681 4461
rect 1778 4458 1790 4461
rect 1846 4458 1854 4461
rect 1998 4461 2001 4468
rect 1986 4458 2001 4461
rect 2030 4462 2033 4468
rect 2066 4458 2153 4461
rect 1430 4452 1433 4458
rect 1494 4452 1497 4458
rect 1622 4452 1625 4458
rect 1846 4452 1849 4458
rect 2150 4452 2153 4458
rect 2246 4458 2270 4461
rect 2362 4458 2366 4461
rect 2410 4458 2422 4461
rect 2426 4458 2518 4461
rect 2550 4461 2553 4468
rect 2522 4458 2553 4461
rect 2730 4458 2734 4461
rect 2774 4461 2777 4468
rect 2774 4458 2894 4461
rect 2950 4458 2998 4461
rect 3002 4458 3030 4461
rect 3218 4458 3230 4461
rect 3258 4458 3262 4461
rect 3458 4458 3542 4461
rect 3570 4458 3726 4461
rect 3782 4461 3785 4468
rect 3762 4458 3785 4461
rect 3866 4458 3878 4461
rect 3938 4458 3966 4461
rect 4026 4458 4049 4461
rect 4082 4458 4086 4461
rect 4170 4458 4278 4461
rect 4330 4458 4414 4461
rect 4418 4458 4430 4461
rect 4466 4458 4718 4461
rect 4754 4458 4758 4461
rect 4810 4458 4814 4461
rect 4842 4458 5046 4461
rect 5050 4458 5054 4461
rect 2246 4452 2249 4458
rect 2294 4452 2297 4458
rect 2950 4452 2953 4458
rect 3134 4452 3137 4458
rect 3902 4452 3905 4458
rect 4046 4452 4049 4458
rect 290 4448 449 4451
rect 594 4448 630 4451
rect 978 4448 998 4451
rect 1202 4448 1230 4451
rect 1234 4448 1238 4451
rect 1642 4448 1694 4451
rect 1786 4448 1830 4451
rect 1890 4448 1894 4451
rect 1914 4448 2030 4451
rect 2034 4448 2062 4451
rect 2386 4448 2510 4451
rect 2514 4448 2886 4451
rect 2978 4448 2982 4451
rect 3090 4448 3110 4451
rect 3238 4448 3246 4451
rect 3250 4448 3358 4451
rect 3506 4448 3558 4451
rect 3602 4448 3742 4451
rect 3746 4448 3862 4451
rect 4162 4448 4206 4451
rect 4282 4448 4294 4451
rect 4394 4448 4422 4451
rect 4610 4448 4670 4451
rect 4694 4448 4713 4451
rect 4818 4448 4846 4451
rect 4922 4448 4990 4451
rect 5054 4448 5110 4451
rect 262 4442 265 4448
rect 602 4438 614 4441
rect 698 4438 814 4441
rect 862 4441 865 4448
rect 902 4441 905 4448
rect 862 4438 905 4441
rect 934 4442 937 4448
rect 986 4438 990 4441
rect 1418 4438 1478 4441
rect 1562 4438 1854 4441
rect 1862 4438 1934 4441
rect 1962 4438 1966 4441
rect 2186 4438 2262 4441
rect 2330 4438 2334 4441
rect 2338 4438 2390 4441
rect 2478 4438 2614 4441
rect 2786 4438 2798 4441
rect 3058 4438 3174 4441
rect 3538 4438 3566 4441
rect 3590 4441 3593 4448
rect 4694 4442 4697 4448
rect 4710 4442 4713 4448
rect 5054 4442 5057 4448
rect 3590 4438 3662 4441
rect 3682 4438 3838 4441
rect 3890 4438 3910 4441
rect 3914 4438 4134 4441
rect 4162 4438 4326 4441
rect 4338 4438 4414 4441
rect 4506 4438 4582 4441
rect 4586 4438 4654 4441
rect 4834 4438 5038 4441
rect 810 4428 881 4431
rect 890 4428 1166 4431
rect 1862 4431 1865 4438
rect 1826 4428 1865 4431
rect 1882 4428 1950 4431
rect 2302 4431 2305 4438
rect 2026 4428 2305 4431
rect 2478 4432 2481 4438
rect 2498 4428 2694 4431
rect 2698 4428 2750 4431
rect 2950 4431 2953 4438
rect 2770 4428 2953 4431
rect 3546 4428 3806 4431
rect 3850 4428 4518 4431
rect 4522 4428 4814 4431
rect 4818 4428 4862 4431
rect 878 4422 881 4428
rect 58 4418 102 4421
rect 1018 4418 1558 4421
rect 1566 4421 1569 4428
rect 1566 4418 1582 4421
rect 1586 4418 1686 4421
rect 1714 4418 1734 4421
rect 1738 4418 1838 4421
rect 1874 4418 1942 4421
rect 1946 4418 2086 4421
rect 2170 4418 2526 4421
rect 2546 4418 2710 4421
rect 2762 4418 2790 4421
rect 2794 4418 2958 4421
rect 2962 4418 3214 4421
rect 3242 4418 3942 4421
rect 4050 4418 4494 4421
rect 4498 4418 4518 4421
rect 4538 4418 4902 4421
rect 4906 4418 4950 4421
rect 102 4412 105 4418
rect 578 4408 590 4411
rect 602 4408 1270 4411
rect 1274 4408 1334 4411
rect 1946 4408 1958 4411
rect 2754 4408 3126 4411
rect 3130 4408 3510 4411
rect 3826 4408 3926 4411
rect 3930 4408 3982 4411
rect 4010 4408 4054 4411
rect 4106 4408 4158 4411
rect 4266 4408 4270 4411
rect 4282 4408 4446 4411
rect 4538 4408 4542 4411
rect 4554 4408 4606 4411
rect 4738 4408 4782 4411
rect 4834 4408 4838 4411
rect 536 4403 538 4407
rect 542 4403 545 4407
rect 550 4403 552 4407
rect 1560 4403 1562 4407
rect 1566 4403 1569 4407
rect 1574 4403 1576 4407
rect 2584 4403 2586 4407
rect 2590 4403 2593 4407
rect 2598 4403 2600 4407
rect 3608 4403 3610 4407
rect 3614 4403 3617 4407
rect 3622 4403 3624 4407
rect 4632 4403 4634 4407
rect 4638 4403 4641 4407
rect 4646 4403 4648 4407
rect 626 4398 694 4401
rect 698 4398 758 4401
rect 1042 4398 1086 4401
rect 1090 4398 1094 4401
rect 1210 4398 1222 4401
rect 1802 4398 2246 4401
rect 2266 4398 2494 4401
rect 2826 4398 3062 4401
rect 3154 4398 3174 4401
rect 3194 4398 3206 4401
rect 3218 4398 3526 4401
rect 3746 4398 3854 4401
rect 4066 4398 4542 4401
rect 4706 4398 4750 4401
rect 4866 4398 4966 4401
rect 570 4388 838 4391
rect 874 4388 1038 4391
rect 1130 4388 1190 4391
rect 1218 4388 1222 4391
rect 1370 4388 1510 4391
rect 1954 4388 2094 4391
rect 2098 4388 2302 4391
rect 2666 4388 2806 4391
rect 2850 4388 3054 4391
rect 3378 4388 3406 4391
rect 3554 4388 3646 4391
rect 3650 4388 3686 4391
rect 3714 4388 4094 4391
rect 4102 4388 4110 4391
rect 4114 4388 4134 4391
rect 4154 4388 4230 4391
rect 4234 4388 4358 4391
rect 4522 4388 5017 4391
rect 5014 4382 5017 4388
rect 738 4378 798 4381
rect 802 4378 1030 4381
rect 1810 4378 1814 4381
rect 1826 4378 1926 4381
rect 1930 4378 1998 4381
rect 2002 4378 2062 4381
rect 2146 4378 2446 4381
rect 2514 4378 2534 4381
rect 2890 4378 3262 4381
rect 3626 4378 3750 4381
rect 3762 4378 3830 4381
rect 3834 4378 3854 4381
rect 3858 4378 3966 4381
rect 4034 4378 4222 4381
rect 4250 4378 4374 4381
rect 4514 4378 4758 4381
rect 4850 4378 4918 4381
rect 58 4368 94 4371
rect 98 4368 158 4371
rect 162 4368 286 4371
rect 962 4368 1022 4371
rect 1470 4371 1473 4378
rect 3494 4372 3497 4378
rect 1470 4368 1486 4371
rect 1602 4368 1790 4371
rect 1818 4368 1849 4371
rect 1906 4368 1910 4371
rect 2082 4368 2118 4371
rect 2138 4368 2190 4371
rect 2194 4368 2214 4371
rect 2370 4368 2390 4371
rect 2418 4368 2694 4371
rect 2706 4368 2710 4371
rect 2722 4368 2726 4371
rect 2794 4368 2814 4371
rect 2898 4368 2910 4371
rect 3026 4368 3134 4371
rect 3194 4368 3302 4371
rect 3442 4368 3462 4371
rect 3762 4368 3798 4371
rect 4034 4368 4206 4371
rect 4218 4368 4422 4371
rect 4434 4368 4926 4371
rect 4930 4368 4934 4371
rect 4938 4368 5078 4371
rect 10 4358 46 4361
rect 154 4358 182 4361
rect 298 4358 302 4361
rect 378 4358 398 4361
rect 574 4361 577 4368
rect 1846 4362 1849 4368
rect 474 4358 577 4361
rect 770 4358 822 4361
rect 994 4358 998 4361
rect 1226 4358 1286 4361
rect 1338 4358 1478 4361
rect 1482 4358 1582 4361
rect 1906 4358 2262 4361
rect 2282 4358 2286 4361
rect 2290 4358 2462 4361
rect 2482 4358 2486 4361
rect 2530 4358 2534 4361
rect 2546 4358 3142 4361
rect 3150 4361 3153 4368
rect 3150 4358 3270 4361
rect 3282 4358 3310 4361
rect 3346 4358 3438 4361
rect 3450 4358 3550 4361
rect 3562 4358 3966 4361
rect 3970 4358 3974 4361
rect 4070 4358 4078 4361
rect 4082 4358 4166 4361
rect 4322 4358 4382 4361
rect 4482 4358 4502 4361
rect 4514 4358 4598 4361
rect 4698 4358 4702 4361
rect 4738 4358 4766 4361
rect 4810 4358 4862 4361
rect 4874 4358 4881 4361
rect 4902 4358 4910 4361
rect 4914 4358 4974 4361
rect 5026 4358 5046 4361
rect 5050 4358 5182 4361
rect 86 4351 89 4358
rect 34 4348 89 4351
rect 242 4348 246 4351
rect 274 4348 278 4351
rect 398 4348 446 4351
rect 586 4348 598 4351
rect 698 4348 806 4351
rect 994 4348 1014 4351
rect 1174 4351 1177 4358
rect 1106 4348 1177 4351
rect 1234 4348 1265 4351
rect 398 4342 401 4348
rect 1262 4342 1265 4348
rect 1450 4348 1470 4351
rect 1634 4348 1638 4351
rect 1642 4348 1670 4351
rect 1750 4351 1753 4358
rect 1750 4348 1838 4351
rect 2122 4348 2158 4351
rect 2162 4348 2406 4351
rect 2450 4348 2470 4351
rect 2506 4348 2750 4351
rect 2778 4348 2782 4351
rect 2794 4348 2798 4351
rect 2818 4348 3006 4351
rect 3090 4348 3134 4351
rect 3146 4348 3150 4351
rect 3170 4348 3174 4351
rect 3418 4348 3470 4351
rect 3474 4348 3502 4351
rect 3554 4348 3670 4351
rect 3778 4348 3782 4351
rect 3898 4348 3958 4351
rect 4070 4351 4073 4358
rect 4310 4352 4313 4358
rect 3970 4348 4073 4351
rect 4082 4348 4094 4351
rect 4146 4348 4230 4351
rect 4330 4348 4334 4351
rect 4430 4351 4433 4358
rect 4378 4348 4433 4351
rect 4450 4348 4502 4351
rect 4594 4348 4766 4351
rect 4798 4351 4801 4358
rect 4878 4352 4881 4358
rect 4798 4348 4822 4351
rect 4898 4348 5030 4351
rect 5070 4348 5121 4351
rect 258 4338 262 4341
rect 334 4338 350 4341
rect 466 4338 614 4341
rect 618 4338 630 4341
rect 642 4338 774 4341
rect 842 4338 854 4341
rect 1002 4338 1006 4341
rect 1170 4338 1214 4341
rect 1366 4341 1369 4348
rect 1298 4338 1369 4341
rect 1394 4338 1486 4341
rect 1602 4338 1646 4341
rect 2054 4341 2057 4348
rect 1986 4338 2057 4341
rect 2066 4338 2145 4341
rect 334 4332 337 4338
rect 194 4328 238 4331
rect 434 4328 742 4331
rect 746 4328 870 4331
rect 962 4328 990 4331
rect 1122 4328 1142 4331
rect 1146 4328 1158 4331
rect 1226 4328 1342 4331
rect 1538 4328 1550 4331
rect 1554 4328 1630 4331
rect 1886 4331 1889 4338
rect 2142 4332 2145 4338
rect 2194 4338 2510 4341
rect 2514 4338 2542 4341
rect 2554 4338 2630 4341
rect 2802 4338 2830 4341
rect 2890 4338 3142 4341
rect 3162 4338 3190 4341
rect 3294 4341 3297 4348
rect 3294 4338 3366 4341
rect 3402 4338 3462 4341
rect 3482 4338 3486 4341
rect 3490 4338 3598 4341
rect 3778 4338 3782 4341
rect 3834 4338 3918 4341
rect 3938 4338 3942 4341
rect 3962 4338 3990 4341
rect 3994 4338 4014 4341
rect 4026 4338 4030 4341
rect 4058 4338 4262 4341
rect 4266 4338 4294 4341
rect 4358 4341 4361 4348
rect 5070 4342 5073 4348
rect 5118 4342 5121 4348
rect 4358 4338 4454 4341
rect 4698 4338 4758 4341
rect 4786 4338 4918 4341
rect 2174 4332 2177 4338
rect 2878 4332 2881 4338
rect 4558 4332 4561 4338
rect 1698 4328 1889 4331
rect 2450 4328 2454 4331
rect 2466 4328 2486 4331
rect 2570 4328 2646 4331
rect 2786 4328 2878 4331
rect 2922 4328 2966 4331
rect 2970 4328 3326 4331
rect 3426 4328 3486 4331
rect 3850 4328 3886 4331
rect 3962 4328 4158 4331
rect 4170 4328 4278 4331
rect 4290 4328 4350 4331
rect 4754 4328 4854 4331
rect 4874 4328 5030 4331
rect 26 4318 142 4321
rect 418 4318 422 4321
rect 858 4318 862 4321
rect 922 4318 966 4321
rect 970 4318 998 4321
rect 1002 4318 1110 4321
rect 1186 4318 1230 4321
rect 1458 4318 1694 4321
rect 2038 4321 2041 4328
rect 2038 4318 2174 4321
rect 2282 4318 2302 4321
rect 2346 4318 2502 4321
rect 2562 4318 2678 4321
rect 2682 4318 2686 4321
rect 2914 4318 2934 4321
rect 2942 4318 3198 4321
rect 3506 4318 3646 4321
rect 3898 4318 3974 4321
rect 3978 4318 4014 4321
rect 4018 4318 4126 4321
rect 4146 4318 4150 4321
rect 4234 4318 4342 4321
rect 4494 4321 4497 4328
rect 4354 4318 4497 4321
rect 4642 4318 4670 4321
rect 4674 4318 4726 4321
rect 4778 4318 5014 4321
rect 5018 4318 5086 4321
rect 586 4308 750 4311
rect 1098 4308 1246 4311
rect 1578 4308 1686 4311
rect 1690 4308 1910 4311
rect 1970 4308 1998 4311
rect 2426 4308 2718 4311
rect 2942 4311 2945 4318
rect 2738 4308 2945 4311
rect 3466 4308 3590 4311
rect 3890 4308 3926 4311
rect 4002 4308 4006 4311
rect 4138 4308 4278 4311
rect 4282 4308 4366 4311
rect 4370 4308 4502 4311
rect 4578 4308 4702 4311
rect 4706 4308 4790 4311
rect 4874 4308 4918 4311
rect 1048 4303 1050 4307
rect 1054 4303 1057 4307
rect 1062 4303 1064 4307
rect 2072 4303 2074 4307
rect 2078 4303 2081 4307
rect 2086 4303 2088 4307
rect 3096 4303 3098 4307
rect 3102 4303 3105 4307
rect 3110 4303 3112 4307
rect 4102 4302 4105 4308
rect 4112 4303 4114 4307
rect 4118 4303 4121 4307
rect 4126 4303 4128 4307
rect 666 4298 926 4301
rect 1234 4298 1374 4301
rect 1378 4298 1462 4301
rect 1474 4298 1646 4301
rect 1650 4298 1694 4301
rect 1770 4298 1846 4301
rect 1850 4298 1958 4301
rect 2194 4298 2246 4301
rect 2274 4298 2398 4301
rect 2410 4298 2606 4301
rect 2634 4298 2702 4301
rect 2706 4298 2830 4301
rect 2842 4298 2982 4301
rect 3330 4298 3334 4301
rect 3338 4298 3886 4301
rect 3914 4298 3934 4301
rect 3994 4298 4046 4301
rect 4138 4298 4150 4301
rect 4162 4298 4710 4301
rect 4770 4298 4822 4301
rect 578 4288 606 4291
rect 610 4288 694 4291
rect 770 4288 774 4291
rect 778 4288 1166 4291
rect 1346 4288 1406 4291
rect 1410 4288 1430 4291
rect 1586 4288 1622 4291
rect 1626 4288 1686 4291
rect 1754 4288 1798 4291
rect 1922 4288 2206 4291
rect 2218 4288 2222 4291
rect 2274 4288 2382 4291
rect 2666 4288 2686 4291
rect 2714 4288 2718 4291
rect 2850 4288 2854 4291
rect 2858 4288 3126 4291
rect 3142 4288 3310 4291
rect 3314 4288 3470 4291
rect 3514 4288 3526 4291
rect 3610 4288 3958 4291
rect 4050 4288 4070 4291
rect 4250 4288 4334 4291
rect 4482 4288 4566 4291
rect 4570 4288 4662 4291
rect 4818 4288 4958 4291
rect 146 4278 262 4281
rect 850 4278 894 4281
rect 906 4278 966 4281
rect 1170 4278 1190 4281
rect 1266 4278 1326 4281
rect 1618 4278 1782 4281
rect 2138 4278 2142 4281
rect 2154 4278 2166 4281
rect 2170 4278 2222 4281
rect 2354 4278 2366 4281
rect 2438 4281 2441 4288
rect 2434 4278 2441 4281
rect 3142 4281 3145 4288
rect 2498 4278 3145 4281
rect 3154 4278 3222 4281
rect 3242 4278 3310 4281
rect 3314 4278 3321 4281
rect 3426 4278 3454 4281
rect 3562 4278 3582 4281
rect 3794 4278 3806 4281
rect 3874 4278 4246 4281
rect 4258 4278 4526 4281
rect 4830 4278 4918 4281
rect 142 4271 145 4278
rect 74 4268 145 4271
rect 170 4268 246 4271
rect 290 4268 334 4271
rect 370 4268 422 4271
rect 426 4268 430 4271
rect 602 4268 638 4271
rect 726 4271 729 4278
rect 658 4268 729 4271
rect 798 4268 830 4271
rect 882 4268 902 4271
rect 938 4268 950 4271
rect 962 4268 966 4271
rect 1010 4268 1054 4271
rect 1058 4268 1070 4271
rect 1170 4268 1174 4271
rect 1314 4268 1326 4271
rect 1362 4268 1542 4271
rect 1706 4268 1726 4271
rect 2062 4271 2065 4278
rect 3782 4272 3785 4278
rect 3870 4272 3873 4278
rect 1962 4268 2065 4271
rect 2242 4268 2302 4271
rect 2306 4268 2350 4271
rect 2442 4268 2702 4271
rect 2746 4268 2838 4271
rect 3050 4268 3062 4271
rect 3106 4268 3150 4271
rect 3314 4268 3350 4271
rect 3354 4268 3470 4271
rect 3514 4268 3534 4271
rect 3562 4268 3574 4271
rect 3586 4268 3598 4271
rect 3722 4268 3758 4271
rect 3790 4268 3814 4271
rect 3850 4268 3862 4271
rect 3938 4268 3942 4271
rect 4026 4268 4038 4271
rect 4050 4268 4174 4271
rect 4182 4268 4230 4271
rect 4266 4268 4270 4271
rect 4290 4268 4318 4271
rect 4530 4268 4742 4271
rect 4798 4271 4801 4278
rect 4830 4272 4833 4278
rect 4798 4268 4814 4271
rect 4866 4268 4902 4271
rect 5066 4268 5126 4271
rect 5130 4268 5150 4271
rect 782 4262 785 4268
rect 798 4262 801 4268
rect 878 4262 881 4268
rect 66 4258 110 4261
rect 114 4258 366 4261
rect 378 4258 390 4261
rect 554 4258 558 4261
rect 710 4258 734 4261
rect 810 4258 814 4261
rect 934 4261 937 4268
rect 922 4258 937 4261
rect 998 4261 1001 4268
rect 998 4258 1014 4261
rect 1042 4259 1102 4261
rect 1042 4258 1105 4259
rect 1154 4258 1206 4261
rect 1210 4258 1217 4261
rect 1226 4258 1246 4261
rect 1290 4258 1318 4261
rect 1322 4258 1438 4261
rect 1590 4261 1593 4268
rect 1822 4262 1825 4268
rect 2150 4262 2153 4268
rect 2374 4262 2377 4268
rect 1506 4258 1593 4261
rect 1698 4258 1734 4261
rect 1890 4258 1966 4261
rect 1994 4258 2038 4261
rect 2202 4258 2278 4261
rect 2666 4258 2670 4261
rect 2714 4258 2726 4261
rect 2746 4258 2750 4261
rect 2922 4258 2926 4261
rect 2962 4258 2966 4261
rect 3146 4258 3150 4261
rect 3158 4261 3161 4268
rect 3158 4258 3182 4261
rect 3202 4258 3342 4261
rect 3434 4258 3478 4261
rect 3538 4258 3569 4261
rect 710 4252 713 4258
rect 290 4248 438 4251
rect 786 4248 854 4251
rect 874 4248 1006 4251
rect 1034 4248 1054 4251
rect 1058 4248 1166 4251
rect 1194 4248 1206 4251
rect 1214 4251 1217 4258
rect 1814 4252 1817 4258
rect 2182 4252 2185 4258
rect 2286 4252 2289 4258
rect 2310 4252 2313 4258
rect 2342 4252 2345 4258
rect 2382 4252 2385 4258
rect 3566 4252 3569 4258
rect 3602 4258 3654 4261
rect 3790 4261 3793 4268
rect 3878 4262 3881 4268
rect 3918 4262 3921 4268
rect 3754 4258 3793 4261
rect 3802 4258 3806 4261
rect 3866 4258 3870 4261
rect 4042 4258 4073 4261
rect 4182 4261 4185 4268
rect 4238 4262 4241 4268
rect 4090 4258 4185 4261
rect 4314 4258 4398 4261
rect 4494 4261 4497 4268
rect 4434 4258 4497 4261
rect 4506 4258 4558 4261
rect 4610 4258 4622 4261
rect 4674 4258 4678 4261
rect 4742 4261 4745 4268
rect 4742 4258 4798 4261
rect 4850 4258 4998 4261
rect 3598 4252 3601 4258
rect 4022 4252 4025 4258
rect 4070 4252 4073 4258
rect 1214 4248 1222 4251
rect 1314 4248 1382 4251
rect 1554 4248 1614 4251
rect 1686 4248 1694 4251
rect 1698 4248 1758 4251
rect 1842 4248 2110 4251
rect 2726 4248 2782 4251
rect 2918 4248 2990 4251
rect 3026 4248 3150 4251
rect 3330 4248 3342 4251
rect 3482 4248 3526 4251
rect 3634 4248 3638 4251
rect 3658 4248 3662 4251
rect 3746 4248 3766 4251
rect 3770 4248 3870 4251
rect 3874 4248 3878 4251
rect 3898 4248 3926 4251
rect 3930 4248 3950 4251
rect 330 4238 350 4241
rect 370 4238 590 4241
rect 778 4238 934 4241
rect 938 4238 990 4241
rect 1014 4241 1017 4248
rect 2302 4242 2305 4248
rect 2726 4242 2729 4248
rect 2918 4242 2921 4248
rect 1014 4238 1150 4241
rect 1154 4238 1206 4241
rect 1386 4238 1614 4241
rect 1618 4238 1638 4241
rect 1642 4238 1678 4241
rect 1682 4238 1918 4241
rect 2090 4238 2182 4241
rect 2462 4238 2494 4241
rect 2522 4238 2542 4241
rect 2930 4238 3366 4241
rect 3370 4238 3718 4241
rect 3794 4238 3798 4241
rect 3890 4238 3982 4241
rect 4206 4241 4209 4258
rect 4234 4248 4238 4251
rect 4322 4248 4366 4251
rect 4466 4248 4486 4251
rect 4490 4248 4558 4251
rect 4626 4248 4670 4251
rect 4698 4248 4974 4251
rect 4978 4248 5022 4251
rect 3986 4238 4209 4241
rect 4226 4238 4441 4241
rect 4482 4238 4718 4241
rect 4722 4238 4814 4241
rect 5006 4238 5070 4241
rect 130 4228 446 4231
rect 450 4228 454 4231
rect 706 4228 822 4231
rect 826 4228 1078 4231
rect 1666 4228 1686 4231
rect 1690 4228 1694 4231
rect 1930 4228 1990 4231
rect 2462 4231 2465 4238
rect 1994 4228 2465 4231
rect 2602 4228 2726 4231
rect 2754 4228 2806 4231
rect 2810 4228 2849 4231
rect 3082 4228 3526 4231
rect 3530 4228 3822 4231
rect 3834 4228 3910 4231
rect 4010 4228 4014 4231
rect 4222 4231 4225 4238
rect 4438 4232 4441 4238
rect 5006 4232 5009 4238
rect 4202 4228 4225 4231
rect 4434 4228 4438 4231
rect 4498 4228 4510 4231
rect 4786 4228 4878 4231
rect 138 4218 326 4221
rect 550 4221 553 4228
rect 2846 4222 2849 4228
rect 550 4218 670 4221
rect 1434 4218 1574 4221
rect 1586 4218 1958 4221
rect 1966 4218 2046 4221
rect 2050 4218 2454 4221
rect 3034 4218 3070 4221
rect 3074 4218 3422 4221
rect 3450 4218 3462 4221
rect 3562 4218 3646 4221
rect 3650 4218 3814 4221
rect 3874 4218 4158 4221
rect 4306 4218 4438 4221
rect 4442 4218 4462 4221
rect 4630 4221 4633 4228
rect 4626 4218 4633 4221
rect 4674 4218 4822 4221
rect 4826 4218 4854 4221
rect 98 4208 270 4211
rect 738 4208 942 4211
rect 946 4208 1230 4211
rect 1330 4208 1406 4211
rect 1618 4208 1734 4211
rect 1966 4211 1969 4218
rect 1754 4208 1969 4211
rect 2106 4208 2358 4211
rect 2418 4208 2510 4211
rect 2706 4208 2782 4211
rect 2826 4208 2966 4211
rect 3258 4208 3582 4211
rect 3634 4208 3846 4211
rect 3858 4208 3894 4211
rect 3898 4208 4126 4211
rect 4218 4208 4518 4211
rect 536 4203 538 4207
rect 542 4203 545 4207
rect 550 4203 552 4207
rect 1560 4203 1562 4207
rect 1566 4203 1569 4207
rect 1574 4203 1576 4207
rect 2584 4203 2586 4207
rect 2590 4203 2593 4207
rect 2598 4203 2600 4207
rect 3608 4203 3610 4207
rect 3614 4203 3617 4207
rect 3622 4203 3624 4207
rect 4632 4203 4634 4207
rect 4638 4203 4641 4207
rect 4646 4203 4648 4207
rect 98 4198 382 4201
rect 762 4198 886 4201
rect 914 4198 974 4201
rect 978 4198 1233 4201
rect 1634 4198 1638 4201
rect 1730 4198 1822 4201
rect 1874 4198 2206 4201
rect 2362 4198 2366 4201
rect 2370 4198 2526 4201
rect 2610 4198 2694 4201
rect 2698 4198 2854 4201
rect 2882 4198 3598 4201
rect 3778 4198 3782 4201
rect 3818 4198 4358 4201
rect 4362 4198 4382 4201
rect 4450 4198 4478 4201
rect 4482 4198 4598 4201
rect 26 4188 86 4191
rect 210 4188 262 4191
rect 418 4188 806 4191
rect 930 4188 1126 4191
rect 1178 4188 1222 4191
rect 1230 4191 1233 4198
rect 1230 4188 1974 4191
rect 2274 4188 2374 4191
rect 2394 4188 2846 4191
rect 2874 4188 2998 4191
rect 3090 4188 3134 4191
rect 3290 4188 3846 4191
rect 4458 4188 4486 4191
rect 4490 4188 4870 4191
rect 4874 4188 4886 4191
rect 4214 4182 4217 4188
rect 226 4178 358 4181
rect 434 4178 494 4181
rect 498 4178 518 4181
rect 522 4178 718 4181
rect 722 4178 1334 4181
rect 1338 4178 1910 4181
rect 2310 4178 2398 4181
rect 2490 4178 3398 4181
rect 3410 4178 3422 4181
rect 3426 4178 3526 4181
rect 3546 4178 3638 4181
rect 3794 4178 3822 4181
rect 3954 4178 3974 4181
rect 3994 4178 3998 4181
rect 4458 4178 4526 4181
rect 4570 4178 4710 4181
rect 218 4168 382 4171
rect 746 4168 766 4171
rect 954 4168 1046 4171
rect 1826 4168 1886 4171
rect 1918 4171 1921 4178
rect 2310 4172 2313 4178
rect 1918 4168 1942 4171
rect 1966 4168 1998 4171
rect 2202 4168 2262 4171
rect 2330 4168 2454 4171
rect 2458 4168 2478 4171
rect 2754 4168 2910 4171
rect 2914 4168 2918 4171
rect 2930 4168 3174 4171
rect 3226 4168 3246 4171
rect 3250 4168 3302 4171
rect 3418 4168 3438 4171
rect 3650 4168 3790 4171
rect 3922 4168 3969 4171
rect 3998 4168 4006 4171
rect 4010 4168 4078 4171
rect 4082 4168 4190 4171
rect 4202 4168 4222 4171
rect 4238 4168 4374 4171
rect 5054 4171 5057 4178
rect 4458 4168 5049 4171
rect 5054 4168 5118 4171
rect 226 4158 246 4161
rect 250 4158 254 4161
rect 322 4158 470 4161
rect 514 4158 566 4161
rect 722 4158 838 4161
rect 930 4158 950 4161
rect 986 4158 998 4161
rect 1182 4161 1185 4168
rect 1114 4158 1185 4161
rect 1198 4161 1201 4168
rect 1526 4162 1529 4168
rect 1198 4158 1222 4161
rect 1458 4158 1494 4161
rect 1710 4161 1713 4168
rect 1966 4162 1969 4168
rect 2318 4162 2321 4168
rect 3966 4162 3969 4168
rect 4238 4162 4241 4168
rect 5046 4162 5049 4168
rect 1690 4158 1713 4161
rect 1866 4158 1966 4161
rect 1990 4158 1998 4161
rect 2002 4158 2062 4161
rect 2234 4158 2286 4161
rect 2434 4158 2438 4161
rect 2474 4158 2534 4161
rect 2578 4158 2622 4161
rect 2674 4158 2678 4161
rect 2798 4158 3038 4161
rect 3042 4158 3254 4161
rect 3402 4158 3478 4161
rect 3482 4158 3638 4161
rect 3698 4158 3750 4161
rect 3850 4158 3953 4161
rect 3978 4158 4174 4161
rect 4178 4158 4238 4161
rect 4426 4158 4574 4161
rect 4658 4158 4678 4161
rect 4698 4158 4894 4161
rect 4934 4158 4942 4161
rect 4946 4158 5006 4161
rect 5050 4158 5086 4161
rect 62 4151 65 4158
rect 302 4152 305 4158
rect 2366 4152 2369 4158
rect 2798 4152 2801 4158
rect 3950 4152 3953 4158
rect 62 4148 142 4151
rect 210 4148 294 4151
rect 370 4148 374 4151
rect 426 4148 430 4151
rect 530 4148 582 4151
rect 682 4148 753 4151
rect 794 4148 798 4151
rect 850 4148 926 4151
rect 986 4148 1006 4151
rect 1014 4148 1022 4151
rect 1178 4148 1214 4151
rect 1458 4148 1526 4151
rect 1634 4148 1654 4151
rect 1714 4148 1718 4151
rect 1738 4148 1998 4151
rect 2002 4148 2158 4151
rect 2170 4148 2174 4151
rect 2178 4148 2270 4151
rect 2282 4148 2286 4151
rect 2306 4148 2318 4151
rect 2418 4148 2422 4151
rect 2442 4148 2470 4151
rect 2482 4148 2710 4151
rect 2722 4148 2726 4151
rect 2730 4148 2750 4151
rect 2794 4148 2798 4151
rect 2850 4148 2950 4151
rect 2970 4148 3078 4151
rect 3082 4148 3214 4151
rect 3250 4148 3254 4151
rect 3434 4148 3438 4151
rect 3474 4148 3558 4151
rect 3562 4148 3566 4151
rect 3602 4148 3766 4151
rect 4066 4148 4078 4151
rect 750 4142 753 4148
rect 138 4138 238 4141
rect 274 4138 278 4141
rect 286 4138 318 4141
rect 426 4138 430 4141
rect 482 4138 638 4141
rect 822 4141 825 4148
rect 1014 4142 1017 4148
rect 1310 4142 1313 4148
rect 1358 4142 1361 4148
rect 822 4138 894 4141
rect 994 4138 998 4141
rect 1042 4138 1166 4141
rect 1170 4138 1182 4141
rect 1222 4138 1230 4141
rect 1402 4138 1494 4141
rect 1610 4138 1638 4141
rect 1702 4141 1705 4148
rect 2334 4142 2337 4148
rect 4154 4148 4230 4151
rect 4350 4151 4353 4158
rect 4250 4148 4353 4151
rect 4378 4148 4526 4151
rect 4546 4148 4566 4151
rect 4626 4148 4630 4151
rect 4698 4148 4766 4151
rect 4802 4148 4822 4151
rect 4946 4148 4950 4151
rect 5058 4148 5062 4151
rect 5090 4148 5182 4151
rect 4246 4142 4249 4148
rect 1674 4138 1705 4141
rect 1722 4138 1870 4141
rect 1874 4138 1886 4141
rect 1938 4138 1966 4141
rect 2130 4138 2326 4141
rect 2394 4138 2446 4141
rect 2618 4138 2814 4141
rect 2826 4138 2862 4141
rect 2926 4138 2998 4141
rect 3090 4138 3134 4141
rect 3242 4138 3246 4141
rect 3330 4138 3454 4141
rect 3466 4138 3486 4141
rect 3586 4138 3598 4141
rect 3746 4138 3750 4141
rect 3762 4138 3782 4141
rect 3970 4138 3974 4141
rect 3978 4138 3998 4141
rect 4090 4138 4094 4141
rect 4290 4138 4398 4141
rect 4538 4138 4542 4141
rect 4554 4138 4558 4141
rect 4714 4138 4718 4141
rect 4738 4138 4870 4141
rect 5030 4138 5174 4141
rect 286 4132 289 4138
rect 342 4132 345 4138
rect 390 4132 393 4138
rect 1222 4132 1225 4138
rect 2926 4132 2929 4138
rect 3270 4132 3273 4138
rect 602 4128 830 4131
rect 890 4128 918 4131
rect 954 4128 1006 4131
rect 1250 4128 1310 4131
rect 1330 4128 1342 4131
rect 1346 4128 1358 4131
rect 1514 4128 1518 4131
rect 1698 4128 1718 4131
rect 1842 4128 2022 4131
rect 2138 4128 2142 4131
rect 2298 4128 2366 4131
rect 2450 4128 2606 4131
rect 2674 4128 2689 4131
rect 2698 4128 2710 4131
rect 2754 4128 2766 4131
rect 2778 4128 2846 4131
rect 3074 4128 3102 4131
rect 3394 4128 3478 4131
rect 3606 4131 3609 4138
rect 4478 4132 4481 4138
rect 5030 4132 5033 4138
rect 3606 4128 3766 4131
rect 3770 4128 3814 4131
rect 4210 4128 4262 4131
rect 4398 4128 4406 4131
rect 4410 4128 4422 4131
rect 4490 4128 4510 4131
rect 4754 4128 4910 4131
rect 4914 4128 4950 4131
rect 1750 4122 1753 4128
rect 346 4118 374 4121
rect 514 4118 526 4121
rect 970 4118 1262 4121
rect 1266 4118 1286 4121
rect 1298 4118 1366 4121
rect 1386 4118 1398 4121
rect 1514 4118 1566 4121
rect 1758 4121 1761 4128
rect 2686 4122 2689 4128
rect 1758 4118 1798 4121
rect 1802 4118 1854 4121
rect 1882 4118 1934 4121
rect 2042 4118 2142 4121
rect 2266 4118 2438 4121
rect 2442 4118 2502 4121
rect 2706 4118 2894 4121
rect 2906 4118 2950 4121
rect 3026 4118 3182 4121
rect 3450 4118 3478 4121
rect 3506 4118 3590 4121
rect 3594 4118 3630 4121
rect 3906 4118 3958 4121
rect 3962 4118 3982 4121
rect 3990 4121 3993 4128
rect 4430 4121 4433 4128
rect 3990 4118 4433 4121
rect 4450 4118 4566 4121
rect 466 4108 950 4111
rect 1218 4108 1294 4111
rect 1298 4108 1302 4111
rect 1314 4108 1422 4111
rect 1610 4108 1670 4111
rect 1706 4108 1982 4111
rect 1986 4108 1990 4111
rect 2274 4108 2342 4111
rect 2474 4108 2654 4111
rect 2810 4108 3030 4111
rect 3034 4108 3070 4111
rect 3146 4108 3198 4111
rect 3218 4108 3390 4111
rect 3402 4108 3470 4111
rect 3474 4108 3582 4111
rect 3666 4108 3734 4111
rect 3938 4108 4006 4111
rect 4058 4108 4086 4111
rect 4210 4108 4302 4111
rect 4338 4108 4414 4111
rect 4418 4108 4654 4111
rect 4658 4108 4814 4111
rect 1048 4103 1050 4107
rect 1054 4103 1057 4107
rect 1062 4103 1064 4107
rect 2072 4103 2074 4107
rect 2078 4103 2081 4107
rect 2086 4103 2088 4107
rect 3096 4103 3098 4107
rect 3102 4103 3105 4107
rect 3110 4103 3112 4107
rect 4112 4103 4114 4107
rect 4118 4103 4121 4107
rect 4126 4103 4128 4107
rect 490 4098 694 4101
rect 698 4098 1038 4101
rect 1290 4098 1462 4101
rect 1642 4098 1678 4101
rect 1746 4098 1846 4101
rect 2162 4098 2214 4101
rect 2266 4098 2294 4101
rect 2510 4098 2566 4101
rect 2618 4098 2702 4101
rect 2706 4098 2774 4101
rect 2794 4098 2822 4101
rect 2834 4098 2870 4101
rect 2994 4098 3006 4101
rect 3210 4098 3358 4101
rect 3538 4098 3550 4101
rect 3578 4098 3638 4101
rect 4562 4098 4646 4101
rect 4658 4098 4742 4101
rect 4882 4098 5062 4101
rect 1998 4092 2001 4098
rect 2222 4092 2225 4098
rect 106 4088 150 4091
rect 154 4088 478 4091
rect 490 4088 494 4091
rect 594 4088 630 4091
rect 666 4088 774 4091
rect 866 4088 878 4091
rect 1146 4088 1182 4091
rect 1210 4088 1222 4091
rect 1234 4088 1374 4091
rect 1378 4088 1382 4091
rect 1386 4088 1393 4091
rect 1402 4088 1646 4091
rect 1810 4088 1822 4091
rect 1918 4088 1990 4091
rect 2178 4088 2190 4091
rect 2302 4088 2305 4098
rect 2310 4092 2313 4098
rect 2510 4091 2513 4098
rect 2314 4088 2513 4091
rect 2522 4088 2526 4091
rect 2530 4088 2638 4091
rect 2762 4088 2814 4091
rect 2818 4088 2902 4091
rect 2906 4088 2982 4091
rect 3034 4088 3054 4091
rect 3058 4088 3078 4091
rect 3090 4088 3198 4091
rect 3206 4088 3214 4091
rect 3218 4088 3222 4091
rect 3226 4088 3334 4091
rect 3398 4088 3406 4091
rect 3410 4088 3446 4091
rect 3530 4088 3566 4091
rect 3578 4088 3742 4091
rect 3938 4088 3950 4091
rect 4034 4088 4062 4091
rect 4066 4088 4073 4091
rect 4082 4088 4262 4091
rect 4274 4088 4318 4091
rect 4442 4088 4702 4091
rect 4706 4088 4870 4091
rect 4890 4088 5102 4091
rect 1918 4082 1921 4088
rect 282 4078 422 4081
rect 506 4078 710 4081
rect 714 4078 1342 4081
rect 1490 4078 1518 4081
rect 1522 4078 1630 4081
rect 1730 4078 1918 4081
rect 1986 4078 2046 4081
rect 2050 4078 2246 4081
rect 2250 4078 2350 4081
rect 2426 4078 3022 4081
rect 3026 4078 3222 4081
rect 3234 4078 3742 4081
rect 3946 4078 4430 4081
rect 4586 4078 4590 4081
rect 4738 4078 4742 4081
rect 4890 4078 5030 4081
rect 42 4068 118 4071
rect 166 4071 169 4078
rect 494 4072 497 4078
rect 146 4068 169 4071
rect 458 4068 486 4071
rect 546 4068 574 4071
rect 610 4068 614 4071
rect 666 4068 670 4071
rect 690 4068 790 4071
rect 802 4068 854 4071
rect 866 4068 902 4071
rect 922 4068 926 4071
rect 962 4068 966 4071
rect 1010 4068 1046 4071
rect 1066 4068 1126 4071
rect 1154 4068 1158 4071
rect 1266 4068 1366 4071
rect 1406 4071 1409 4078
rect 1370 4068 1409 4071
rect 1418 4068 1430 4071
rect 1538 4068 1758 4071
rect 1786 4068 1886 4071
rect 1898 4068 1902 4071
rect 1938 4068 2446 4071
rect 2450 4068 2518 4071
rect 2546 4068 2582 4071
rect 2610 4068 2654 4071
rect 2762 4068 2838 4071
rect 2842 4068 2854 4071
rect 2938 4068 2961 4071
rect 310 4062 313 4068
rect 334 4062 337 4068
rect 382 4062 385 4068
rect 518 4062 521 4068
rect 582 4062 585 4068
rect 250 4058 270 4061
rect 274 4058 302 4061
rect 458 4058 462 4061
rect 466 4058 518 4061
rect 586 4058 870 4061
rect 946 4058 1014 4061
rect 1018 4058 1158 4061
rect 1194 4058 1222 4061
rect 1242 4058 1246 4061
rect 1410 4058 1414 4061
rect 1518 4061 1521 4068
rect 2958 4062 2961 4068
rect 3058 4068 3158 4071
rect 3182 4068 3246 4071
rect 3378 4068 3390 4071
rect 3410 4068 3446 4071
rect 3450 4068 3454 4071
rect 3506 4068 3510 4071
rect 3562 4068 3574 4071
rect 3578 4068 3686 4071
rect 3690 4068 3726 4071
rect 3730 4068 3758 4071
rect 3766 4068 3782 4071
rect 3994 4068 3998 4071
rect 4010 4068 4014 4071
rect 4042 4068 4070 4071
rect 4194 4068 4222 4071
rect 4234 4068 4238 4071
rect 4274 4068 4302 4071
rect 4314 4068 4318 4071
rect 4346 4068 4446 4071
rect 4490 4068 4766 4071
rect 4770 4068 4790 4071
rect 4982 4068 5001 4071
rect 1498 4058 1521 4061
rect 1530 4058 1550 4061
rect 1698 4058 1718 4061
rect 1746 4058 1766 4061
rect 1834 4058 1838 4061
rect 1898 4058 2158 4061
rect 2162 4058 2190 4061
rect 2282 4058 2302 4061
rect 2322 4058 2350 4061
rect 2394 4058 2398 4061
rect 2434 4058 2438 4061
rect 2474 4058 2678 4061
rect 2742 4058 2758 4061
rect 2818 4058 2822 4061
rect 3014 4061 3017 4068
rect 3182 4062 3185 4068
rect 3486 4062 3489 4068
rect 3550 4062 3553 4068
rect 3766 4062 3769 4068
rect 3950 4062 3953 4068
rect 4982 4062 4985 4068
rect 4998 4062 5001 4068
rect 3014 4058 3046 4061
rect 3050 4058 3094 4061
rect 3202 4058 3278 4061
rect 3386 4058 3414 4061
rect 3490 4058 3542 4061
rect 3634 4058 3654 4061
rect 3682 4058 3702 4061
rect 3730 4058 3758 4061
rect 3794 4058 3798 4061
rect 3858 4058 3902 4061
rect 3978 4058 4054 4061
rect 4058 4058 4246 4061
rect 4266 4058 4278 4061
rect 4282 4058 4334 4061
rect 4362 4058 4422 4061
rect 4426 4058 4478 4061
rect 4586 4058 4606 4061
rect 4778 4058 4854 4061
rect 102 4052 105 4058
rect 918 4052 921 4058
rect 1614 4052 1617 4058
rect 2358 4052 2361 4058
rect 2742 4052 2745 4058
rect 194 4048 281 4051
rect 330 4048 334 4051
rect 498 4048 526 4051
rect 574 4048 646 4051
rect 738 4048 902 4051
rect 1010 4048 1070 4051
rect 1074 4048 1534 4051
rect 1546 4048 1558 4051
rect 1618 4048 1934 4051
rect 1962 4048 2006 4051
rect 2026 4048 2078 4051
rect 2210 4048 2353 4051
rect 2458 4048 2574 4051
rect 2578 4048 2638 4051
rect 2642 4048 2654 4051
rect 2682 4048 2710 4051
rect 2822 4048 2830 4051
rect 2834 4048 2894 4051
rect 2934 4051 2937 4058
rect 3758 4052 3761 4058
rect 3806 4052 3809 4058
rect 2922 4048 2937 4051
rect 2954 4048 3014 4051
rect 3074 4048 3310 4051
rect 3330 4048 3334 4051
rect 3338 4048 3390 4051
rect 3474 4048 3550 4051
rect 4090 4048 4097 4051
rect 4170 4048 4174 4051
rect 4178 4048 4286 4051
rect 4302 4048 4310 4051
rect 4314 4048 4390 4051
rect 4402 4048 4614 4051
rect 4618 4048 4654 4051
rect 4682 4048 5086 4051
rect 278 4042 281 4048
rect 574 4042 577 4048
rect 2350 4042 2353 4048
rect 386 4038 438 4041
rect 474 4038 510 4041
rect 722 4038 734 4041
rect 746 4038 750 4041
rect 754 4038 878 4041
rect 882 4038 886 4041
rect 946 4038 966 4041
rect 978 4038 1230 4041
rect 1254 4038 1294 4041
rect 1314 4038 1382 4041
rect 1546 4038 1774 4041
rect 2138 4038 2142 4041
rect 2466 4038 2590 4041
rect 2594 4038 2622 4041
rect 2798 4041 2801 4048
rect 2798 4038 2830 4041
rect 3474 4038 3518 4041
rect 3634 4038 3638 4041
rect 3790 4041 3793 4048
rect 4046 4042 4049 4048
rect 4094 4042 4097 4048
rect 3790 4038 3838 4041
rect 4154 4038 4182 4041
rect 4434 4038 4446 4041
rect 4722 4038 4870 4041
rect 1254 4032 1257 4038
rect 322 4028 630 4031
rect 762 4028 814 4031
rect 818 4028 1222 4031
rect 1474 4028 1566 4031
rect 1658 4028 1814 4031
rect 1866 4028 1886 4031
rect 1914 4028 1918 4031
rect 1946 4028 1950 4031
rect 1954 4028 2150 4031
rect 2154 4028 2270 4031
rect 2338 4028 2662 4031
rect 2670 4028 3521 4031
rect 642 4018 910 4021
rect 914 4018 1022 4021
rect 1170 4018 1294 4021
rect 1626 4018 1982 4021
rect 1986 4018 2054 4021
rect 2146 4018 2230 4021
rect 2346 4018 2526 4021
rect 2534 4018 2542 4021
rect 2546 4018 2606 4021
rect 2670 4021 2673 4028
rect 3518 4022 3521 4028
rect 3758 4031 3761 4038
rect 4022 4032 4025 4038
rect 3758 4028 3814 4031
rect 3946 4028 3950 4031
rect 4154 4028 4446 4031
rect 4514 4028 4598 4031
rect 3670 4022 3673 4028
rect 2618 4018 2673 4021
rect 2690 4018 2702 4021
rect 2722 4018 2838 4021
rect 2850 4018 2990 4021
rect 2994 4018 3001 4021
rect 3010 4018 3414 4021
rect 3418 4018 3502 4021
rect 3754 4018 4134 4021
rect 4194 4018 4214 4021
rect 4218 4018 4270 4021
rect 4274 4018 4526 4021
rect 4930 4018 4958 4021
rect 146 4008 310 4011
rect 378 4008 486 4011
rect 1002 4008 1022 4011
rect 1234 4008 1270 4011
rect 1866 4008 1958 4011
rect 1962 4008 2022 4011
rect 2202 4008 2206 4011
rect 2554 4008 2558 4011
rect 2642 4008 2958 4011
rect 2962 4008 2974 4011
rect 3066 4008 3118 4011
rect 3122 4008 3214 4011
rect 3346 4008 3366 4011
rect 3370 4008 3398 4011
rect 3490 4008 3590 4011
rect 3690 4008 4286 4011
rect 4290 4008 4518 4011
rect 536 4003 538 4007
rect 542 4003 545 4007
rect 550 4003 552 4007
rect 1560 4003 1562 4007
rect 1566 4003 1569 4007
rect 1574 4003 1576 4007
rect 2584 4003 2586 4007
rect 2590 4003 2593 4007
rect 2598 4003 2600 4007
rect 3608 4003 3610 4007
rect 3614 4003 3617 4007
rect 3622 4003 3624 4007
rect 4632 4003 4634 4007
rect 4638 4003 4641 4007
rect 4646 4003 4648 4007
rect 1146 3998 1278 4001
rect 1914 3998 2374 4001
rect 2658 3998 2878 4001
rect 3290 3998 3542 4001
rect 3978 3998 3998 4001
rect 4050 3998 4126 4001
rect 4146 3998 4254 4001
rect 4266 3998 4286 4001
rect 4290 3998 4406 4001
rect 4570 3998 4590 4001
rect 4658 3998 5110 4001
rect 410 3988 742 3991
rect 826 3988 846 3991
rect 986 3988 1054 3991
rect 1242 3988 1257 3991
rect 1426 3988 1534 3991
rect 1602 3988 1726 3991
rect 1930 3988 1934 3991
rect 1970 3988 2302 3991
rect 2306 3988 2366 3991
rect 2370 3988 2542 3991
rect 2546 3988 2638 3991
rect 2658 3988 2694 3991
rect 2810 3988 2830 3991
rect 2834 3988 2974 3991
rect 3394 3988 3430 3991
rect 3594 3988 3718 3991
rect 3930 3988 4006 3991
rect 4122 3988 4278 3991
rect 4298 3988 4486 3991
rect 4538 3988 4753 3991
rect 1198 3982 1201 3988
rect 1254 3982 1257 3988
rect 362 3978 382 3981
rect 594 3978 846 3981
rect 898 3978 1014 3981
rect 1018 3978 1142 3981
rect 1154 3978 1174 3981
rect 1234 3978 1246 3981
rect 1458 3978 1502 3981
rect 1546 3978 1606 3981
rect 1610 3978 1662 3981
rect 1778 3978 1854 3981
rect 1906 3978 1926 3981
rect 1978 3978 2086 3981
rect 2226 3978 2254 3981
rect 2258 3978 2462 3981
rect 2602 3978 2902 3981
rect 3218 3978 3846 3981
rect 3850 3978 3950 3981
rect 3994 3978 3998 3981
rect 4294 3981 4297 3988
rect 4750 3982 4753 3988
rect 4218 3978 4297 3981
rect 4506 3978 4678 3981
rect 4874 3978 4926 3981
rect 5018 3978 5086 3981
rect 1142 3972 1145 3978
rect 106 3968 150 3971
rect 154 3968 593 3971
rect 590 3962 593 3968
rect 838 3968 870 3971
rect 874 3968 881 3971
rect 946 3968 950 3971
rect 1018 3968 1022 3971
rect 1042 3968 1102 3971
rect 1154 3968 1158 3971
rect 1170 3968 1174 3971
rect 1186 3968 1198 3971
rect 1210 3968 1214 3971
rect 1450 3968 1518 3971
rect 1546 3968 1550 3971
rect 1686 3971 1689 3978
rect 4102 3972 4105 3978
rect 1674 3968 1689 3971
rect 1738 3968 1902 3971
rect 1906 3968 2025 3971
rect 2162 3968 2342 3971
rect 2354 3968 2390 3971
rect 2418 3968 2606 3971
rect 2726 3968 2742 3971
rect 2762 3968 2790 3971
rect 2870 3968 2918 3971
rect 3514 3968 3518 3971
rect 4186 3968 4297 3971
rect 4306 3968 4414 3971
rect 4574 3968 4582 3971
rect 4586 3968 4598 3971
rect 4734 3971 4737 3978
rect 4734 3968 4753 3971
rect 4762 3968 4881 3971
rect 4922 3968 5046 3971
rect 838 3962 841 3968
rect 2022 3962 2025 3968
rect 250 3958 366 3961
rect 402 3958 406 3961
rect 458 3958 542 3961
rect 602 3958 678 3961
rect 858 3958 1198 3961
rect 1210 3958 1278 3961
rect 1346 3958 1726 3961
rect 1730 3958 1742 3961
rect 1778 3958 1785 3961
rect 1810 3958 1822 3961
rect 1850 3958 1862 3961
rect 1962 3958 1998 3961
rect 2170 3958 2270 3961
rect 2274 3958 2302 3961
rect 2306 3958 2398 3961
rect 2402 3958 2486 3961
rect 2662 3961 2665 3968
rect 2634 3958 2665 3961
rect 2726 3962 2729 3968
rect 2870 3962 2873 3968
rect 2738 3958 2774 3961
rect 2778 3958 2814 3961
rect 2834 3958 2838 3961
rect 2882 3958 2886 3961
rect 3406 3961 3409 3968
rect 3346 3958 3409 3961
rect 3574 3961 3577 3968
rect 3490 3958 3577 3961
rect 3850 3958 3854 3961
rect 4114 3958 4142 3961
rect 4166 3961 4169 3968
rect 4166 3958 4190 3961
rect 4234 3958 4238 3961
rect 4294 3961 4297 3968
rect 4294 3958 4305 3961
rect 4354 3958 4382 3961
rect 4386 3958 4390 3961
rect 4402 3958 4478 3961
rect 4526 3961 4529 3968
rect 4526 3958 4702 3961
rect 4706 3958 4734 3961
rect 4750 3961 4753 3968
rect 4878 3962 4881 3968
rect 4750 3958 4822 3961
rect 5098 3958 5118 3961
rect 5122 3958 5142 3961
rect 94 3952 97 3958
rect 1782 3952 1785 3958
rect 3038 3952 3041 3958
rect 114 3948 134 3951
rect 138 3948 142 3951
rect 170 3948 174 3951
rect 370 3948 406 3951
rect 450 3948 462 3951
rect 594 3948 614 3951
rect 618 3948 734 3951
rect 794 3948 870 3951
rect 950 3948 1038 3951
rect 1050 3948 1054 3951
rect 1062 3948 1078 3951
rect 1182 3948 1190 3951
rect 1306 3948 1318 3951
rect 1498 3948 1577 3951
rect 1586 3948 1678 3951
rect 1818 3948 1838 3951
rect 1890 3948 1942 3951
rect 1994 3948 2014 3951
rect 2042 3948 2046 3951
rect 2186 3948 2670 3951
rect 2674 3948 2766 3951
rect 2786 3948 2982 3951
rect 3074 3948 3182 3951
rect 3250 3948 3254 3951
rect 3274 3948 3398 3951
rect 3578 3948 3598 3951
rect 3662 3951 3665 3958
rect 3634 3948 3665 3951
rect 3766 3952 3769 3958
rect 4302 3952 4305 3958
rect 3978 3948 3990 3951
rect 4026 3948 4134 3951
rect 4178 3948 4198 3951
rect 4226 3948 4246 3951
rect 4318 3948 4326 3951
rect 4362 3948 4374 3951
rect 4442 3948 4446 3951
rect 4458 3948 4462 3951
rect 4546 3948 4550 3951
rect 4626 3948 4654 3951
rect 4690 3948 4766 3951
rect 4770 3948 4782 3951
rect 4834 3948 4886 3951
rect 4918 3951 4921 3958
rect 4918 3948 4942 3951
rect 5014 3951 5017 3958
rect 5014 3948 5070 3951
rect 734 3942 737 3948
rect 942 3942 945 3948
rect 950 3942 953 3948
rect 1062 3942 1065 3948
rect 42 3938 118 3941
rect 170 3938 190 3941
rect 330 3938 334 3941
rect 378 3938 414 3941
rect 426 3938 590 3941
rect 594 3938 710 3941
rect 858 3938 862 3941
rect 1110 3941 1113 3948
rect 1182 3942 1185 3948
rect 1098 3938 1113 3941
rect 1174 3938 1182 3941
rect 1282 3938 1390 3941
rect 1394 3938 1486 3941
rect 1490 3938 1494 3941
rect 1562 3938 1566 3941
rect 1574 3941 1577 3948
rect 1574 3938 1622 3941
rect 1646 3938 1750 3941
rect 1754 3938 1814 3941
rect 1818 3938 2006 3941
rect 2018 3938 2022 3941
rect 2058 3938 2118 3941
rect 2202 3938 2286 3941
rect 2370 3938 2374 3941
rect 2510 3938 2574 3941
rect 2578 3938 2598 3941
rect 2634 3938 2646 3941
rect 2762 3938 3014 3941
rect 3246 3941 3249 3948
rect 3018 3938 3249 3941
rect 3346 3938 3422 3941
rect 3426 3938 3462 3941
rect 3514 3938 3670 3941
rect 3814 3941 3817 3948
rect 3934 3942 3937 3948
rect 4318 3942 4321 3948
rect 4390 3942 4393 3948
rect 3814 3938 3934 3941
rect 3978 3938 4118 3941
rect 4246 3938 4254 3941
rect 4258 3938 4262 3941
rect 4558 3941 4561 3948
rect 4402 3938 4561 3941
rect 4594 3938 4638 3941
rect 4698 3938 4702 3941
rect 4906 3938 4921 3941
rect 5058 3938 5070 3941
rect 5126 3941 5129 3948
rect 5106 3938 5129 3941
rect 166 3932 169 3938
rect 1174 3932 1177 3938
rect 1646 3932 1649 3938
rect 2510 3932 2513 3938
rect 4678 3932 4681 3938
rect 4766 3932 4769 3938
rect 4918 3932 4921 3938
rect 402 3928 438 3931
rect 570 3928 670 3931
rect 1002 3928 1078 3931
rect 1082 3928 1102 3931
rect 1218 3928 1262 3931
rect 1266 3928 1374 3931
rect 1394 3928 1462 3931
rect 1466 3928 1646 3931
rect 1658 3928 1662 3931
rect 1730 3928 1766 3931
rect 1882 3928 2126 3931
rect 2130 3928 2190 3931
rect 2370 3928 2430 3931
rect 2610 3928 2726 3931
rect 2738 3928 2806 3931
rect 2858 3928 2878 3931
rect 2906 3928 3046 3931
rect 3050 3928 3390 3931
rect 3394 3928 3398 3931
rect 3418 3928 3446 3931
rect 3514 3928 3790 3931
rect 3834 3928 3838 3931
rect 3858 3928 3958 3931
rect 3994 3928 4254 3931
rect 4258 3928 4350 3931
rect 4418 3928 4502 3931
rect 4506 3928 4526 3931
rect 4586 3928 4614 3931
rect 5074 3928 5174 3931
rect 174 3921 177 3928
rect 1766 3922 1769 3928
rect 42 3918 177 3921
rect 314 3918 334 3921
rect 442 3918 478 3921
rect 746 3918 1238 3921
rect 1498 3918 1550 3921
rect 1594 3918 1686 3921
rect 1790 3912 1793 3928
rect 1810 3918 2022 3921
rect 2082 3918 2110 3921
rect 2254 3921 2257 3928
rect 2254 3918 2318 3921
rect 2338 3918 2406 3921
rect 2442 3918 2470 3921
rect 2634 3918 2654 3921
rect 2682 3918 2766 3921
rect 2822 3921 2825 3928
rect 2770 3918 2825 3921
rect 2858 3918 2862 3921
rect 3010 3918 3094 3921
rect 3138 3918 3254 3921
rect 3258 3918 3486 3921
rect 3698 3918 3894 3921
rect 3982 3921 3985 3928
rect 3922 3918 3985 3921
rect 4074 3918 4102 3921
rect 4186 3918 4190 3921
rect 4202 3918 4206 3921
rect 4242 3918 4270 3921
rect 4362 3918 4590 3921
rect 4626 3918 4902 3921
rect 4906 3918 4910 3921
rect 5098 3918 5134 3921
rect 130 3908 470 3911
rect 842 3908 918 3911
rect 1082 3908 1118 3911
rect 1122 3908 1318 3911
rect 1322 3908 1334 3911
rect 1354 3908 1590 3911
rect 1602 3908 1606 3911
rect 1642 3908 1702 3911
rect 2218 3908 2422 3911
rect 2530 3908 2774 3911
rect 2794 3908 2806 3911
rect 3018 3908 3022 3911
rect 3378 3908 3382 3911
rect 3402 3908 3502 3911
rect 3506 3908 3734 3911
rect 3762 3908 4038 3911
rect 4178 3908 4334 3911
rect 4346 3908 4654 3911
rect 5026 3908 5102 3911
rect 958 3902 961 3908
rect 1048 3903 1050 3907
rect 1054 3903 1057 3907
rect 1062 3903 1064 3907
rect 2072 3903 2074 3907
rect 2078 3903 2081 3907
rect 2086 3903 2088 3907
rect 3096 3903 3098 3907
rect 3102 3903 3105 3907
rect 3110 3903 3112 3907
rect 4112 3903 4114 3907
rect 4118 3903 4121 3907
rect 4126 3903 4128 3907
rect 98 3898 206 3901
rect 210 3898 342 3901
rect 666 3898 742 3901
rect 1154 3898 1310 3901
rect 1314 3898 1342 3901
rect 1370 3898 1398 3901
rect 1434 3898 1470 3901
rect 1506 3898 1798 3901
rect 2106 3898 2262 3901
rect 2290 3898 2518 3901
rect 2562 3898 2982 3901
rect 3146 3898 3238 3901
rect 3378 3898 3558 3901
rect 3882 3898 3974 3901
rect 4138 3898 4174 3901
rect 4182 3898 4366 3901
rect 4378 3898 4534 3901
rect 4546 3898 4558 3901
rect 4562 3898 4662 3901
rect 114 3888 198 3891
rect 274 3888 1102 3891
rect 1106 3888 1113 3891
rect 1122 3888 1142 3891
rect 1194 3888 1238 3891
rect 1266 3888 1374 3891
rect 1538 3888 1825 3891
rect 1938 3888 2022 3891
rect 2066 3888 2814 3891
rect 2818 3888 3662 3891
rect 3682 3888 3702 3891
rect 3798 3888 3806 3891
rect 3810 3888 4054 3891
rect 4182 3891 4185 3898
rect 4066 3888 4185 3891
rect 4226 3888 4254 3891
rect 4458 3888 4462 3891
rect 4482 3888 4494 3891
rect 4550 3888 4702 3891
rect 4818 3888 4878 3891
rect 4882 3888 4934 3891
rect 4954 3888 4990 3891
rect 4994 3888 5078 3891
rect 266 3878 366 3881
rect 410 3878 414 3881
rect 906 3878 910 3881
rect 914 3878 1158 3881
rect 1162 3878 1166 3881
rect 1202 3878 1334 3881
rect 1338 3878 1446 3881
rect 1462 3881 1465 3888
rect 1822 3882 1825 3888
rect 4550 3882 4553 3888
rect 1462 3878 1614 3881
rect 1638 3878 1646 3881
rect 1650 3878 1654 3881
rect 1698 3878 1710 3881
rect 1746 3878 1750 3881
rect 1850 3878 1870 3881
rect 1882 3878 1886 3881
rect 2242 3878 2262 3881
rect 2330 3878 2342 3881
rect 2414 3878 2422 3881
rect 2490 3878 2510 3881
rect 2538 3878 2614 3881
rect 2626 3878 2737 3881
rect 2762 3878 2846 3881
rect 2850 3878 2950 3881
rect 3018 3878 3270 3881
rect 3434 3878 3438 3881
rect 3754 3878 3838 3881
rect 4090 3878 4134 3881
rect 4170 3878 4214 3881
rect 4266 3878 4550 3881
rect 4578 3878 4598 3881
rect 4818 3878 4918 3881
rect 182 3871 185 3878
rect 182 3868 281 3871
rect 378 3868 430 3871
rect 498 3868 566 3871
rect 730 3868 774 3871
rect 838 3871 841 3878
rect 2734 3872 2737 3878
rect 4230 3872 4233 3878
rect 4246 3872 4249 3878
rect 778 3868 841 3871
rect 882 3868 926 3871
rect 970 3868 974 3871
rect 1002 3868 1022 3871
rect 1034 3868 1062 3871
rect 1146 3868 1150 3871
rect 1162 3868 1302 3871
rect 1370 3868 1414 3871
rect 1442 3868 1446 3871
rect 1482 3868 1558 3871
rect 1578 3868 1622 3871
rect 1626 3868 1798 3871
rect 1818 3868 1854 3871
rect 1882 3868 1886 3871
rect 1994 3868 2062 3871
rect 2130 3868 2142 3871
rect 2250 3868 2334 3871
rect 2346 3868 2630 3871
rect 2778 3868 2782 3871
rect 2922 3868 2958 3871
rect 2962 3868 2969 3871
rect 2978 3868 2998 3871
rect 3042 3868 3046 3871
rect 3066 3868 3070 3871
rect 3226 3868 3254 3871
rect 3266 3868 3270 3871
rect 3474 3868 3542 3871
rect 3610 3868 3614 3871
rect 3714 3868 3750 3871
rect 3946 3868 3982 3871
rect 3986 3868 3993 3871
rect 4058 3868 4150 3871
rect 4250 3868 4270 3871
rect 4322 3868 4374 3871
rect 4378 3868 4398 3871
rect 4434 3868 4582 3871
rect 4634 3868 4662 3871
rect 4770 3868 4830 3871
rect 4858 3868 4934 3871
rect 5018 3868 5094 3871
rect 278 3862 281 3868
rect 1022 3862 1025 3868
rect 1094 3862 1097 3868
rect 2198 3862 2201 3868
rect 234 3858 246 3861
rect 266 3858 270 3861
rect 330 3858 486 3861
rect 610 3858 718 3861
rect 770 3858 782 3861
rect 874 3858 1006 3861
rect 1054 3858 1070 3861
rect 1114 3858 1358 3861
rect 1482 3858 1486 3861
rect 1502 3858 1526 3861
rect 1554 3858 1590 3861
rect 1594 3858 1638 3861
rect 1734 3858 1758 3861
rect 1786 3858 1870 3861
rect 1874 3858 2038 3861
rect 2042 3858 2086 3861
rect 2090 3858 2126 3861
rect 2306 3858 2374 3861
rect 2418 3858 2425 3861
rect 2434 3858 2438 3861
rect 2562 3858 2569 3861
rect 2594 3858 2598 3861
rect 2646 3861 2649 3868
rect 3382 3862 3385 3868
rect 2626 3858 2649 3861
rect 2778 3858 2782 3861
rect 2810 3858 2942 3861
rect 2954 3858 2958 3861
rect 2962 3858 2990 3861
rect 3002 3858 3006 3861
rect 3082 3858 3246 3861
rect 3250 3858 3294 3861
rect 3370 3858 3374 3861
rect 3414 3861 3417 3868
rect 3446 3861 3449 3868
rect 3414 3858 3449 3861
rect 3498 3858 3526 3861
rect 3774 3861 3777 3868
rect 3690 3858 3777 3861
rect 3994 3858 4014 3861
rect 4022 3858 4070 3861
rect 4074 3858 4134 3861
rect 4162 3858 4214 3861
rect 4218 3858 4286 3861
rect 4378 3858 4398 3861
rect 4434 3858 4438 3861
rect 4446 3858 4462 3861
rect 4474 3858 4478 3861
rect 4490 3858 4526 3861
rect 4530 3858 4758 3861
rect 4762 3858 4822 3861
rect 4826 3858 4886 3861
rect 5014 3861 5017 3868
rect 4898 3858 5017 3861
rect 5082 3858 5086 3861
rect 822 3852 825 3858
rect 1054 3852 1057 3858
rect 1502 3852 1505 3858
rect 170 3848 225 3851
rect 322 3848 406 3851
rect 1002 3848 1014 3851
rect 1066 3848 1078 3851
rect 1162 3848 1206 3851
rect 1330 3848 1334 3851
rect 1350 3848 1358 3851
rect 1410 3848 1438 3851
rect 1734 3851 1737 3858
rect 2158 3852 2161 3858
rect 2422 3852 2425 3858
rect 2566 3852 2569 3858
rect 2726 3852 2729 3858
rect 3334 3852 3337 3858
rect 3342 3852 3345 3858
rect 4022 3852 4025 3858
rect 1582 3848 1737 3851
rect 1746 3848 1878 3851
rect 2330 3848 2358 3851
rect 2402 3848 2406 3851
rect 2746 3848 2766 3851
rect 2994 3848 3054 3851
rect 3074 3848 3214 3851
rect 3242 3848 3254 3851
rect 3682 3848 3718 3851
rect 3778 3848 3822 3851
rect 3946 3848 3998 3851
rect 4106 3848 4166 3851
rect 4246 3848 4254 3851
rect 4258 3848 4318 3851
rect 4446 3851 4449 3858
rect 4394 3848 4449 3851
rect 4466 3848 4502 3851
rect 4810 3848 4870 3851
rect 4874 3848 4918 3851
rect 5078 3848 5150 3851
rect 222 3842 225 3848
rect 1350 3842 1353 3848
rect 1582 3842 1585 3848
rect 930 3838 974 3841
rect 1074 3838 1118 3841
rect 1154 3838 1174 3841
rect 1418 3838 1510 3841
rect 1642 3838 1702 3841
rect 1802 3838 1814 3841
rect 2042 3838 2342 3841
rect 2346 3838 2606 3841
rect 2746 3838 2870 3841
rect 3230 3841 3233 3848
rect 3654 3842 3657 3848
rect 4542 3842 4545 3848
rect 5054 3842 5057 3848
rect 5078 3842 5081 3848
rect 3210 3838 3233 3841
rect 3250 3838 3350 3841
rect 3490 3838 3494 3841
rect 3586 3838 3638 3841
rect 4002 3838 4142 3841
rect 4146 3838 4198 3841
rect 4418 3838 4422 3841
rect 4754 3838 4846 3841
rect 4850 3838 4878 3841
rect 206 3831 209 3838
rect 206 3828 390 3831
rect 706 3828 918 3831
rect 1034 3828 1334 3831
rect 1338 3828 1430 3831
rect 1510 3828 1606 3831
rect 1714 3828 1806 3831
rect 2074 3828 2110 3831
rect 2306 3828 2446 3831
rect 2546 3828 2702 3831
rect 2722 3828 2750 3831
rect 2754 3828 2918 3831
rect 2946 3828 3022 3831
rect 3090 3828 3398 3831
rect 3402 3828 3414 3831
rect 3418 3828 3494 3831
rect 3498 3828 3574 3831
rect 3602 3828 3782 3831
rect 3850 3828 3862 3831
rect 3874 3828 4254 3831
rect 4262 3831 4265 3838
rect 4262 3828 4382 3831
rect 4402 3828 4726 3831
rect 5058 3828 5086 3831
rect 306 3818 334 3821
rect 362 3818 366 3821
rect 426 3818 462 3821
rect 482 3818 686 3821
rect 1510 3821 1513 3828
rect 810 3818 1513 3821
rect 1522 3818 1830 3821
rect 1866 3818 1926 3821
rect 1930 3818 2310 3821
rect 2338 3818 2374 3821
rect 2378 3818 2398 3821
rect 2690 3818 2790 3821
rect 3362 3818 3718 3821
rect 3898 3818 3902 3821
rect 3962 3818 4014 3821
rect 4018 3818 4086 3821
rect 4090 3818 4174 3821
rect 4362 3818 4462 3821
rect 4586 3818 4966 3821
rect 4970 3818 5070 3821
rect 2542 3812 2545 3818
rect 378 3808 526 3811
rect 938 3808 1094 3811
rect 1170 3808 1206 3811
rect 1218 3808 1534 3811
rect 1586 3808 1846 3811
rect 1850 3808 2110 3811
rect 2258 3808 2310 3811
rect 2322 3808 2374 3811
rect 2386 3808 2414 3811
rect 2634 3808 2838 3811
rect 2842 3808 2950 3811
rect 3266 3808 3382 3811
rect 3666 3808 4190 3811
rect 4386 3808 4422 3811
rect 4450 3808 4486 3811
rect 536 3803 538 3807
rect 542 3803 545 3807
rect 550 3803 552 3807
rect 1560 3803 1562 3807
rect 1566 3803 1569 3807
rect 1574 3803 1576 3807
rect 2584 3803 2586 3807
rect 2590 3803 2593 3807
rect 2598 3803 2600 3807
rect 3608 3803 3610 3807
rect 3614 3803 3617 3807
rect 3622 3803 3624 3807
rect 4632 3803 4634 3807
rect 4638 3803 4641 3807
rect 4646 3803 4648 3807
rect 250 3798 430 3801
rect 890 3798 910 3801
rect 914 3798 934 3801
rect 938 3798 1142 3801
rect 1170 3798 1350 3801
rect 1858 3798 1862 3801
rect 1870 3798 2166 3801
rect 2194 3798 2534 3801
rect 2634 3798 2798 3801
rect 3714 3798 3718 3801
rect 3794 3798 3950 3801
rect 3954 3798 4006 3801
rect 4130 3798 4198 3801
rect 4202 3798 4238 3801
rect 418 3788 742 3791
rect 898 3788 1462 3791
rect 1490 3788 1753 3791
rect 1870 3791 1873 3798
rect 1858 3788 1873 3791
rect 1898 3788 2278 3791
rect 2282 3788 2382 3791
rect 2394 3788 2606 3791
rect 2666 3788 2806 3791
rect 2834 3788 2966 3791
rect 3370 3788 3446 3791
rect 3578 3788 4470 3791
rect 4474 3788 4694 3791
rect 4698 3788 4734 3791
rect 4882 3788 4982 3791
rect 406 3781 409 3788
rect 1750 3782 1753 3788
rect 138 3778 409 3781
rect 530 3778 766 3781
rect 810 3778 838 3781
rect 954 3778 1078 3781
rect 1306 3778 1350 3781
rect 1450 3778 1697 3781
rect 1770 3778 1782 3781
rect 1826 3778 2273 3781
rect 1694 3772 1697 3778
rect 2270 3772 2273 3778
rect 2554 3778 2662 3781
rect 2786 3778 2878 3781
rect 3002 3778 3390 3781
rect 3538 3778 3814 3781
rect 3898 3778 4350 3781
rect 4358 3778 4710 3781
rect 4770 3778 4990 3781
rect 362 3768 654 3771
rect 778 3768 902 3771
rect 906 3768 1022 3771
rect 1106 3768 1286 3771
rect 1330 3768 1358 3771
rect 1698 3768 1726 3771
rect 1730 3768 1737 3771
rect 1762 3768 1766 3771
rect 1894 3768 2014 3771
rect 2018 3768 2246 3771
rect 2390 3771 2393 3778
rect 2354 3768 2393 3771
rect 2762 3768 3014 3771
rect 3026 3768 3286 3771
rect 3330 3768 3366 3771
rect 3546 3768 3638 3771
rect 3642 3768 3686 3771
rect 3714 3768 3886 3771
rect 3994 3768 4238 3771
rect 4358 3771 4361 3778
rect 4330 3768 4361 3771
rect 4366 3768 5086 3771
rect 5090 3768 5134 3771
rect 106 3758 310 3761
rect 354 3758 422 3761
rect 594 3758 750 3761
rect 754 3758 814 3761
rect 954 3758 958 3761
rect 970 3758 1006 3761
rect 1034 3758 1118 3761
rect 1138 3758 1262 3761
rect 1326 3761 1329 3768
rect 1894 3762 1897 3768
rect 3374 3762 3377 3768
rect 4366 3762 4369 3768
rect 1306 3758 1329 3761
rect 1594 3758 1750 3761
rect 1754 3758 1878 3761
rect 2034 3758 2038 3761
rect 2058 3758 2174 3761
rect 2202 3758 2206 3761
rect 2234 3758 2518 3761
rect 2522 3758 2534 3761
rect 2578 3758 2598 3761
rect 2602 3758 2670 3761
rect 2706 3758 2854 3761
rect 2898 3758 2902 3761
rect 2914 3758 3030 3761
rect 3250 3758 3334 3761
rect 3594 3758 3606 3761
rect 3642 3758 3678 3761
rect 3682 3758 3814 3761
rect 3874 3758 4126 3761
rect 4226 3758 4294 3761
rect 4314 3758 4342 3761
rect 4594 3758 4609 3761
rect 4714 3758 4734 3761
rect 5002 3758 5014 3761
rect 418 3748 430 3751
rect 434 3748 686 3751
rect 690 3748 710 3751
rect 890 3748 982 3751
rect 994 3748 1134 3751
rect 1154 3748 1302 3751
rect 1342 3748 1414 3751
rect 1626 3748 1646 3751
rect 1810 3748 1814 3751
rect 1910 3751 1913 3758
rect 1958 3751 1961 3758
rect 2230 3752 2233 3758
rect 1858 3748 1865 3751
rect 1910 3748 1961 3751
rect 1986 3748 2118 3751
rect 2138 3748 2214 3751
rect 2266 3748 2270 3751
rect 2386 3748 2414 3751
rect 2466 3748 2478 3751
rect 2482 3748 2486 3751
rect 2498 3748 2638 3751
rect 2642 3748 2822 3751
rect 2842 3748 2865 3751
rect 2882 3748 2918 3751
rect 3130 3748 3206 3751
rect 3210 3748 3230 3751
rect 3402 3748 3406 3751
rect 3530 3748 3574 3751
rect 3586 3748 3617 3751
rect 382 3742 385 3748
rect 686 3742 689 3748
rect 1342 3742 1345 3748
rect 322 3738 350 3741
rect 802 3738 894 3741
rect 906 3738 942 3741
rect 978 3738 1070 3741
rect 1142 3738 1150 3741
rect 1314 3738 1318 3741
rect 1370 3738 1390 3741
rect 1494 3741 1497 3748
rect 1670 3742 1673 3748
rect 1418 3738 1497 3741
rect 1522 3738 1638 3741
rect 1686 3741 1689 3748
rect 1862 3742 1865 3748
rect 1682 3738 1689 3741
rect 1714 3738 1718 3741
rect 1722 3738 1838 3741
rect 1866 3738 2382 3741
rect 2426 3738 2430 3741
rect 2446 3741 2449 3748
rect 2862 3742 2865 3748
rect 2446 3738 2518 3741
rect 2570 3738 2574 3741
rect 2618 3738 2622 3741
rect 2666 3738 2766 3741
rect 2850 3738 2854 3741
rect 2866 3738 2894 3741
rect 2906 3738 2974 3741
rect 2998 3741 3001 3748
rect 2998 3738 3078 3741
rect 3110 3741 3113 3748
rect 3082 3738 3113 3741
rect 3262 3741 3265 3748
rect 3162 3738 3265 3741
rect 3322 3738 3358 3741
rect 3510 3741 3513 3748
rect 3614 3742 3617 3748
rect 3706 3748 3710 3751
rect 3722 3748 3726 3751
rect 3738 3748 3742 3751
rect 3754 3748 3798 3751
rect 3670 3742 3673 3748
rect 3810 3748 3830 3751
rect 3898 3748 3902 3751
rect 3970 3748 3985 3751
rect 3994 3748 4198 3751
rect 4314 3748 4318 3751
rect 4410 3748 4510 3751
rect 4606 3751 4609 3758
rect 4606 3748 4710 3751
rect 5038 3751 5041 3758
rect 4986 3748 5041 3751
rect 5126 3751 5129 3758
rect 5082 3748 5129 3751
rect 3982 3742 3985 3748
rect 4574 3742 4577 3748
rect 4598 3742 4601 3748
rect 3510 3738 3598 3741
rect 3858 3738 3862 3741
rect 4050 3738 4054 3741
rect 4082 3738 4118 3741
rect 4154 3738 4206 3741
rect 4266 3738 4558 3741
rect 4650 3738 4686 3741
rect 4726 3741 4729 3748
rect 4726 3738 4750 3741
rect 4762 3738 5102 3741
rect 206 3731 209 3738
rect 670 3732 673 3738
rect 1142 3732 1145 3738
rect 1174 3732 1177 3738
rect 2646 3732 2649 3738
rect 3662 3732 3665 3738
rect 3934 3732 3937 3738
rect 4606 3732 4609 3738
rect 4686 3732 4689 3738
rect 206 3728 398 3731
rect 450 3728 590 3731
rect 594 3728 646 3731
rect 778 3728 1094 3731
rect 1234 3728 2030 3731
rect 2058 3728 2094 3731
rect 2178 3728 2262 3731
rect 2266 3728 2342 3731
rect 2370 3728 2502 3731
rect 2698 3728 2782 3731
rect 3214 3728 3278 3731
rect 3522 3728 3526 3731
rect 3546 3728 3558 3731
rect 3562 3728 3654 3731
rect 3802 3728 3870 3731
rect 4290 3728 4390 3731
rect 4738 3728 4742 3731
rect 4906 3728 5038 3731
rect 274 3718 294 3721
rect 354 3718 358 3721
rect 398 3721 401 3728
rect 3214 3722 3217 3728
rect 3846 3722 3849 3728
rect 398 3718 718 3721
rect 866 3718 990 3721
rect 1018 3718 1110 3721
rect 1130 3718 1294 3721
rect 1450 3718 1478 3721
rect 1482 3718 1542 3721
rect 1698 3718 1718 3721
rect 1738 3718 1766 3721
rect 1770 3718 1870 3721
rect 2034 3718 2126 3721
rect 2210 3718 2230 3721
rect 2282 3718 2382 3721
rect 2402 3718 2438 3721
rect 2466 3718 2478 3721
rect 2634 3718 2870 3721
rect 2874 3718 3198 3721
rect 3234 3718 3406 3721
rect 3430 3718 3438 3721
rect 3498 3718 3526 3721
rect 4338 3718 4398 3721
rect 4426 3718 4662 3721
rect 4674 3718 4694 3721
rect 4826 3718 4974 3721
rect 2606 3712 2609 3718
rect 3430 3712 3433 3718
rect 306 3708 670 3711
rect 1074 3708 1278 3711
rect 1330 3708 1398 3711
rect 1730 3708 1934 3711
rect 2202 3708 2590 3711
rect 2642 3708 3030 3711
rect 3146 3708 3190 3711
rect 3338 3708 3414 3711
rect 3538 3708 3590 3711
rect 3698 3708 3718 3711
rect 3882 3708 4094 3711
rect 4194 3708 4438 3711
rect 4922 3708 5190 3711
rect 1048 3703 1050 3707
rect 1054 3703 1057 3707
rect 1062 3703 1064 3707
rect 2072 3703 2074 3707
rect 2078 3703 2081 3707
rect 2086 3703 2088 3707
rect 3096 3703 3098 3707
rect 3102 3703 3105 3707
rect 3110 3703 3112 3707
rect 4112 3703 4114 3707
rect 4118 3703 4121 3707
rect 4126 3703 4128 3707
rect 338 3698 358 3701
rect 370 3698 382 3701
rect 514 3698 542 3701
rect 578 3698 630 3701
rect 634 3698 726 3701
rect 730 3698 766 3701
rect 794 3698 822 3701
rect 1034 3698 1038 3701
rect 1106 3698 1118 3701
rect 1206 3698 1350 3701
rect 1354 3698 1398 3701
rect 1514 3698 1606 3701
rect 1722 3698 1742 3701
rect 1810 3698 1910 3701
rect 2138 3698 2262 3701
rect 2266 3698 2318 3701
rect 2378 3698 2566 3701
rect 2570 3698 2622 3701
rect 2626 3698 2806 3701
rect 2826 3698 2894 3701
rect 2898 3698 3014 3701
rect 3258 3698 3374 3701
rect 3394 3698 3398 3701
rect 3426 3698 3553 3701
rect 3642 3698 3766 3701
rect 3770 3698 3998 3701
rect 4266 3698 4270 3701
rect 4282 3698 4342 3701
rect 4370 3698 4382 3701
rect 4418 3698 4686 3701
rect 4706 3698 4734 3701
rect 4786 3698 4990 3701
rect 10 3688 374 3691
rect 402 3688 406 3691
rect 466 3688 782 3691
rect 786 3688 838 3691
rect 1206 3691 1209 3698
rect 3550 3692 3553 3698
rect 1026 3688 1209 3691
rect 1306 3688 1582 3691
rect 1594 3688 1726 3691
rect 1762 3688 1798 3691
rect 1850 3688 1878 3691
rect 1890 3688 2102 3691
rect 2266 3688 2550 3691
rect 2658 3688 2734 3691
rect 2818 3688 3086 3691
rect 3094 3688 3102 3691
rect 3106 3688 3134 3691
rect 3390 3688 3398 3691
rect 3402 3688 3430 3691
rect 3466 3688 3470 3691
rect 3554 3688 3566 3691
rect 3570 3688 3630 3691
rect 3650 3688 3662 3691
rect 3666 3688 3694 3691
rect 3850 3688 3854 3691
rect 3922 3688 3926 3691
rect 3978 3688 4014 3691
rect 4226 3688 4270 3691
rect 4666 3688 4710 3691
rect 4778 3688 4830 3691
rect 4962 3688 5054 3691
rect 98 3678 174 3681
rect 314 3678 478 3681
rect 818 3678 854 3681
rect 938 3678 974 3681
rect 1006 3681 1009 3688
rect 1002 3678 1009 3681
rect 1082 3678 1102 3681
rect 1170 3678 1310 3681
rect 1394 3678 1470 3681
rect 1586 3678 1590 3681
rect 1698 3678 1702 3681
rect 1722 3678 1782 3681
rect 1818 3678 1854 3681
rect 1898 3678 1902 3681
rect 2034 3678 2150 3681
rect 2402 3678 2462 3681
rect 2482 3678 2574 3681
rect 2794 3678 3102 3681
rect 3122 3678 3718 3681
rect 3858 3678 3942 3681
rect 3978 3678 4046 3681
rect 4186 3678 4358 3681
rect 4682 3678 4774 3681
rect 4802 3678 4878 3681
rect 4882 3678 4926 3681
rect 58 3668 158 3671
rect 226 3668 446 3671
rect 482 3668 486 3671
rect 578 3668 646 3671
rect 650 3668 678 3671
rect 762 3668 910 3671
rect 954 3668 1038 3671
rect 1098 3668 1158 3671
rect 1366 3671 1369 3678
rect 1598 3672 1601 3678
rect 2358 3672 2361 3678
rect 2750 3672 2753 3678
rect 1266 3668 1369 3671
rect 1466 3668 1470 3671
rect 1530 3668 1534 3671
rect 1562 3668 1593 3671
rect 1618 3668 1846 3671
rect 1930 3668 1982 3671
rect 2010 3668 2046 3671
rect 2282 3668 2286 3671
rect 2314 3668 2334 3671
rect 2394 3668 2462 3671
rect 2522 3668 2526 3671
rect 2530 3668 2542 3671
rect 2626 3668 2654 3671
rect 2786 3668 2801 3671
rect 2914 3668 2942 3671
rect 2954 3668 2966 3671
rect 3098 3668 3126 3671
rect 3250 3668 3270 3671
rect 3298 3668 3390 3671
rect 3402 3668 3422 3671
rect 3450 3668 3462 3671
rect 3514 3668 3534 3671
rect 3570 3668 3718 3671
rect 3734 3671 3737 3678
rect 3734 3668 3814 3671
rect 3818 3668 3830 3671
rect 3834 3668 3910 3671
rect 3914 3668 3990 3671
rect 4018 3668 4070 3671
rect 4242 3668 4254 3671
rect 4358 3671 4361 3678
rect 4358 3668 4502 3671
rect 4606 3671 4609 3678
rect 5086 3672 5089 3678
rect 4606 3668 4750 3671
rect 4826 3668 4846 3671
rect 4898 3668 4982 3671
rect 5026 3668 5046 3671
rect 5106 3668 5110 3671
rect 5154 3668 5166 3671
rect 1078 3662 1081 3668
rect 1222 3662 1225 3668
rect 34 3658 46 3661
rect 50 3658 166 3661
rect 170 3658 230 3661
rect 234 3658 254 3661
rect 258 3658 318 3661
rect 322 3658 358 3661
rect 362 3658 462 3661
rect 474 3658 502 3661
rect 570 3658 606 3661
rect 770 3658 886 3661
rect 962 3658 974 3661
rect 1018 3658 1038 3661
rect 1114 3658 1118 3661
rect 1130 3658 1142 3661
rect 1170 3658 1206 3661
rect 1474 3658 1574 3661
rect 1590 3661 1593 3668
rect 1902 3662 1905 3668
rect 1578 3658 1585 3661
rect 1590 3658 1614 3661
rect 1650 3658 1662 3661
rect 1738 3658 1750 3661
rect 1782 3658 1790 3661
rect 1818 3658 1822 3661
rect 1838 3658 1894 3661
rect 1938 3658 1953 3661
rect 718 3652 721 3658
rect 942 3652 945 3658
rect 1782 3652 1785 3658
rect 1838 3652 1841 3658
rect 1950 3652 1953 3658
rect 1974 3658 1982 3661
rect 2166 3661 2169 3668
rect 2114 3659 2169 3661
rect 2110 3658 2169 3659
rect 2330 3658 2422 3661
rect 2450 3658 2526 3661
rect 2714 3658 2790 3661
rect 2798 3661 2801 3668
rect 2798 3658 2902 3661
rect 2962 3659 2998 3661
rect 2962 3658 3001 3659
rect 3074 3658 3238 3661
rect 3250 3658 3254 3661
rect 3330 3658 3390 3661
rect 3410 3658 3438 3661
rect 3442 3658 3446 3661
rect 3458 3658 3470 3661
rect 3522 3658 3542 3661
rect 3570 3658 3694 3661
rect 3698 3658 3846 3661
rect 3874 3658 3878 3661
rect 3930 3658 3990 3661
rect 4002 3658 4009 3661
rect 4066 3658 4150 3661
rect 4266 3658 4270 3661
rect 4362 3658 4377 3661
rect 4450 3658 4454 3661
rect 4474 3658 4486 3661
rect 4706 3658 4710 3661
rect 4850 3658 4854 3661
rect 4882 3658 4910 3661
rect 4914 3658 5030 3661
rect 5034 3658 5062 3661
rect 5066 3658 5110 3661
rect 1974 3652 1977 3658
rect 2614 3652 2617 3658
rect 4006 3652 4009 3658
rect 4374 3652 4377 3658
rect 4622 3652 4625 3658
rect 282 3648 446 3651
rect 450 3648 454 3651
rect 650 3648 694 3651
rect 882 3648 926 3651
rect 994 3648 1014 3651
rect 1078 3648 1086 3651
rect 1090 3648 1150 3651
rect 1186 3648 1318 3651
rect 1322 3648 1406 3651
rect 1490 3648 1494 3651
rect 1530 3648 1582 3651
rect 1594 3648 1678 3651
rect 2002 3648 2038 3651
rect 2162 3648 2182 3651
rect 2186 3648 2190 3651
rect 2242 3648 2366 3651
rect 2370 3648 2406 3651
rect 2650 3648 2662 3651
rect 2682 3648 2774 3651
rect 2938 3648 3046 3651
rect 3186 3648 3422 3651
rect 3450 3648 3454 3651
rect 3578 3648 3686 3651
rect 3706 3648 3854 3651
rect 3874 3648 3942 3651
rect 4258 3648 4318 3651
rect 4458 3648 4462 3651
rect 4494 3648 4582 3651
rect 4698 3648 4798 3651
rect 4826 3648 4841 3651
rect 150 3641 153 3648
rect 190 3641 193 3648
rect 4494 3642 4497 3648
rect 4838 3642 4841 3648
rect 150 3638 193 3641
rect 306 3638 398 3641
rect 442 3638 470 3641
rect 530 3638 614 3641
rect 690 3638 766 3641
rect 882 3638 998 3641
rect 1002 3638 1278 3641
rect 1282 3638 1958 3641
rect 2338 3638 2454 3641
rect 2554 3638 2686 3641
rect 2730 3638 3062 3641
rect 3066 3638 3430 3641
rect 3594 3638 3598 3641
rect 3686 3638 3694 3641
rect 3698 3638 3758 3641
rect 3770 3638 3886 3641
rect 3946 3638 4094 3641
rect 4098 3638 4206 3641
rect 4258 3638 4406 3641
rect 4690 3638 4702 3641
rect 4714 3638 4726 3641
rect 4730 3638 4806 3641
rect 122 3628 166 3631
rect 394 3628 406 3631
rect 458 3628 654 3631
rect 658 3628 870 3631
rect 898 3628 934 3631
rect 1214 3628 1254 3631
rect 1442 3628 1526 3631
rect 1594 3628 1702 3631
rect 1978 3628 2374 3631
rect 3082 3628 3118 3631
rect 3122 3628 3310 3631
rect 3430 3631 3433 3638
rect 3430 3628 4086 3631
rect 4106 3628 4110 3631
rect 4186 3628 4190 3631
rect 4362 3628 4406 3631
rect 4630 3628 4638 3631
rect 4642 3628 4654 3631
rect 4666 3628 4726 3631
rect 1214 3622 1217 3628
rect 418 3618 729 3621
rect 738 3618 902 3621
rect 906 3618 1038 3621
rect 1234 3618 1526 3621
rect 1582 3621 1585 3628
rect 1582 3618 1590 3621
rect 1602 3618 1822 3621
rect 1826 3618 1918 3621
rect 1922 3618 2166 3621
rect 2330 3618 2494 3621
rect 2498 3618 2702 3621
rect 2706 3618 3406 3621
rect 3410 3618 3430 3621
rect 3586 3618 3745 3621
rect 3754 3618 3958 3621
rect 4322 3618 4478 3621
rect 4482 3618 4670 3621
rect 5082 3618 5134 3621
rect 194 3608 374 3611
rect 726 3611 729 3618
rect 726 3608 1030 3611
rect 1282 3608 1310 3611
rect 1658 3608 1942 3611
rect 1946 3608 1998 3611
rect 2130 3608 2398 3611
rect 2522 3608 2558 3611
rect 2618 3608 2646 3611
rect 3034 3608 3350 3611
rect 3378 3608 3390 3611
rect 3394 3608 3502 3611
rect 3650 3608 3734 3611
rect 3742 3611 3745 3618
rect 3742 3608 3934 3611
rect 3938 3608 4366 3611
rect 4658 3608 4774 3611
rect 536 3603 538 3607
rect 542 3603 545 3607
rect 550 3603 552 3607
rect 1560 3603 1562 3607
rect 1566 3603 1569 3607
rect 1574 3603 1576 3607
rect 2584 3603 2586 3607
rect 2590 3603 2593 3607
rect 2598 3603 2600 3607
rect 3608 3603 3610 3607
rect 3614 3603 3617 3607
rect 3622 3603 3624 3607
rect 4632 3603 4634 3607
rect 4638 3603 4641 3607
rect 4646 3603 4648 3607
rect 10 3598 278 3601
rect 1138 3598 1246 3601
rect 1250 3598 1286 3601
rect 1386 3598 1478 3601
rect 1482 3598 1486 3601
rect 1586 3598 1662 3601
rect 1746 3598 1750 3601
rect 1778 3598 1838 3601
rect 1898 3598 1918 3601
rect 2714 3598 2726 3601
rect 2978 3598 3582 3601
rect 3778 3598 3798 3601
rect 3818 3598 3838 3601
rect 3842 3598 3902 3601
rect 3906 3598 4134 3601
rect 4138 3598 4606 3601
rect 4690 3598 4702 3601
rect 4706 3598 5150 3601
rect 2230 3592 2233 3598
rect 2294 3592 2297 3598
rect 490 3588 598 3591
rect 650 3588 1006 3591
rect 1242 3588 1278 3591
rect 1282 3588 1758 3591
rect 1842 3588 1846 3591
rect 1930 3588 1958 3591
rect 1970 3588 1982 3591
rect 2330 3588 2342 3591
rect 2346 3588 2382 3591
rect 2386 3588 2598 3591
rect 2830 3588 2990 3591
rect 3026 3588 3038 3591
rect 3042 3588 3126 3591
rect 3242 3588 3254 3591
rect 3306 3588 3510 3591
rect 3514 3588 3830 3591
rect 3962 3588 4022 3591
rect 4050 3588 4094 3591
rect 4098 3588 4214 3591
rect 4298 3588 4310 3591
rect 4314 3588 4390 3591
rect 4394 3588 4598 3591
rect 4802 3588 4870 3591
rect 4874 3588 4942 3591
rect 458 3578 726 3581
rect 730 3578 798 3581
rect 1026 3578 1142 3581
rect 1146 3578 1302 3581
rect 1314 3578 2606 3581
rect 2710 3581 2713 3588
rect 2830 3582 2833 3588
rect 2698 3578 2713 3581
rect 2730 3578 2830 3581
rect 2890 3578 2974 3581
rect 2978 3578 3006 3581
rect 3042 3578 3574 3581
rect 3578 3578 3662 3581
rect 3722 3578 4422 3581
rect 4602 3578 4894 3581
rect 4898 3578 4902 3581
rect 318 3571 321 3578
rect 298 3568 321 3571
rect 386 3568 446 3571
rect 514 3568 654 3571
rect 898 3568 918 3571
rect 1134 3568 1142 3571
rect 1146 3568 1182 3571
rect 1350 3568 1358 3571
rect 1362 3568 1382 3571
rect 1386 3568 1422 3571
rect 1454 3568 1462 3571
rect 1466 3568 1486 3571
rect 1490 3568 1606 3571
rect 1874 3568 1926 3571
rect 1970 3568 2001 3571
rect 2114 3568 2174 3571
rect 2314 3568 2398 3571
rect 2426 3568 2462 3571
rect 2466 3568 2582 3571
rect 2586 3568 2734 3571
rect 2738 3568 2790 3571
rect 2794 3568 2838 3571
rect 2842 3568 2934 3571
rect 2938 3568 2974 3571
rect 2978 3568 3190 3571
rect 3226 3568 3289 3571
rect 3498 3568 3502 3571
rect 3962 3568 4054 3571
rect 4082 3568 4118 3571
rect 4210 3568 4222 3571
rect 4426 3568 4430 3571
rect 4450 3568 4510 3571
rect 4546 3568 4582 3571
rect 4730 3568 4750 3571
rect 266 3558 302 3561
rect 306 3558 326 3561
rect 362 3558 406 3561
rect 426 3558 430 3561
rect 626 3558 726 3561
rect 878 3561 881 3568
rect 738 3558 881 3561
rect 922 3558 926 3561
rect 1074 3558 1134 3561
rect 1138 3558 1166 3561
rect 1250 3558 1310 3561
rect 1622 3561 1625 3568
rect 1322 3558 1625 3561
rect 1682 3558 1694 3561
rect 1814 3561 1817 3568
rect 1998 3562 2001 3568
rect 3286 3562 3289 3568
rect 1778 3558 1817 3561
rect 1906 3558 1982 3561
rect 2134 3558 2142 3561
rect 2194 3558 2958 3561
rect 2962 3558 3126 3561
rect 3154 3558 3273 3561
rect 3330 3558 3342 3561
rect 3442 3558 3478 3561
rect 3502 3561 3505 3568
rect 3502 3558 3526 3561
rect 3746 3558 3750 3561
rect 3902 3561 3905 3568
rect 3866 3558 3905 3561
rect 3914 3558 3918 3561
rect 4182 3561 4185 3568
rect 3946 3558 4073 3561
rect 4182 3558 4302 3561
rect 4382 3561 4385 3568
rect 4382 3558 4470 3561
rect 4514 3558 4614 3561
rect 4626 3558 4630 3561
rect 4710 3561 4713 3568
rect 4674 3558 4713 3561
rect 4758 3561 4761 3568
rect 4758 3558 4846 3561
rect 4926 3561 4929 3568
rect 4926 3558 5014 3561
rect -26 3551 -22 3552
rect -26 3548 6 3551
rect 154 3548 182 3551
rect 198 3551 201 3558
rect 1246 3552 1249 3558
rect 3270 3552 3273 3558
rect 198 3548 286 3551
rect 402 3548 582 3551
rect 586 3548 606 3551
rect 610 3548 614 3551
rect 682 3548 686 3551
rect 810 3548 830 3551
rect 834 3548 838 3551
rect 890 3548 902 3551
rect 938 3548 1054 3551
rect 1058 3548 1166 3551
rect 1322 3548 1374 3551
rect 1394 3548 1486 3551
rect 1490 3548 1590 3551
rect 1626 3548 1630 3551
rect 1690 3548 1790 3551
rect 1794 3548 1926 3551
rect 1962 3548 2030 3551
rect 2042 3548 2046 3551
rect 2058 3548 2062 3551
rect 2162 3548 2230 3551
rect 2338 3548 2374 3551
rect 2394 3548 2414 3551
rect 2442 3548 2446 3551
rect 2626 3548 2662 3551
rect 2698 3548 2766 3551
rect 358 3542 361 3548
rect 162 3538 270 3541
rect 402 3538 414 3541
rect 498 3538 582 3541
rect 610 3538 846 3541
rect 850 3538 982 3541
rect 1042 3538 2190 3541
rect 2218 3538 2230 3541
rect 2286 3541 2289 3548
rect 2414 3542 2417 3548
rect 2866 3548 2926 3551
rect 3034 3548 3054 3551
rect 3082 3548 3086 3551
rect 3306 3548 3337 3551
rect 3418 3548 3454 3551
rect 3510 3548 3598 3551
rect 3634 3548 3742 3551
rect 3746 3548 3838 3551
rect 3914 3548 3926 3551
rect 3934 3551 3937 3558
rect 3934 3548 4046 3551
rect 4070 3551 4073 3558
rect 5054 3552 5057 3558
rect 4070 3548 4134 3551
rect 4138 3548 4158 3551
rect 4162 3548 4174 3551
rect 4362 3548 4390 3551
rect 4394 3548 4406 3551
rect 4514 3548 4518 3551
rect 4538 3548 4750 3551
rect 4906 3548 4926 3551
rect 3334 3542 3337 3548
rect 3478 3542 3481 3548
rect 3510 3542 3513 3548
rect 2234 3538 2289 3541
rect 2362 3538 2366 3541
rect 2474 3538 2478 3541
rect 2514 3538 2638 3541
rect 2666 3538 2886 3541
rect 3010 3538 3038 3541
rect 3050 3538 3070 3541
rect 3346 3538 3454 3541
rect 3522 3538 3686 3541
rect 3786 3538 3790 3541
rect 3894 3541 3897 3548
rect 3794 3538 3897 3541
rect 4210 3538 4230 3541
rect 4342 3541 4345 3548
rect 4314 3538 4345 3541
rect 4494 3541 4497 3548
rect 4886 3542 4889 3548
rect 4494 3538 4502 3541
rect 4506 3538 4510 3541
rect 4522 3538 4574 3541
rect 4762 3538 4854 3541
rect 5098 3538 5110 3541
rect 5154 3538 5158 3541
rect 270 3532 273 3538
rect 478 3532 481 3538
rect 170 3528 198 3531
rect 530 3528 598 3531
rect 618 3528 638 3531
rect 802 3528 822 3531
rect 990 3531 993 3538
rect 3750 3532 3753 3538
rect 874 3528 993 3531
rect 1122 3528 1126 3531
rect 1130 3528 1470 3531
rect 1482 3528 1494 3531
rect 1594 3528 1686 3531
rect 1714 3528 1718 3531
rect 1722 3528 1838 3531
rect 1866 3528 1902 3531
rect 1906 3528 1958 3531
rect 1970 3528 2174 3531
rect 2178 3528 2486 3531
rect 2514 3528 2550 3531
rect 2570 3528 2633 3531
rect 2650 3528 2657 3531
rect 2674 3528 2830 3531
rect 2834 3528 2862 3531
rect 2866 3528 2942 3531
rect 3130 3528 3134 3531
rect 3266 3528 3318 3531
rect 3410 3528 3414 3531
rect 3434 3528 3438 3531
rect 3442 3528 3534 3531
rect 3546 3528 3694 3531
rect 3906 3528 3942 3531
rect 3954 3528 3974 3531
rect 4002 3528 4094 3531
rect 4122 3528 4142 3531
rect 4146 3528 4214 3531
rect 4394 3528 4534 3531
rect 4738 3528 4934 3531
rect 5154 3528 5166 3531
rect 178 3518 278 3521
rect 370 3518 422 3521
rect 514 3518 566 3521
rect 570 3518 598 3521
rect 638 3521 641 3528
rect 2630 3522 2633 3528
rect 2654 3522 2657 3528
rect 638 3518 910 3521
rect 946 3518 974 3521
rect 978 3518 1022 3521
rect 1042 3518 1126 3521
rect 1274 3518 1302 3521
rect 1314 3518 1350 3521
rect 1434 3518 1438 3521
rect 1458 3518 1550 3521
rect 1778 3518 1814 3521
rect 1818 3518 1974 3521
rect 2002 3518 2030 3521
rect 2170 3518 2310 3521
rect 2378 3518 2430 3521
rect 2538 3518 2550 3521
rect 2714 3518 2870 3521
rect 2946 3518 3150 3521
rect 3170 3518 3310 3521
rect 3354 3518 3382 3521
rect 3450 3518 3950 3521
rect 3954 3518 3982 3521
rect 3986 3518 4086 3521
rect 4110 3521 4113 3528
rect 4090 3518 4142 3521
rect 4402 3518 4526 3521
rect 4530 3518 4542 3521
rect 4570 3518 4598 3521
rect 4610 3518 4710 3521
rect 4714 3518 4966 3521
rect 4970 3518 5078 3521
rect 2094 3512 2097 3518
rect 10 3508 454 3511
rect 458 3508 542 3511
rect 546 3508 646 3511
rect 794 3508 854 3511
rect 866 3508 990 3511
rect 1098 3508 1118 3511
rect 1122 3508 1270 3511
rect 1338 3508 1462 3511
rect 1514 3508 1686 3511
rect 1858 3508 2014 3511
rect 2482 3508 2550 3511
rect 2674 3508 2862 3511
rect 2866 3508 2974 3511
rect 2986 3508 3022 3511
rect 3266 3508 3422 3511
rect 3578 3508 3670 3511
rect 3674 3508 3694 3511
rect 3810 3508 3814 3511
rect 3970 3508 3998 3511
rect 4522 3508 4750 3511
rect 4754 3508 4774 3511
rect 130 3498 142 3501
rect 146 3498 222 3501
rect 386 3498 470 3501
rect 646 3501 649 3508
rect 1048 3503 1050 3507
rect 1054 3503 1057 3507
rect 1062 3503 1064 3507
rect 2072 3503 2074 3507
rect 2078 3503 2081 3507
rect 2086 3503 2088 3507
rect 3096 3503 3098 3507
rect 3102 3503 3105 3507
rect 3110 3503 3112 3507
rect 4112 3503 4114 3507
rect 4118 3503 4121 3507
rect 4126 3503 4128 3507
rect 646 3498 950 3501
rect 954 3498 1038 3501
rect 1194 3498 1270 3501
rect 1298 3498 1334 3501
rect 1394 3498 1414 3501
rect 1426 3498 1446 3501
rect 1506 3498 1814 3501
rect 2162 3498 2278 3501
rect 2282 3498 2390 3501
rect 2450 3498 2678 3501
rect 2826 3498 2894 3501
rect 3210 3498 3262 3501
rect 3298 3498 3710 3501
rect 3714 3498 3750 3501
rect 3770 3498 3902 3501
rect 3970 3498 4102 3501
rect 4578 3498 4590 3501
rect 4930 3498 4982 3501
rect 5130 3498 5150 3501
rect 114 3488 193 3491
rect 190 3482 193 3488
rect 238 3488 646 3491
rect 850 3488 942 3491
rect 986 3488 1046 3491
rect 1258 3488 1286 3491
rect 1314 3488 1358 3491
rect 1398 3488 1406 3491
rect 1410 3488 1582 3491
rect 1698 3488 1886 3491
rect 1954 3488 2038 3491
rect 2066 3488 2166 3491
rect 2354 3488 2470 3491
rect 2474 3488 2534 3491
rect 2618 3488 2622 3491
rect 2634 3488 2710 3491
rect 2818 3488 3286 3491
rect 3298 3488 3438 3491
rect 3666 3488 3678 3491
rect 4426 3488 4470 3491
rect 4694 3491 4697 3498
rect 4610 3488 4697 3491
rect 5066 3488 5118 3491
rect 238 3482 241 3488
rect 170 3478 174 3481
rect 226 3478 230 3481
rect 250 3478 278 3481
rect 294 3478 326 3481
rect 418 3478 585 3481
rect 642 3478 774 3481
rect 930 3478 1238 3481
rect 1242 3478 1358 3481
rect 1378 3478 1382 3481
rect 1386 3478 1502 3481
rect 1602 3478 1606 3481
rect 1682 3478 2654 3481
rect 2730 3478 2790 3481
rect 2946 3478 3046 3481
rect 3106 3478 3110 3481
rect 3130 3478 3406 3481
rect 3458 3478 3534 3481
rect 3546 3478 3582 3481
rect 3642 3478 3766 3481
rect 3826 3478 3870 3481
rect 3898 3478 3910 3481
rect 3994 3478 4358 3481
rect 4442 3478 4622 3481
rect 4674 3478 4782 3481
rect 4786 3478 4798 3481
rect 5162 3478 5190 3481
rect 154 3468 158 3471
rect 162 3468 214 3471
rect 226 3468 230 3471
rect 294 3471 297 3478
rect 234 3468 297 3471
rect 306 3468 390 3471
rect 450 3468 454 3471
rect 466 3468 494 3471
rect 582 3471 585 3478
rect 582 3468 1334 3471
rect 1362 3468 1366 3471
rect 1410 3468 1414 3471
rect 1434 3468 1990 3471
rect 1994 3468 2006 3471
rect 2018 3468 2022 3471
rect 2026 3468 2062 3471
rect 2090 3468 2118 3471
rect 2122 3468 2334 3471
rect 2530 3468 2614 3471
rect 2618 3468 2630 3471
rect 2674 3468 2678 3471
rect 2754 3468 2894 3471
rect 3058 3468 3134 3471
rect 3362 3468 3414 3471
rect 3426 3468 3430 3471
rect 3538 3468 3574 3471
rect 3626 3468 3662 3471
rect 3782 3471 3785 3478
rect 3674 3468 3785 3471
rect 3810 3468 3822 3471
rect 3890 3468 3894 3471
rect 4098 3468 4153 3471
rect 4202 3468 4206 3471
rect 4362 3468 4398 3471
rect 4458 3468 4462 3471
rect 4610 3468 4694 3471
rect 5030 3468 5086 3471
rect 5138 3468 5150 3471
rect 70 3461 73 3468
rect 70 3458 110 3461
rect 386 3458 398 3461
rect 442 3458 534 3461
rect 674 3458 846 3461
rect 866 3458 870 3461
rect 962 3458 982 3461
rect 994 3458 998 3461
rect 1042 3458 1046 3461
rect 1066 3458 1246 3461
rect 1266 3458 1302 3461
rect 1306 3458 1310 3461
rect 1314 3458 1438 3461
rect 1442 3458 1454 3461
rect 1506 3458 1550 3461
rect 1610 3458 1630 3461
rect 1878 3458 1934 3461
rect 1986 3458 1990 3461
rect 2002 3458 2014 3461
rect 2018 3458 2046 3461
rect 2050 3458 2158 3461
rect 2226 3458 2302 3461
rect 2454 3461 2457 3468
rect 2402 3459 2457 3461
rect 2398 3458 2457 3459
rect 2494 3458 2526 3461
rect 2538 3458 2678 3461
rect 2874 3458 2878 3461
rect 2994 3458 3078 3461
rect 3154 3458 3158 3461
rect 3186 3458 3190 3461
rect 3230 3458 3238 3461
rect 3270 3461 3273 3468
rect 3242 3458 3273 3461
rect 3362 3458 3382 3461
rect 3406 3458 3478 3461
rect 3498 3458 3926 3461
rect 3930 3458 4014 3461
rect 4150 3462 4153 3468
rect 4718 3462 4721 3468
rect 5030 3462 5033 3468
rect 4034 3459 4094 3461
rect 4030 3458 4094 3459
rect 4202 3458 4206 3461
rect 4338 3458 4382 3461
rect 4386 3458 4430 3461
rect 4474 3458 4670 3461
rect 4730 3458 4750 3461
rect 4770 3458 4846 3461
rect 4906 3458 4910 3461
rect 4914 3458 4918 3461
rect 262 3452 265 3458
rect 398 3452 401 3458
rect 958 3452 961 3458
rect 1694 3452 1697 3458
rect 1734 3452 1737 3458
rect 1838 3452 1841 3458
rect 1878 3452 1881 3458
rect 2494 3452 2497 3458
rect 3406 3452 3409 3458
rect 10 3448 134 3451
rect 138 3448 230 3451
rect 410 3448 566 3451
rect 602 3448 614 3451
rect 682 3448 686 3451
rect 746 3448 750 3451
rect 754 3448 806 3451
rect 834 3448 838 3451
rect 874 3448 902 3451
rect 1322 3448 1326 3451
rect 1346 3448 1382 3451
rect 1394 3448 1398 3451
rect 1450 3448 1502 3451
rect 1506 3448 1614 3451
rect 1618 3448 1678 3451
rect 1890 3448 2038 3451
rect 2082 3448 2086 3451
rect 2102 3448 2110 3451
rect 2114 3448 2142 3451
rect 2178 3448 2238 3451
rect 2274 3448 2318 3451
rect 2378 3448 2446 3451
rect 2506 3448 2614 3451
rect 2650 3448 2774 3451
rect 2890 3448 2926 3451
rect 3002 3448 3254 3451
rect 3290 3448 3318 3451
rect 3346 3448 3369 3451
rect 3394 3448 3398 3451
rect 3438 3448 3590 3451
rect 3594 3448 3638 3451
rect 3666 3448 3742 3451
rect 3770 3448 3798 3451
rect 3850 3448 3910 3451
rect 3914 3448 3921 3451
rect 3930 3448 3974 3451
rect 4086 3448 4094 3451
rect 4198 3451 4201 3458
rect 4122 3448 4201 3451
rect 4410 3448 4446 3451
rect 4570 3448 4673 3451
rect 4746 3448 4758 3451
rect 4918 3448 5006 3451
rect 5162 3448 5174 3451
rect 106 3438 153 3441
rect 198 3438 206 3441
rect 210 3438 246 3441
rect 266 3438 422 3441
rect 578 3438 614 3441
rect 658 3438 678 3441
rect 690 3438 1030 3441
rect 1114 3438 1134 3441
rect 1342 3441 1345 3448
rect 1138 3438 1345 3441
rect 1354 3438 1366 3441
rect 1430 3441 1433 3448
rect 1386 3438 1433 3441
rect 1490 3438 1678 3441
rect 1706 3438 1942 3441
rect 1946 3438 2014 3441
rect 2054 3441 2057 3448
rect 2034 3438 2057 3441
rect 2066 3438 2134 3441
rect 2162 3438 2286 3441
rect 2290 3438 2334 3441
rect 2338 3438 2438 3441
rect 2442 3438 2494 3441
rect 2570 3438 2622 3441
rect 2630 3441 2633 3448
rect 2630 3438 2654 3441
rect 2670 3438 2710 3441
rect 3050 3438 3070 3441
rect 3074 3438 3078 3441
rect 3138 3438 3358 3441
rect 3366 3441 3369 3448
rect 3438 3442 3441 3448
rect 4086 3442 4089 3448
rect 3366 3438 3433 3441
rect 3450 3438 3454 3441
rect 3658 3438 3662 3441
rect 3786 3438 3790 3441
rect 3914 3438 3918 3441
rect 3946 3438 3990 3441
rect 4146 3438 4166 3441
rect 4198 3438 4254 3441
rect 4370 3438 4558 3441
rect 4562 3438 4662 3441
rect 4670 3441 4673 3448
rect 4918 3442 4921 3448
rect 4670 3438 4798 3441
rect 4938 3438 5182 3441
rect 150 3432 153 3438
rect 2670 3432 2673 3438
rect 2782 3432 2785 3438
rect 162 3428 214 3431
rect 218 3428 278 3431
rect 282 3428 318 3431
rect 654 3428 734 3431
rect 1234 3428 1350 3431
rect 1362 3428 1454 3431
rect 1482 3428 1654 3431
rect 1690 3428 1702 3431
rect 1866 3428 2030 3431
rect 2034 3428 2094 3431
rect 2122 3428 2654 3431
rect 3042 3428 3094 3431
rect 3178 3428 3374 3431
rect 3378 3428 3422 3431
rect 3430 3431 3433 3438
rect 3462 3431 3465 3438
rect 4174 3432 4177 3438
rect 4198 3432 4201 3438
rect 3430 3428 3465 3431
rect 3538 3428 3558 3431
rect 3562 3428 4054 3431
rect 4322 3428 4622 3431
rect 4762 3428 5166 3431
rect 654 3422 657 3428
rect 122 3418 238 3421
rect 1162 3418 1414 3421
rect 1418 3418 1518 3421
rect 1550 3418 1710 3421
rect 1726 3421 1729 3428
rect 1726 3418 1833 3421
rect 1842 3418 1998 3421
rect 2450 3418 2470 3421
rect 2506 3418 2838 3421
rect 2882 3418 2910 3421
rect 2914 3418 2942 3421
rect 3010 3418 3262 3421
rect 3266 3418 3350 3421
rect 3586 3418 3902 3421
rect 3906 3418 4310 3421
rect 562 3408 1110 3411
rect 1146 3408 1198 3411
rect 1550 3411 1553 3418
rect 1290 3408 1553 3411
rect 1642 3408 1782 3411
rect 1830 3411 1833 3418
rect 1830 3408 1918 3411
rect 2874 3408 2902 3411
rect 2906 3408 3054 3411
rect 3250 3408 3398 3411
rect 3666 3408 3830 3411
rect 3922 3408 3966 3411
rect 3978 3408 4006 3411
rect 4010 3408 4070 3411
rect 4178 3408 4214 3411
rect 4226 3408 4438 3411
rect 536 3403 538 3407
rect 542 3403 545 3407
rect 550 3403 552 3407
rect 1560 3403 1562 3407
rect 1566 3403 1569 3407
rect 1574 3403 1576 3407
rect 2584 3403 2586 3407
rect 2590 3403 2593 3407
rect 2598 3403 2600 3407
rect 3608 3403 3610 3407
rect 3614 3403 3617 3407
rect 3622 3403 3624 3407
rect 4632 3403 4634 3407
rect 4638 3403 4641 3407
rect 4646 3403 4648 3407
rect 730 3398 902 3401
rect 970 3398 974 3401
rect 986 3398 1174 3401
rect 1322 3398 1390 3401
rect 1434 3398 1534 3401
rect 1602 3398 1630 3401
rect 1778 3398 1974 3401
rect 2162 3398 2494 3401
rect 2554 3398 2574 3401
rect 3146 3398 3518 3401
rect 3650 3398 3830 3401
rect 4106 3398 4390 3401
rect 410 3388 838 3391
rect 850 3388 1542 3391
rect 1546 3388 2606 3391
rect 2610 3388 2774 3391
rect 2826 3388 3302 3391
rect 3322 3388 3518 3391
rect 3722 3388 3782 3391
rect 4338 3388 4358 3391
rect 4618 3388 5001 3391
rect 4998 3382 5001 3388
rect 234 3378 262 3381
rect 698 3378 710 3381
rect 714 3378 742 3381
rect 834 3378 878 3381
rect 1026 3378 1142 3381
rect 1158 3378 1414 3381
rect 1466 3378 1470 3381
rect 1530 3378 1550 3381
rect 1578 3378 1662 3381
rect 1666 3378 1678 3381
rect 1754 3378 1782 3381
rect 1786 3378 1830 3381
rect 2114 3378 2958 3381
rect 2962 3378 2966 3381
rect 3090 3378 3166 3381
rect 3386 3378 3614 3381
rect 3642 3378 3878 3381
rect 3946 3378 3974 3381
rect 4210 3378 4262 3381
rect 4642 3378 4726 3381
rect 4938 3378 4950 3381
rect 5174 3381 5177 3388
rect 5002 3378 5177 3381
rect 394 3368 406 3371
rect 498 3368 510 3371
rect 514 3368 542 3371
rect 554 3368 806 3371
rect 866 3368 870 3371
rect 958 3371 961 3378
rect 958 3368 982 3371
rect 1158 3371 1161 3378
rect 1090 3368 1161 3371
rect 1258 3368 1294 3371
rect 1410 3368 1582 3371
rect 1642 3368 1830 3371
rect 1834 3368 1841 3371
rect 2038 3371 2041 3378
rect 1954 3368 2041 3371
rect 2162 3368 2206 3371
rect 2302 3368 2422 3371
rect 2546 3368 2558 3371
rect 2618 3368 2782 3371
rect 2826 3368 2854 3371
rect 2930 3368 2990 3371
rect 3050 3368 3094 3371
rect 3210 3368 3278 3371
rect 3310 3371 3313 3378
rect 3310 3368 3374 3371
rect 3418 3368 3478 3371
rect 3546 3368 3566 3371
rect 3602 3368 3702 3371
rect 3970 3368 3974 3371
rect 4062 3368 4070 3371
rect 4074 3368 4174 3371
rect 4178 3368 4350 3371
rect 4634 3368 4654 3371
rect 4914 3368 4998 3371
rect 5170 3368 5174 3371
rect 238 3361 241 3368
rect 1158 3362 1161 3368
rect 2302 3362 2305 3368
rect 178 3358 241 3361
rect 330 3358 422 3361
rect 450 3358 510 3361
rect 514 3358 521 3361
rect 530 3358 558 3361
rect 666 3358 782 3361
rect 786 3358 878 3361
rect 882 3358 998 3361
rect 1026 3358 1102 3361
rect 1106 3358 1113 3361
rect 1130 3358 1150 3361
rect 1282 3358 1318 3361
rect 1362 3358 1398 3361
rect 1410 3358 1494 3361
rect 1506 3358 1678 3361
rect 1786 3358 1854 3361
rect 2010 3358 2022 3361
rect 2058 3358 2062 3361
rect 2194 3358 2214 3361
rect 2326 3358 2334 3361
rect 2338 3358 2366 3361
rect 2458 3358 2462 3361
rect 2518 3361 2521 3368
rect 2534 3361 2537 3368
rect 2518 3358 2537 3361
rect 2554 3358 2614 3361
rect 2762 3358 2838 3361
rect 2866 3358 2886 3361
rect 3090 3358 3278 3361
rect 3282 3358 3326 3361
rect 3522 3358 3550 3361
rect 3582 3361 3585 3368
rect 3578 3358 3585 3361
rect 3714 3358 4038 3361
rect 4042 3358 4086 3361
rect 4170 3358 4190 3361
rect 4402 3358 4406 3361
rect 4430 3361 4433 3368
rect 4430 3358 4502 3361
rect 4558 3361 4561 3368
rect 4558 3358 4566 3361
rect 4618 3358 4654 3361
rect 4762 3358 4766 3361
rect 4786 3358 4790 3361
rect 4846 3361 4849 3368
rect 4910 3361 4913 3368
rect 4846 3358 4913 3361
rect 4922 3358 4934 3361
rect 4958 3358 4966 3361
rect 4986 3358 5110 3361
rect 5130 3358 5142 3361
rect 5162 3358 5166 3361
rect 98 3348 230 3351
rect 426 3348 526 3351
rect 530 3348 598 3351
rect 650 3348 686 3351
rect 726 3348 798 3351
rect 898 3348 926 3351
rect 1074 3348 1102 3351
rect 1106 3348 1422 3351
rect 1434 3348 1734 3351
rect 1798 3348 1806 3351
rect 1810 3348 1870 3351
rect 1906 3348 2006 3351
rect 2010 3348 2174 3351
rect 2178 3348 2230 3351
rect 2270 3351 2273 3358
rect 2270 3348 2278 3351
rect 2354 3348 2526 3351
rect 2538 3348 2670 3351
rect 2682 3348 2686 3351
rect 2738 3348 2830 3351
rect 2938 3348 2974 3351
rect 3090 3348 3126 3351
rect 3138 3348 3262 3351
rect 3266 3348 3574 3351
rect 3626 3348 3630 3351
rect 3682 3348 3710 3351
rect 3722 3348 3726 3351
rect 3738 3348 3742 3351
rect 3970 3348 3974 3351
rect 4146 3348 4166 3351
rect 4186 3348 4246 3351
rect 4258 3348 4294 3351
rect 4386 3348 4390 3351
rect 4442 3348 4558 3351
rect 4562 3348 4574 3351
rect 4594 3348 4598 3351
rect 4690 3348 4718 3351
rect 4722 3348 4734 3351
rect 4738 3348 4822 3351
rect 4826 3348 4846 3351
rect 4874 3348 4886 3351
rect 4922 3348 4950 3351
rect 5002 3348 5006 3351
rect 5058 3348 5062 3351
rect 98 3338 118 3341
rect 398 3341 401 3348
rect 726 3342 729 3348
rect 2334 3342 2337 3348
rect 306 3338 401 3341
rect 522 3338 526 3341
rect 578 3338 646 3341
rect 746 3338 750 3341
rect 862 3338 1070 3341
rect 1114 3338 1126 3341
rect 1170 3338 1182 3341
rect 1302 3338 1358 3341
rect 1458 3338 1462 3341
rect 1498 3338 1502 3341
rect 1530 3338 1606 3341
rect 1714 3338 1742 3341
rect 1754 3338 1934 3341
rect 2034 3338 2038 3341
rect 2074 3338 2102 3341
rect 2106 3338 2198 3341
rect 2218 3338 2262 3341
rect 2266 3338 2286 3341
rect 2458 3338 2630 3341
rect 2818 3338 2822 3341
rect 2906 3338 2910 3341
rect 3078 3341 3081 3348
rect 3838 3342 3841 3348
rect 5134 3342 5137 3348
rect 2978 3338 3081 3341
rect 3154 3338 3254 3341
rect 3314 3338 3358 3341
rect 3362 3338 3454 3341
rect 3458 3338 3494 3341
rect 3586 3338 3782 3341
rect 3866 3338 3886 3341
rect 3930 3338 3958 3341
rect 3978 3338 4030 3341
rect 4074 3338 4078 3341
rect 4098 3338 4222 3341
rect 4226 3338 4246 3341
rect 4266 3338 4366 3341
rect 4370 3338 4702 3341
rect 4794 3338 4822 3341
rect 4898 3338 4958 3341
rect 4962 3338 5078 3341
rect 5090 3338 5102 3341
rect 862 3332 865 3338
rect 1302 3332 1305 3338
rect 2014 3332 2017 3338
rect 2454 3332 2457 3338
rect 170 3328 230 3331
rect 242 3328 342 3331
rect 346 3328 422 3331
rect 498 3328 670 3331
rect 682 3328 710 3331
rect 922 3328 966 3331
rect 986 3328 1206 3331
rect 1218 3328 1230 3331
rect 1234 3328 1270 3331
rect 1426 3328 1510 3331
rect 1690 3328 1766 3331
rect 2018 3328 2278 3331
rect 2518 3328 2526 3331
rect 2530 3328 2550 3331
rect 2562 3328 2566 3331
rect 2882 3328 3030 3331
rect 3046 3328 3062 3331
rect 3082 3328 3222 3331
rect 3354 3328 3550 3331
rect 3566 3331 3569 3338
rect 4750 3332 4753 3338
rect 3566 3328 3654 3331
rect 3738 3328 3742 3331
rect 3826 3328 3902 3331
rect 3910 3328 4062 3331
rect 4162 3328 4190 3331
rect 4250 3328 4302 3331
rect 4386 3328 4398 3331
rect 4530 3328 4566 3331
rect 4578 3328 4665 3331
rect 4826 3328 5046 3331
rect 5074 3328 5078 3331
rect 5106 3328 5158 3331
rect 3046 3322 3049 3328
rect 162 3318 286 3321
rect 290 3318 382 3321
rect 386 3318 478 3321
rect 482 3318 582 3321
rect 586 3318 910 3321
rect 914 3318 982 3321
rect 1074 3318 1238 3321
rect 1362 3318 1446 3321
rect 1474 3318 1542 3321
rect 2802 3318 2886 3321
rect 3146 3318 3150 3321
rect 3274 3318 3590 3321
rect 3766 3321 3769 3328
rect 3594 3318 3769 3321
rect 3910 3322 3913 3328
rect 4150 3322 4153 3328
rect 4662 3322 4665 3328
rect 4106 3318 4118 3321
rect 4162 3318 4198 3321
rect 4370 3318 4582 3321
rect 4594 3318 4614 3321
rect 5146 3318 5158 3321
rect 4918 3312 4921 3318
rect 82 3308 398 3311
rect 658 3308 686 3311
rect 1258 3308 1430 3311
rect 1730 3308 1766 3311
rect 1770 3308 1806 3311
rect 1818 3308 1822 3311
rect 1826 3308 2062 3311
rect 2122 3308 2134 3311
rect 2138 3308 2214 3311
rect 2234 3308 2366 3311
rect 2826 3308 3078 3311
rect 3402 3308 3406 3311
rect 3554 3308 3558 3311
rect 3722 3308 3806 3311
rect 3810 3308 3846 3311
rect 4290 3308 4446 3311
rect 4594 3308 4598 3311
rect 4602 3308 4638 3311
rect 4706 3308 4766 3311
rect 1048 3303 1050 3307
rect 1054 3303 1057 3307
rect 1062 3303 1064 3307
rect 2072 3303 2074 3307
rect 2078 3303 2081 3307
rect 2086 3303 2088 3307
rect 3096 3303 3098 3307
rect 3102 3303 3105 3307
rect 3110 3303 3112 3307
rect 4112 3303 4114 3307
rect 4118 3303 4121 3307
rect 4126 3303 4128 3307
rect 18 3298 78 3301
rect 130 3298 222 3301
rect 258 3298 318 3301
rect 322 3298 390 3301
rect 426 3298 606 3301
rect 610 3298 630 3301
rect 634 3298 726 3301
rect 938 3298 974 3301
rect 1074 3298 2038 3301
rect 2106 3298 2166 3301
rect 2242 3298 2286 3301
rect 2402 3298 2438 3301
rect 2466 3298 2678 3301
rect 2682 3298 2790 3301
rect 2866 3298 2926 3301
rect 3010 3298 3038 3301
rect 3050 3298 3086 3301
rect 3314 3298 3318 3301
rect 3322 3298 3326 3301
rect 3338 3298 3398 3301
rect 3546 3298 3574 3301
rect 3658 3298 3790 3301
rect 3794 3298 3990 3301
rect 4138 3298 4246 3301
rect 4266 3298 4398 3301
rect 4434 3298 4438 3301
rect 4490 3298 4542 3301
rect 4746 3298 4870 3301
rect 4874 3298 4974 3301
rect 122 3288 182 3291
rect 214 3288 254 3291
rect 346 3288 414 3291
rect 418 3288 494 3291
rect 498 3288 598 3291
rect 626 3288 686 3291
rect 722 3288 902 3291
rect 954 3288 1118 3291
rect 1122 3288 1134 3291
rect 1178 3288 1254 3291
rect 1274 3288 1478 3291
rect 1506 3288 1598 3291
rect 1698 3288 1710 3291
rect 2282 3288 2326 3291
rect 2330 3288 2478 3291
rect 2498 3288 2550 3291
rect 2554 3288 2566 3291
rect 2570 3288 2713 3291
rect 2754 3288 2774 3291
rect 2794 3288 2910 3291
rect 3034 3288 3270 3291
rect 3378 3288 3406 3291
rect 3490 3288 3614 3291
rect 3770 3288 3774 3291
rect 3778 3288 4038 3291
rect 4042 3288 4046 3291
rect 4186 3288 4214 3291
rect 4766 3288 4854 3291
rect 4866 3288 4974 3291
rect 214 3282 217 3288
rect 286 3281 289 3288
rect 266 3278 289 3281
rect 602 3278 606 3281
rect 626 3278 654 3281
rect 658 3278 870 3281
rect 950 3281 953 3288
rect 874 3278 953 3281
rect 982 3278 1182 3281
rect 1258 3278 1334 3281
rect 1538 3278 1670 3281
rect 1874 3278 1958 3281
rect 2042 3278 2190 3281
rect 2242 3278 2310 3281
rect 2322 3278 2361 3281
rect 2442 3278 2582 3281
rect 2710 3281 2713 3288
rect 2710 3278 3118 3281
rect 3146 3278 3217 3281
rect 3258 3278 3262 3281
rect 3354 3278 3422 3281
rect 3490 3278 3502 3281
rect 3538 3278 3558 3281
rect 3602 3278 3726 3281
rect 4026 3278 4190 3281
rect 4210 3278 4398 3281
rect 4454 3281 4457 3288
rect 4766 3282 4769 3288
rect 4402 3278 4457 3281
rect 4574 3278 4582 3281
rect 4586 3278 4606 3281
rect 4610 3278 4662 3281
rect 4810 3278 4830 3281
rect 4866 3278 4886 3281
rect 4930 3278 4934 3281
rect 134 3271 137 3278
rect 66 3268 137 3271
rect 226 3268 286 3271
rect 298 3268 326 3271
rect 382 3271 385 3278
rect 982 3272 985 3278
rect 2358 3272 2361 3278
rect 3214 3272 3217 3278
rect 3966 3272 3969 3278
rect 382 3268 446 3271
rect 738 3268 774 3271
rect 858 3268 878 3271
rect 930 3268 958 3271
rect 962 3268 966 3271
rect 994 3268 1078 3271
rect 1082 3268 1182 3271
rect 1194 3268 1310 3271
rect 1314 3268 1342 3271
rect 1482 3268 1486 3271
rect 1514 3268 1758 3271
rect 1802 3268 1910 3271
rect 2018 3268 2078 3271
rect 2138 3268 2142 3271
rect 2258 3268 2286 3271
rect 2290 3268 2350 3271
rect 2366 3268 2502 3271
rect 2630 3268 2638 3271
rect 2658 3268 2662 3271
rect 2666 3268 2718 3271
rect 2890 3268 2902 3271
rect 2938 3268 2982 3271
rect 2994 3268 3030 3271
rect 3034 3268 3094 3271
rect 3098 3268 3134 3271
rect 3266 3268 3550 3271
rect 3586 3268 3662 3271
rect 3674 3268 3726 3271
rect 3730 3268 3734 3271
rect 3754 3268 3798 3271
rect 3986 3268 3990 3271
rect 4154 3268 4161 3271
rect 4178 3268 4214 3271
rect 4386 3268 4502 3271
rect 4538 3268 4574 3271
rect 4742 3271 4745 3278
rect 4742 3268 4998 3271
rect 70 3258 110 3261
rect 122 3258 126 3261
rect 170 3258 238 3261
rect 258 3258 329 3261
rect 354 3258 398 3261
rect 614 3261 617 3268
rect 886 3262 889 3268
rect 530 3258 617 3261
rect 674 3258 694 3261
rect 698 3258 702 3261
rect 746 3258 854 3261
rect 1010 3258 1086 3261
rect 1142 3258 1150 3261
rect 1154 3258 1174 3261
rect 1194 3258 1222 3261
rect 1290 3258 1382 3261
rect 1418 3258 1494 3261
rect 1610 3259 1654 3261
rect 1606 3258 1654 3259
rect 1674 3258 1726 3261
rect 1790 3258 1798 3261
rect 1802 3258 1841 3261
rect 1954 3258 1958 3261
rect 2074 3258 2182 3261
rect 2366 3261 2369 3268
rect 2614 3262 2617 3268
rect 2630 3262 2633 3268
rect 2314 3258 2369 3261
rect 2378 3258 2382 3261
rect 2498 3258 2574 3261
rect 2658 3258 2694 3261
rect 2734 3261 2737 3268
rect 2734 3258 2774 3261
rect 2818 3258 2846 3261
rect 2962 3258 2966 3261
rect 3114 3258 3118 3261
rect 3182 3261 3185 3268
rect 3130 3258 3185 3261
rect 3198 3261 3201 3268
rect 3198 3258 3206 3261
rect 3210 3258 3310 3261
rect 3330 3258 3374 3261
rect 3402 3258 3438 3261
rect 3458 3258 3462 3261
rect 3474 3258 3502 3261
rect 3658 3258 3990 3261
rect 3994 3258 3998 3261
rect 4058 3258 4110 3261
rect 4142 3261 4145 3268
rect 4138 3258 4145 3261
rect 4158 3262 4161 3268
rect 4238 3262 4241 3268
rect 4410 3258 4414 3261
rect 4418 3258 4430 3261
rect 4442 3258 4510 3261
rect 4530 3258 4558 3261
rect 4562 3258 4622 3261
rect 4642 3258 4710 3261
rect 4786 3258 4790 3261
rect 4794 3258 4806 3261
rect 4930 3258 5006 3261
rect 5098 3258 5182 3261
rect 6 3252 9 3258
rect 70 3252 73 3258
rect 90 3248 110 3251
rect 326 3251 329 3258
rect 1142 3252 1145 3258
rect 1838 3252 1841 3258
rect 2310 3252 2313 3258
rect 2798 3252 2801 3258
rect 2894 3252 2897 3258
rect 2990 3252 2993 3258
rect 3542 3252 3545 3258
rect 114 3248 313 3251
rect 326 3248 358 3251
rect 666 3248 745 3251
rect 890 3248 918 3251
rect 970 3248 1006 3251
rect 1098 3248 1118 3251
rect 1178 3248 1182 3251
rect 1282 3248 1286 3251
rect 1290 3248 1470 3251
rect 1522 3248 1614 3251
rect 1666 3248 1742 3251
rect 1778 3248 1806 3251
rect 1906 3248 1950 3251
rect 2130 3248 2134 3251
rect 2546 3248 2598 3251
rect 2602 3248 2622 3251
rect 2698 3248 2734 3251
rect 2738 3248 2742 3251
rect 2770 3248 2774 3251
rect 2802 3248 2822 3251
rect 2914 3248 2958 3251
rect 2962 3248 2969 3251
rect 3274 3248 3438 3251
rect 3474 3248 3478 3251
rect 3562 3248 3670 3251
rect 3690 3248 3734 3251
rect 3794 3248 3806 3251
rect 3814 3248 3902 3251
rect 3978 3248 4022 3251
rect 4198 3248 4206 3251
rect 4210 3248 4246 3251
rect 4430 3251 4433 3258
rect 4430 3248 4574 3251
rect 4578 3248 4862 3251
rect 4866 3248 4886 3251
rect 4914 3248 4934 3251
rect 5186 3248 5190 3251
rect 310 3242 313 3248
rect 250 3238 273 3241
rect 314 3238 374 3241
rect 630 3241 633 3248
rect 586 3238 734 3241
rect 742 3241 745 3248
rect 1126 3241 1129 3248
rect 742 3238 1190 3241
rect 1202 3238 1238 3241
rect 1518 3241 1521 3248
rect 1774 3242 1777 3248
rect 1242 3238 1521 3241
rect 1610 3238 1646 3241
rect 1958 3241 1961 3248
rect 1958 3238 1966 3241
rect 1970 3238 2094 3241
rect 2326 3241 2329 3248
rect 3814 3242 3817 3248
rect 2298 3238 2329 3241
rect 2506 3238 2670 3241
rect 2762 3238 2854 3241
rect 3362 3238 3582 3241
rect 4218 3238 4222 3241
rect 4226 3238 4470 3241
rect 4810 3238 4830 3241
rect 4882 3238 4926 3241
rect 270 3232 273 3238
rect 282 3228 374 3231
rect 530 3228 550 3231
rect 706 3228 990 3231
rect 1018 3228 1358 3231
rect 1362 3228 1366 3231
rect 1474 3228 1502 3231
rect 1674 3228 2046 3231
rect 2150 3231 2153 3238
rect 2150 3228 2350 3231
rect 2354 3228 2534 3231
rect 2642 3228 2902 3231
rect 2906 3228 3014 3231
rect 3018 3228 3318 3231
rect 3338 3228 3374 3231
rect 3430 3228 3510 3231
rect 3594 3228 3694 3231
rect 3766 3231 3769 3238
rect 3766 3228 3846 3231
rect 3898 3228 4470 3231
rect 4570 3228 4606 3231
rect 4610 3228 4814 3231
rect 4818 3228 4862 3231
rect 3430 3222 3433 3228
rect 330 3218 670 3221
rect 674 3218 806 3221
rect 810 3218 1758 3221
rect 1946 3218 1982 3221
rect 2514 3218 2750 3221
rect 2754 3218 3398 3221
rect 3530 3218 3718 3221
rect 3754 3218 3934 3221
rect 3938 3218 4142 3221
rect 4234 3218 4254 3221
rect 4258 3218 4310 3221
rect 4442 3218 4446 3221
rect 4554 3218 4782 3221
rect 330 3208 430 3211
rect 458 3208 478 3211
rect 570 3208 934 3211
rect 994 3208 1302 3211
rect 1666 3208 1806 3211
rect 1810 3208 1974 3211
rect 1978 3208 2278 3211
rect 2642 3208 2782 3211
rect 2818 3208 3198 3211
rect 3250 3208 3542 3211
rect 3682 3208 3742 3211
rect 3794 3208 3950 3211
rect 4306 3208 4486 3211
rect 4746 3208 4774 3211
rect 536 3203 538 3207
rect 542 3203 545 3207
rect 550 3203 552 3207
rect 934 3201 937 3208
rect 1560 3203 1562 3207
rect 1566 3203 1569 3207
rect 1574 3203 1576 3207
rect 2584 3203 2586 3207
rect 2590 3203 2593 3207
rect 2598 3203 2600 3207
rect 3608 3203 3610 3207
rect 3614 3203 3617 3207
rect 3622 3203 3624 3207
rect 4632 3203 4634 3207
rect 4638 3203 4641 3207
rect 4646 3203 4648 3207
rect 346 3198 529 3201
rect 934 3198 1094 3201
rect 1114 3198 1198 3201
rect 1202 3198 1486 3201
rect 1618 3198 1686 3201
rect 1706 3198 1902 3201
rect 1906 3198 2214 3201
rect 2218 3198 2270 3201
rect 2434 3198 2486 3201
rect 2610 3198 2718 3201
rect 2778 3198 2854 3201
rect 2954 3198 3086 3201
rect 3090 3198 3214 3201
rect 3346 3198 3390 3201
rect 3698 3198 3814 3201
rect 4178 3198 4190 3201
rect 4690 3198 4838 3201
rect 4890 3198 4966 3201
rect 5098 3198 5110 3201
rect 234 3188 350 3191
rect 526 3191 529 3198
rect 526 3188 798 3191
rect 906 3188 1102 3191
rect 1106 3188 1222 3191
rect 1226 3188 1374 3191
rect 1466 3188 1478 3191
rect 1482 3188 1662 3191
rect 1682 3188 1750 3191
rect 1770 3188 1998 3191
rect 2162 3188 2454 3191
rect 2562 3188 2718 3191
rect 2730 3188 2886 3191
rect 2890 3188 3062 3191
rect 3098 3188 3222 3191
rect 3642 3188 3950 3191
rect 3954 3188 3982 3191
rect 4194 3188 4534 3191
rect 4698 3188 4910 3191
rect 4914 3188 4982 3191
rect 5066 3188 5166 3191
rect 3390 3182 3393 3188
rect 458 3178 902 3181
rect 1058 3178 1118 3181
rect 1138 3178 1145 3181
rect 1162 3178 1222 3181
rect 1278 3178 1286 3181
rect 1290 3178 1318 3181
rect 1538 3178 1638 3181
rect 1642 3178 2102 3181
rect 2226 3178 2318 3181
rect 2330 3178 2550 3181
rect 2826 3178 2910 3181
rect 2922 3178 2942 3181
rect 2986 3178 3046 3181
rect 3050 3178 3094 3181
rect 3238 3178 3246 3181
rect 3250 3178 3278 3181
rect 3426 3178 3566 3181
rect 3698 3178 4038 3181
rect 4162 3178 4310 3181
rect 4706 3178 4846 3181
rect 4954 3178 5094 3181
rect 66 3168 110 3171
rect 342 3171 345 3178
rect 282 3168 345 3171
rect 570 3168 646 3171
rect 866 3168 1302 3171
rect 1498 3168 1798 3171
rect 1914 3168 1990 3171
rect 1994 3168 2126 3171
rect 2130 3168 2150 3171
rect 2154 3168 2230 3171
rect 2322 3168 2366 3171
rect 2442 3168 2446 3171
rect 2522 3168 2606 3171
rect 2618 3168 2638 3171
rect 2806 3171 2809 3178
rect 2794 3168 2809 3171
rect 2842 3168 3070 3171
rect 3074 3168 3694 3171
rect 3758 3168 3766 3171
rect 3770 3168 3790 3171
rect 3794 3168 3822 3171
rect 3834 3168 4198 3171
rect 4918 3171 4921 3178
rect 4730 3168 4921 3171
rect 5146 3168 5150 3171
rect 74 3158 198 3161
rect 330 3158 334 3161
rect 566 3161 569 3168
rect 814 3162 817 3168
rect 4934 3162 4937 3168
rect 474 3158 569 3161
rect 770 3158 774 3161
rect 834 3158 838 3161
rect 842 3158 854 3161
rect 922 3158 926 3161
rect 930 3158 982 3161
rect 1050 3158 1166 3161
rect 1170 3158 1174 3161
rect 1186 3158 1238 3161
rect 1254 3158 1262 3161
rect 1266 3158 1382 3161
rect 1386 3158 1470 3161
rect 1498 3158 1502 3161
rect 1554 3158 1582 3161
rect 1586 3158 1590 3161
rect 1674 3158 1678 3161
rect 1738 3158 1854 3161
rect 1866 3158 1934 3161
rect 1946 3158 1966 3161
rect 2082 3158 2110 3161
rect 2218 3158 2334 3161
rect 2354 3158 2446 3161
rect 2458 3158 2766 3161
rect 2770 3158 2862 3161
rect 2866 3158 3446 3161
rect 3450 3158 3574 3161
rect 3578 3158 3878 3161
rect 4210 3158 4246 3161
rect 4250 3158 4262 3161
rect 4658 3158 4702 3161
rect 4730 3158 4734 3161
rect 4738 3158 4782 3161
rect 4802 3158 4806 3161
rect 4982 3161 4985 3168
rect 4982 3158 5054 3161
rect -26 3151 -22 3152
rect -26 3148 14 3151
rect 354 3148 422 3151
rect 498 3148 526 3151
rect 642 3148 686 3151
rect 722 3148 878 3151
rect 882 3148 950 3151
rect 994 3148 998 3151
rect 1122 3148 1126 3151
rect 1138 3148 1150 3151
rect 1194 3148 1198 3151
rect 1290 3148 1334 3151
rect 1506 3148 1526 3151
rect 1554 3148 1622 3151
rect 1674 3148 1694 3151
rect 1770 3148 1886 3151
rect 1954 3148 1958 3151
rect 2018 3148 2134 3151
rect 2170 3148 2174 3151
rect 2178 3148 2206 3151
rect 2250 3148 2430 3151
rect 2434 3148 2502 3151
rect 2546 3148 2566 3151
rect 2610 3148 2694 3151
rect 2802 3148 2934 3151
rect 2938 3148 2942 3151
rect 2958 3148 3022 3151
rect 3062 3148 3150 3151
rect 3218 3148 3230 3151
rect 3250 3148 3350 3151
rect 3370 3148 3374 3151
rect 3418 3148 3470 3151
rect 3618 3148 3694 3151
rect 3886 3151 3889 3158
rect 3926 3152 3929 3158
rect 3806 3148 3889 3151
rect 4046 3151 4049 3158
rect 3962 3148 4049 3151
rect 4210 3148 4297 3151
rect 4506 3148 4510 3151
rect 4538 3148 4726 3151
rect 4730 3148 4822 3151
rect 4898 3148 4974 3151
rect 4994 3148 4998 3151
rect 5002 3148 5033 3151
rect 5050 3148 5142 3151
rect 102 3142 105 3148
rect 950 3142 953 3148
rect 1726 3142 1729 3148
rect 2958 3142 2961 3148
rect 3062 3142 3065 3148
rect 3806 3142 3809 3148
rect 26 3138 54 3141
rect 122 3138 374 3141
rect 394 3138 406 3141
rect 490 3138 622 3141
rect 690 3138 702 3141
rect 738 3138 742 3141
rect 762 3138 766 3141
rect 810 3138 814 3141
rect 1018 3138 1078 3141
rect 1114 3138 1142 3141
rect 1202 3138 1238 3141
rect 1242 3138 1294 3141
rect 1474 3138 1510 3141
rect 1530 3138 1582 3141
rect 1586 3138 1606 3141
rect 1906 3138 1934 3141
rect 1938 3138 1974 3141
rect 2194 3138 2254 3141
rect 2346 3138 2358 3141
rect 2362 3138 2430 3141
rect 2506 3138 2534 3141
rect 2634 3138 2758 3141
rect 2762 3138 2806 3141
rect 2810 3138 2902 3141
rect 2938 3138 2942 3141
rect 2970 3138 2982 3141
rect 3034 3138 3038 3141
rect 3182 3138 3241 3141
rect 3290 3138 3358 3141
rect 3402 3138 3430 3141
rect 3474 3138 3534 3141
rect 3586 3138 3622 3141
rect 3834 3138 3838 3141
rect 3894 3141 3897 3148
rect 4294 3142 4297 3148
rect 3894 3138 4006 3141
rect 4066 3138 4262 3141
rect 4518 3141 4521 3148
rect 5030 3142 5033 3148
rect 4302 3138 4505 3141
rect 4518 3138 4566 3141
rect 4666 3138 4670 3141
rect 4682 3138 4686 3141
rect 4754 3138 4758 3141
rect 4774 3138 4782 3141
rect 4786 3138 4870 3141
rect 4914 3138 4918 3141
rect 4946 3138 4998 3141
rect 5002 3138 5006 3141
rect 382 3132 385 3138
rect 1686 3132 1689 3138
rect 2094 3132 2097 3138
rect 98 3128 118 3131
rect 394 3128 470 3131
rect 474 3128 582 3131
rect 586 3128 838 3131
rect 898 3128 1014 3131
rect 1034 3128 1182 3131
rect 1194 3128 1286 3131
rect 1290 3128 1326 3131
rect 1386 3128 1422 3131
rect 1442 3128 1446 3131
rect 1450 3128 1526 3131
rect 1834 3128 1846 3131
rect 1850 3128 2014 3131
rect 2550 3131 2553 3138
rect 3182 3132 3185 3138
rect 3238 3132 3241 3138
rect 3462 3132 3465 3138
rect 2550 3128 2654 3131
rect 2682 3128 2790 3131
rect 2882 3128 2966 3131
rect 2970 3128 2974 3131
rect 3002 3128 3142 3131
rect 3242 3128 3294 3131
rect 3298 3128 3406 3131
rect 3430 3128 3438 3131
rect 3442 3128 3446 3131
rect 3634 3128 3665 3131
rect 3738 3128 3742 3131
rect 3746 3128 4054 3131
rect 4098 3128 4102 3131
rect 4138 3128 4174 3131
rect 4302 3131 4305 3138
rect 4290 3128 4305 3131
rect 4502 3131 4505 3138
rect 4502 3128 4718 3131
rect 4762 3128 5078 3131
rect 362 3118 390 3121
rect 482 3118 598 3121
rect 690 3118 710 3121
rect 786 3118 878 3121
rect 898 3118 958 3121
rect 978 3118 982 3121
rect 1002 3118 1118 3121
rect 1122 3118 1270 3121
rect 1402 3118 1406 3121
rect 1418 3118 1534 3121
rect 1750 3121 1753 3128
rect 1714 3118 1753 3121
rect 1834 3118 1910 3121
rect 1946 3118 1974 3121
rect 2066 3118 2126 3121
rect 2186 3118 2294 3121
rect 2298 3118 2302 3121
rect 2374 3121 2377 3128
rect 2374 3118 2518 3121
rect 2546 3118 2638 3121
rect 2642 3118 2798 3121
rect 2874 3118 3134 3121
rect 3314 3118 3358 3121
rect 3662 3121 3665 3128
rect 3662 3118 3734 3121
rect 3738 3118 3806 3121
rect 3818 3118 3878 3121
rect 3882 3118 3974 3121
rect 3978 3118 4158 3121
rect 4494 3121 4497 3128
rect 4494 3118 4518 3121
rect 4866 3118 4950 3121
rect 4994 3118 5014 3121
rect 122 3108 214 3111
rect 410 3108 526 3111
rect 578 3108 614 3111
rect 842 3108 1030 3111
rect 1210 3108 1238 3111
rect 1250 3108 1278 3111
rect 1314 3108 1318 3111
rect 1330 3108 1654 3111
rect 1730 3108 1790 3111
rect 1802 3108 1966 3111
rect 1970 3108 2062 3111
rect 2274 3108 2510 3111
rect 2530 3108 2742 3111
rect 2746 3108 3030 3111
rect 3586 3108 3982 3111
rect 4170 3108 4214 3111
rect 4266 3108 4654 3111
rect 4914 3108 5086 3111
rect 290 3098 414 3101
rect 426 3098 430 3101
rect 434 3098 550 3101
rect 614 3101 617 3108
rect 1048 3103 1050 3107
rect 1054 3103 1057 3107
rect 1062 3103 1064 3107
rect 2072 3103 2074 3107
rect 2078 3103 2081 3107
rect 2086 3103 2088 3107
rect 3096 3103 3098 3107
rect 3102 3103 3105 3107
rect 3110 3103 3112 3107
rect 4112 3103 4114 3107
rect 4118 3103 4121 3107
rect 4126 3103 4128 3107
rect 614 3098 774 3101
rect 778 3098 814 3101
rect 890 3098 894 3101
rect 1178 3098 1598 3101
rect 1602 3098 1782 3101
rect 1866 3098 2054 3101
rect 2458 3098 2486 3101
rect 2490 3098 2662 3101
rect 2722 3098 2742 3101
rect 2758 3098 2774 3101
rect 2778 3098 2830 3101
rect 3018 3098 3070 3101
rect 3186 3098 3478 3101
rect 3690 3098 3846 3101
rect 3850 3098 3870 3101
rect 3906 3098 3942 3101
rect 4218 3098 4230 3101
rect 4426 3098 4462 3101
rect 4466 3098 4470 3101
rect 4514 3098 4678 3101
rect 4682 3098 4718 3101
rect 4778 3098 5142 3101
rect 522 3088 542 3091
rect 706 3088 710 3091
rect 730 3088 758 3091
rect 802 3088 846 3091
rect 890 3088 982 3091
rect 1114 3088 1166 3091
rect 1210 3088 1321 3091
rect 1330 3088 1422 3091
rect 1538 3088 1633 3091
rect 10 3078 126 3081
rect 162 3078 174 3081
rect 178 3078 270 3081
rect 330 3078 390 3081
rect 394 3078 462 3081
rect 506 3078 606 3081
rect 610 3078 630 3081
rect 682 3078 734 3081
rect 738 3078 862 3081
rect 898 3078 942 3081
rect 1146 3078 1278 3081
rect 1318 3081 1321 3088
rect 1630 3082 1633 3088
rect 1658 3088 1678 3091
rect 1750 3088 1846 3091
rect 2266 3088 2574 3091
rect 2758 3091 2761 3098
rect 2578 3088 2761 3091
rect 2778 3088 3062 3091
rect 3082 3088 3310 3091
rect 3362 3088 3446 3091
rect 3498 3088 3822 3091
rect 4242 3088 4270 3091
rect 4290 3088 4838 3091
rect 4842 3088 4870 3091
rect 4890 3088 4894 3091
rect 4898 3088 4942 3091
rect 4978 3088 4990 3091
rect 1318 3078 1358 3081
rect 1402 3078 1430 3081
rect 1482 3078 1486 3081
rect 1546 3078 1606 3081
rect 1610 3078 1622 3081
rect 1638 3081 1641 3088
rect 1750 3082 1753 3088
rect 1638 3078 1654 3081
rect 1706 3078 1710 3081
rect 1786 3078 1806 3081
rect 1834 3078 1846 3081
rect 1958 3081 1961 3088
rect 3830 3082 3833 3088
rect 1958 3078 1966 3081
rect 2074 3078 2102 3081
rect 2354 3078 2473 3081
rect 86 3068 206 3071
rect 290 3068 310 3071
rect 426 3068 486 3071
rect 522 3068 654 3071
rect 658 3068 774 3071
rect 826 3068 870 3071
rect 874 3068 934 3071
rect 938 3068 942 3071
rect 1042 3068 1214 3071
rect 1346 3068 1358 3071
rect 1378 3068 1390 3071
rect 1394 3068 1446 3071
rect 1450 3068 1454 3071
rect 1514 3068 1614 3071
rect 1626 3068 1662 3071
rect 1698 3068 1870 3071
rect 1882 3068 1910 3071
rect 1942 3068 1950 3071
rect 2138 3068 2158 3071
rect 2162 3068 2270 3071
rect 2310 3071 2313 3078
rect 2470 3072 2473 3078
rect 2570 3078 2614 3081
rect 2714 3078 2806 3081
rect 2826 3078 2894 3081
rect 2898 3078 2902 3081
rect 3042 3078 3046 3081
rect 3066 3078 3350 3081
rect 3466 3078 3489 3081
rect 3498 3078 3617 3081
rect 3626 3078 3686 3081
rect 3730 3078 3750 3081
rect 3922 3078 3926 3081
rect 4034 3078 4038 3081
rect 4226 3078 4558 3081
rect 4562 3078 4582 3081
rect 4778 3078 4798 3081
rect 4858 3078 4878 3081
rect 5074 3078 5086 3081
rect 2310 3068 2318 3071
rect 2338 3068 2422 3071
rect 2518 3071 2521 3078
rect 2506 3068 2521 3071
rect 2526 3072 2529 3078
rect 2554 3068 2558 3071
rect 2578 3068 2582 3071
rect 2770 3068 2822 3071
rect 2858 3068 2862 3071
rect 2906 3068 3030 3071
rect 3218 3068 3318 3071
rect 3330 3068 3334 3071
rect 3346 3068 3470 3071
rect 3486 3071 3489 3078
rect 3614 3072 3617 3078
rect 3486 3068 3502 3071
rect 3594 3068 3614 3071
rect 3718 3071 3721 3078
rect 3718 3068 3774 3071
rect 3814 3071 3817 3078
rect 3814 3068 3862 3071
rect 3938 3068 3942 3071
rect 4018 3068 4054 3071
rect 4086 3068 4198 3071
rect 4230 3068 4318 3071
rect 4354 3068 4374 3071
rect 4378 3068 4406 3071
rect 4434 3068 4550 3071
rect 4658 3068 4694 3071
rect 5010 3068 5126 3071
rect 86 3062 89 3068
rect 122 3058 174 3061
rect 178 3058 182 3061
rect 238 3061 241 3068
rect 342 3062 345 3068
rect 238 3058 294 3061
rect 402 3058 414 3061
rect 418 3058 574 3061
rect 578 3058 622 3061
rect 990 3058 1158 3061
rect 1202 3058 1206 3061
rect 1222 3061 1225 3068
rect 1942 3062 1945 3068
rect 2422 3062 2425 3068
rect 1222 3058 1286 3061
rect 1298 3058 1310 3061
rect 1378 3058 1454 3061
rect 1474 3058 1670 3061
rect 1694 3058 1905 3061
rect 1914 3058 1918 3061
rect 1986 3058 2001 3061
rect 2042 3058 2078 3061
rect 2186 3058 2262 3061
rect 2490 3058 2494 3061
rect 2698 3058 2774 3061
rect 2890 3058 2913 3061
rect 2922 3058 3014 3061
rect 3018 3058 3022 3061
rect 3086 3058 3094 3061
rect 3142 3061 3145 3068
rect 3526 3062 3529 3068
rect 3098 3058 3145 3061
rect 3314 3058 3342 3061
rect 3402 3058 3454 3061
rect 3458 3058 3510 3061
rect 3514 3058 3518 3061
rect 3566 3061 3569 3068
rect 3566 3058 3686 3061
rect 3798 3061 3801 3068
rect 3918 3062 3921 3068
rect 3798 3058 3854 3061
rect 3954 3058 3958 3061
rect 3990 3061 3993 3068
rect 4086 3062 4089 3068
rect 3990 3058 3998 3061
rect 4018 3058 4030 3061
rect 4230 3061 4233 3068
rect 4230 3058 4238 3061
rect 4250 3058 4262 3061
rect 4334 3061 4337 3068
rect 4314 3058 4337 3061
rect 4342 3062 4345 3068
rect 4354 3058 4454 3061
rect 4490 3058 4494 3061
rect 4522 3058 4638 3061
rect 4674 3058 4702 3061
rect 4706 3058 4870 3061
rect 5138 3058 5158 3061
rect 378 3048 406 3051
rect 690 3048 694 3051
rect 838 3051 841 3058
rect 826 3048 841 3051
rect 990 3052 993 3058
rect 1350 3052 1353 3058
rect 1098 3048 1182 3051
rect 1186 3048 1206 3051
rect 1362 3048 1478 3051
rect 1490 3048 1582 3051
rect 1594 3048 1646 3051
rect 1694 3051 1697 3058
rect 1650 3048 1697 3051
rect 1706 3048 1718 3051
rect 1738 3048 1766 3051
rect 1786 3048 1838 3051
rect 1902 3051 1905 3058
rect 1926 3051 1929 3058
rect 1902 3048 1929 3051
rect 1998 3052 2001 3058
rect 2286 3052 2289 3058
rect 2018 3048 2134 3051
rect 2234 3048 2273 3051
rect 2502 3051 2505 3058
rect 2314 3048 2505 3051
rect 2510 3052 2513 3058
rect 2542 3051 2545 3058
rect 2542 3048 2574 3051
rect 2602 3048 2710 3051
rect 2730 3048 2878 3051
rect 2910 3051 2913 3058
rect 2886 3048 2905 3051
rect 2910 3048 2950 3051
rect 3114 3048 3142 3051
rect 3146 3048 3246 3051
rect 3474 3048 3486 3051
rect 3490 3048 3518 3051
rect 3530 3048 3542 3051
rect 3546 3048 3574 3051
rect 3650 3048 3686 3051
rect 3946 3048 4110 3051
rect 4114 3048 4134 3051
rect 4146 3048 4241 3051
rect 66 3038 206 3041
rect 210 3038 326 3041
rect 330 3038 606 3041
rect 834 3038 870 3041
rect 938 3038 942 3041
rect 954 3038 1070 3041
rect 1074 3038 1102 3041
rect 1106 3038 1270 3041
rect 1274 3038 1286 3041
rect 1734 3041 1737 3048
rect 2270 3042 2273 3048
rect 2886 3042 2889 3048
rect 2902 3042 2905 3048
rect 4238 3042 4241 3048
rect 4290 3048 4302 3051
rect 4306 3048 4449 3051
rect 4474 3048 4494 3051
rect 4570 3048 4590 3051
rect 4594 3048 4606 3051
rect 4618 3048 4630 3051
rect 4634 3048 4862 3051
rect 4974 3051 4977 3058
rect 4962 3048 4977 3051
rect 5050 3048 5062 3051
rect 5066 3048 5070 3051
rect 5074 3048 5086 3051
rect 5090 3048 5118 3051
rect 5154 3048 5158 3051
rect 1290 3038 1737 3041
rect 1762 3038 1766 3041
rect 1946 3038 2046 3041
rect 2058 3038 2230 3041
rect 2418 3038 2430 3041
rect 2442 3038 2502 3041
rect 2722 3038 2870 3041
rect 3106 3038 3342 3041
rect 3418 3038 3505 3041
rect 3522 3038 3534 3041
rect 3538 3038 3630 3041
rect 3914 3038 3950 3041
rect 4010 3038 4070 3041
rect 4278 3041 4281 3048
rect 4446 3042 4449 3048
rect 4278 3038 4318 3041
rect 4346 3038 4374 3041
rect 4546 3038 4622 3041
rect 4626 3038 4726 3041
rect 4730 3038 4737 3041
rect 4862 3038 4926 3041
rect 5074 3038 5086 3041
rect 5090 3038 5174 3041
rect 250 3028 358 3031
rect 362 3028 430 3031
rect 622 3031 625 3038
rect 3502 3032 3505 3038
rect 622 3028 894 3031
rect 962 3028 1094 3031
rect 1146 3028 1230 3031
rect 1258 3028 1358 3031
rect 1402 3028 1622 3031
rect 1626 3028 1662 3031
rect 1794 3028 1822 3031
rect 1874 3028 2006 3031
rect 2130 3028 2270 3031
rect 2282 3028 2438 3031
rect 2442 3028 2526 3031
rect 2554 3028 2822 3031
rect 2826 3028 2838 3031
rect 2842 3028 2846 3031
rect 3514 3028 3886 3031
rect 3898 3028 4270 3031
rect 4374 3031 4377 3038
rect 4862 3032 4865 3038
rect 4374 3028 4518 3031
rect 4598 3028 4614 3031
rect 4686 3028 4774 3031
rect 394 3018 614 3021
rect 934 3021 937 3028
rect 934 3018 998 3021
rect 1190 3018 1198 3021
rect 1202 3018 1486 3021
rect 1494 3018 1502 3021
rect 1506 3018 1606 3021
rect 1710 3021 1713 3028
rect 4278 3022 4281 3028
rect 4598 3022 4601 3028
rect 4686 3022 4689 3028
rect 1710 3018 1854 3021
rect 2066 3018 2342 3021
rect 2346 3018 2910 3021
rect 2914 3018 3430 3021
rect 3434 3018 4022 3021
rect 4026 3018 4094 3021
rect 4170 3018 4238 3021
rect 4482 3018 4574 3021
rect 4610 3018 4622 3021
rect 4626 3018 4654 3021
rect 978 3008 998 3011
rect 1002 3008 1038 3011
rect 1586 3008 1702 3011
rect 1818 3008 1934 3011
rect 1978 3008 1990 3011
rect 2146 3008 2270 3011
rect 2338 3008 2398 3011
rect 2466 3008 2534 3011
rect 2618 3008 2934 3011
rect 3634 3008 3774 3011
rect 3842 3008 3934 3011
rect 3970 3008 4054 3011
rect 4386 3008 4462 3011
rect 4466 3008 4478 3011
rect 4490 3008 4622 3011
rect 4706 3008 4982 3011
rect 536 3003 538 3007
rect 542 3003 545 3007
rect 550 3003 552 3007
rect 1238 3002 1241 3008
rect 1560 3003 1562 3007
rect 1566 3003 1569 3007
rect 1574 3003 1576 3007
rect 2584 3003 2586 3007
rect 2590 3003 2593 3007
rect 2598 3003 2600 3007
rect 3406 3002 3409 3008
rect 3608 3003 3610 3007
rect 3614 3003 3617 3007
rect 3622 3003 3624 3007
rect 4632 3003 4634 3007
rect 4638 3003 4641 3007
rect 4646 3003 4648 3007
rect 1042 2998 1142 3001
rect 1466 2998 1502 3001
rect 1602 2998 1774 3001
rect 1786 2998 2406 3001
rect 2426 2998 2574 3001
rect 2754 2998 2958 3001
rect 3138 2998 3270 3001
rect 3410 2998 3558 3001
rect 3562 2998 3566 3001
rect 3762 2998 3766 3001
rect 4010 2998 4326 3001
rect 4458 2998 4534 3001
rect 4658 2998 4814 3001
rect 4818 2998 4870 3001
rect 346 2988 358 2991
rect 370 2988 558 2991
rect 562 2988 918 2991
rect 922 2988 974 2991
rect 1370 2988 1422 2991
rect 1538 2988 1758 2991
rect 1826 2988 1870 2991
rect 1922 2988 1982 2991
rect 2026 2988 2182 2991
rect 2282 2988 2838 2991
rect 2954 2988 3022 2991
rect 3026 2988 3630 2991
rect 3634 2988 3710 2991
rect 3718 2988 3974 2991
rect 4002 2988 4025 2991
rect 4210 2988 4462 2991
rect 4466 2988 4654 2991
rect 4718 2988 4766 2991
rect 4794 2988 4798 2991
rect 4802 2988 4990 2991
rect 18 2978 102 2981
rect 154 2978 430 2981
rect 754 2978 806 2981
rect 922 2978 974 2981
rect 1018 2978 1134 2981
rect 1162 2978 1398 2981
rect 1442 2978 1534 2981
rect 1554 2978 1766 2981
rect 1798 2981 1801 2988
rect 2222 2982 2225 2988
rect 3718 2982 3721 2988
rect 4022 2982 4025 2988
rect 1798 2978 1878 2981
rect 2018 2978 2038 2981
rect 2042 2978 2166 2981
rect 2266 2978 2422 2981
rect 2426 2978 2494 2981
rect 2498 2978 3046 2981
rect 3194 2978 3214 2981
rect 3218 2978 3238 2981
rect 3246 2978 3494 2981
rect 3498 2978 3518 2981
rect 3522 2978 3582 2981
rect 3762 2978 3854 2981
rect 4090 2978 4294 2981
rect 4298 2978 4342 2981
rect 4718 2981 4721 2988
rect 4530 2978 4721 2981
rect 4730 2978 5070 2981
rect 346 2968 393 2971
rect 410 2968 486 2971
rect 566 2971 569 2978
rect 3246 2972 3249 2978
rect 566 2968 910 2971
rect 1018 2968 1318 2971
rect 1362 2968 1390 2971
rect 1594 2968 1662 2971
rect 1778 2968 2006 2971
rect 2138 2968 2246 2971
rect 2538 2968 2542 2971
rect 2578 2968 2630 2971
rect 2682 2968 2686 2971
rect 2706 2968 2710 2971
rect 2778 2968 2782 2971
rect 3026 2968 3246 2971
rect 3346 2968 3534 2971
rect 3538 2968 3550 2971
rect 3682 2968 3886 2971
rect 4194 2968 4550 2971
rect 4554 2968 4718 2971
rect 4778 2968 4782 2971
rect 4786 2968 4870 2971
rect 4946 2968 4950 2971
rect 4986 2968 5158 2971
rect 5162 2968 5174 2971
rect 390 2962 393 2968
rect 282 2958 374 2961
rect 494 2961 497 2968
rect 518 2961 521 2968
rect 494 2958 521 2961
rect 562 2958 574 2961
rect 650 2958 662 2961
rect 674 2958 686 2961
rect 774 2958 782 2961
rect 786 2958 1022 2961
rect 1122 2958 1174 2961
rect 1354 2958 1366 2961
rect 1678 2958 1686 2961
rect 1826 2958 1838 2961
rect 1850 2958 1942 2961
rect 2030 2958 2102 2961
rect 2470 2961 2473 2968
rect 2386 2958 2473 2961
rect 2486 2962 2489 2968
rect 3286 2962 3289 2968
rect 2498 2958 2734 2961
rect 2762 2958 2774 2961
rect 2778 2958 2790 2961
rect 2794 2958 2814 2961
rect 2922 2958 2982 2961
rect 2986 2958 3054 2961
rect 3074 2958 3134 2961
rect 3334 2958 3390 2961
rect 3722 2958 3726 2961
rect 3778 2958 3782 2961
rect 3814 2958 3822 2961
rect 3826 2958 3833 2961
rect 3842 2958 3934 2961
rect 3962 2958 3982 2961
rect 4106 2958 4182 2961
rect 4530 2958 4582 2961
rect 4594 2958 4606 2961
rect 4690 2958 4694 2961
rect 4722 2958 5030 2961
rect -26 2951 -22 2952
rect -26 2948 14 2951
rect 70 2951 73 2958
rect 70 2948 126 2951
rect 186 2948 198 2951
rect 202 2948 206 2951
rect 470 2951 473 2958
rect 1806 2952 1809 2958
rect 2030 2952 2033 2958
rect 362 2948 473 2951
rect 490 2948 510 2951
rect 658 2948 678 2951
rect 778 2948 782 2951
rect 826 2948 838 2951
rect 874 2948 878 2951
rect 954 2948 966 2951
rect 1042 2948 1046 2951
rect 1122 2948 1142 2951
rect 1146 2948 1150 2951
rect 1162 2948 1190 2951
rect 1338 2948 1342 2951
rect 1378 2948 1478 2951
rect 1546 2948 1609 2951
rect 1626 2948 1630 2951
rect 1642 2948 1694 2951
rect 1706 2948 1734 2951
rect 1826 2948 2014 2951
rect 2074 2948 2166 2951
rect 2170 2948 2294 2951
rect 2410 2948 2486 2951
rect 2498 2948 2518 2951
rect 2562 2948 2606 2951
rect 2626 2948 2630 2951
rect 2650 2948 2742 2951
rect 2798 2948 2806 2951
rect 2894 2951 2897 2958
rect 2810 2948 2897 2951
rect 2954 2948 2998 2951
rect 3122 2948 3126 2951
rect 3130 2948 3150 2951
rect 3334 2951 3337 2958
rect 3202 2948 3337 2951
rect 3462 2951 3465 2958
rect 3362 2948 3433 2951
rect 3462 2948 3494 2951
rect 3542 2951 3545 2958
rect 3606 2951 3609 2958
rect 3542 2948 3590 2951
rect 566 2942 569 2948
rect 678 2942 681 2948
rect 734 2942 737 2948
rect 154 2938 222 2941
rect 226 2938 230 2941
rect 362 2938 366 2941
rect 426 2938 526 2941
rect 754 2938 790 2941
rect 794 2938 798 2941
rect 810 2938 926 2941
rect 1114 2938 1118 2941
rect 1142 2938 1150 2941
rect 1154 2938 1246 2941
rect 1270 2941 1273 2948
rect 1270 2938 1302 2941
rect 1314 2938 1318 2941
rect 1346 2938 1406 2941
rect 1418 2938 1438 2941
rect 1606 2941 1609 2948
rect 1606 2938 1694 2941
rect 1706 2938 1710 2941
rect 1730 2938 1750 2941
rect 1754 2938 1782 2941
rect 1786 2938 1998 2941
rect 2018 2938 2158 2941
rect 2170 2938 2174 2941
rect 2210 2938 2238 2941
rect 2298 2938 2310 2941
rect 2322 2938 2326 2941
rect 2342 2938 2446 2941
rect 2534 2941 2537 2948
rect 3430 2942 3433 2948
rect 3606 2948 3662 2951
rect 3690 2948 3710 2951
rect 3722 2948 3726 2951
rect 3794 2948 3822 2951
rect 3830 2951 3833 2958
rect 4310 2952 4313 2958
rect 3830 2948 3878 2951
rect 3962 2948 3966 2951
rect 4042 2948 4062 2951
rect 4066 2948 4142 2951
rect 4326 2948 4334 2951
rect 4338 2948 4398 2951
rect 4418 2948 4478 2951
rect 4634 2948 4822 2951
rect 4850 2948 4894 2951
rect 4898 2948 4998 2951
rect 5058 2948 5094 2951
rect 5166 2948 5174 2951
rect 2534 2938 2590 2941
rect 2594 2938 2622 2941
rect 2706 2938 2830 2941
rect 2978 2938 2982 2941
rect 3002 2938 3102 2941
rect 3114 2938 3182 2941
rect 3266 2938 3278 2941
rect 3322 2938 3326 2941
rect 3538 2938 3686 2941
rect 3706 2938 4030 2941
rect 4042 2938 4118 2941
rect 4122 2938 4134 2941
rect 4178 2938 4182 2941
rect 4310 2941 4313 2948
rect 4310 2938 4326 2941
rect 4402 2938 4406 2941
rect 4558 2941 4561 2948
rect 4838 2942 4841 2948
rect 5166 2942 5169 2948
rect 4458 2938 4561 2941
rect 4682 2938 4694 2941
rect 4970 2938 5118 2941
rect 5130 2938 5150 2941
rect 526 2932 529 2938
rect 654 2932 657 2938
rect 2286 2932 2289 2938
rect 2342 2932 2345 2938
rect 4206 2932 4209 2938
rect 4342 2932 4345 2938
rect 18 2928 238 2931
rect 458 2928 462 2931
rect 682 2928 782 2931
rect 962 2928 982 2931
rect 1018 2928 1070 2931
rect 1074 2928 1150 2931
rect 1186 2928 1190 2931
rect 1306 2928 1430 2931
rect 1818 2928 1822 2931
rect 1834 2928 1910 2931
rect 2002 2928 2014 2931
rect 2154 2928 2286 2931
rect 2490 2928 2542 2931
rect 2610 2928 2614 2931
rect 2698 2928 2726 2931
rect 2762 2928 3198 2931
rect 3202 2928 3238 2931
rect 3522 2928 3574 2931
rect 3618 2928 3798 2931
rect 3802 2928 3854 2931
rect 3874 2928 4030 2931
rect 4082 2928 4086 2931
rect 4130 2928 4166 2931
rect 4446 2931 4449 2938
rect 4402 2928 4606 2931
rect 4874 2928 4902 2931
rect 5106 2928 5166 2931
rect 58 2918 118 2921
rect 122 2918 142 2921
rect 146 2918 318 2921
rect 322 2918 414 2921
rect 634 2918 774 2921
rect 862 2921 865 2928
rect 778 2918 865 2921
rect 1010 2918 1014 2921
rect 1074 2918 1222 2921
rect 1298 2918 1350 2921
rect 1354 2918 1414 2921
rect 1830 2921 1833 2928
rect 1682 2918 1833 2921
rect 2050 2918 2254 2921
rect 2282 2918 2502 2921
rect 2626 2918 2662 2921
rect 2762 2918 2766 2921
rect 2770 2918 2814 2921
rect 2858 2918 2950 2921
rect 2954 2918 3022 2921
rect 3154 2918 3174 2921
rect 3178 2918 3193 2921
rect 3230 2918 3238 2921
rect 3242 2918 3318 2921
rect 3330 2918 3534 2921
rect 3538 2918 3766 2921
rect 3770 2918 3830 2921
rect 4118 2921 4121 2928
rect 3954 2918 4121 2921
rect 4262 2922 4265 2928
rect 4578 2918 4582 2921
rect 4586 2918 4598 2921
rect 4690 2918 4966 2921
rect 1462 2912 1465 2918
rect 218 2908 238 2911
rect 250 2908 582 2911
rect 586 2908 774 2911
rect 954 2908 958 2911
rect 1082 2908 1446 2911
rect 1546 2908 1598 2911
rect 1910 2911 1913 2918
rect 1634 2908 1913 2911
rect 2266 2908 2318 2911
rect 2522 2908 2622 2911
rect 2634 2908 2678 2911
rect 2786 2908 2902 2911
rect 3074 2908 3078 2911
rect 3190 2911 3193 2918
rect 4462 2912 4465 2918
rect 3190 2908 3750 2911
rect 3970 2908 4006 2911
rect 4026 2908 4054 2911
rect 4138 2908 4214 2911
rect 4250 2908 4334 2911
rect 4562 2908 4662 2911
rect 4818 2908 5142 2911
rect 1048 2903 1050 2907
rect 1054 2903 1057 2907
rect 1062 2903 1064 2907
rect 2022 2902 2025 2908
rect 2072 2903 2074 2907
rect 2078 2903 2081 2907
rect 2086 2903 2088 2907
rect 3096 2903 3098 2907
rect 3102 2903 3105 2907
rect 3110 2903 3112 2907
rect 4112 2903 4114 2907
rect 4118 2903 4121 2907
rect 4126 2903 4128 2907
rect 74 2898 190 2901
rect 242 2898 246 2901
rect 346 2898 574 2901
rect 642 2898 662 2901
rect 866 2898 958 2901
rect 1098 2898 1374 2901
rect 1378 2898 1782 2901
rect 1930 2898 1958 2901
rect 2162 2898 2462 2901
rect 2466 2898 2486 2901
rect 2602 2898 2662 2901
rect 2770 2898 2774 2901
rect 2778 2898 2870 2901
rect 2890 2898 3030 2901
rect 3122 2898 3166 2901
rect 3170 2898 3750 2901
rect 3850 2898 4078 2901
rect 4146 2898 4182 2901
rect 4226 2898 4678 2901
rect 4698 2898 4846 2901
rect 4906 2898 4950 2901
rect 5026 2898 5030 2901
rect 18 2888 134 2891
rect 138 2888 158 2891
rect 186 2888 326 2891
rect 650 2888 670 2891
rect 706 2888 822 2891
rect 842 2888 942 2891
rect 954 2888 1001 2891
rect 998 2882 1001 2888
rect 1082 2888 1086 2891
rect 1098 2888 1222 2891
rect 1234 2888 1302 2891
rect 1306 2888 1318 2891
rect 1346 2888 1358 2891
rect 1474 2888 1542 2891
rect 1554 2888 1582 2891
rect 1666 2888 1670 2891
rect 1698 2888 1742 2891
rect 1746 2888 1782 2891
rect 1834 2888 1838 2891
rect 1938 2888 1958 2891
rect 1970 2888 2006 2891
rect 2042 2888 2070 2891
rect 2098 2888 2150 2891
rect 2306 2888 2310 2891
rect 2642 2888 2646 2891
rect 2810 2888 2942 2891
rect 3066 2888 3166 2891
rect 3194 2888 3206 2891
rect 3242 2888 3358 2891
rect 3402 2888 3462 2891
rect 3470 2888 3478 2891
rect 3482 2888 3494 2891
rect 3610 2888 3630 2891
rect 3674 2888 3678 2891
rect 3890 2888 4038 2891
rect 4154 2888 4254 2891
rect 4290 2888 4294 2891
rect 4314 2888 4366 2891
rect 4594 2888 4702 2891
rect 4802 2888 5041 2891
rect 5066 2888 5182 2891
rect 1030 2882 1033 2888
rect 90 2878 158 2881
rect 906 2878 910 2881
rect 1058 2878 1094 2881
rect 1098 2878 1105 2881
rect 1450 2878 1486 2881
rect 1538 2878 1582 2881
rect 1626 2878 1630 2881
rect 1666 2878 3278 2881
rect 3322 2878 3342 2881
rect 3398 2881 3401 2888
rect 3362 2878 3401 2881
rect 3450 2878 3654 2881
rect 3682 2878 3958 2881
rect 3962 2878 4158 2881
rect 4170 2878 4190 2881
rect 4458 2878 4614 2881
rect 4626 2878 4670 2881
rect 4750 2881 4753 2888
rect 5038 2882 5041 2888
rect 4674 2878 4753 2881
rect 4890 2878 4918 2881
rect 5046 2878 5054 2881
rect 5058 2878 5086 2881
rect 934 2872 937 2878
rect 282 2868 366 2871
rect 402 2868 526 2871
rect 530 2868 598 2871
rect 762 2868 766 2871
rect 898 2868 902 2871
rect 986 2868 1086 2871
rect 1090 2868 1110 2871
rect 1190 2868 1214 2871
rect 1234 2868 1318 2871
rect 1330 2868 1446 2871
rect 1450 2868 1494 2871
rect 1506 2868 1510 2871
rect 1522 2868 1542 2871
rect 1586 2868 1630 2871
rect 1650 2868 1678 2871
rect 1754 2868 1790 2871
rect 1858 2868 1862 2871
rect 1898 2868 1902 2871
rect 1946 2868 2038 2871
rect 2130 2868 2214 2871
rect 2226 2868 2318 2871
rect 2322 2868 2414 2871
rect 2426 2868 2446 2871
rect 2474 2868 2510 2871
rect 2554 2868 2558 2871
rect 2650 2868 2654 2871
rect 2666 2868 2670 2871
rect 2690 2868 2782 2871
rect 2794 2868 2814 2871
rect 2850 2868 2854 2871
rect 2970 2868 2990 2871
rect 3058 2868 3142 2871
rect 3146 2868 3326 2871
rect 3334 2868 3350 2871
rect 3482 2868 3510 2871
rect 3514 2868 3558 2871
rect 3698 2868 3830 2871
rect 3874 2868 3910 2871
rect 4230 2871 4233 2878
rect 3962 2868 4233 2871
rect 4290 2868 4433 2871
rect 4442 2868 4470 2871
rect 4530 2868 4598 2871
rect 4642 2868 4662 2871
rect 4890 2868 4910 2871
rect 5022 2871 5025 2878
rect 4914 2868 5054 2871
rect 5058 2868 5118 2871
rect 102 2861 105 2868
rect 102 2858 398 2861
rect 466 2858 494 2861
rect 546 2858 574 2861
rect 702 2861 705 2868
rect 1182 2862 1185 2868
rect 1190 2862 1193 2868
rect 594 2858 705 2861
rect 786 2858 814 2861
rect 874 2858 1094 2861
rect 1106 2858 1110 2861
rect 1130 2858 1166 2861
rect 1274 2858 1582 2861
rect 1638 2861 1641 2868
rect 2838 2862 2841 2868
rect 1586 2858 1641 2861
rect 1674 2858 1774 2861
rect 1778 2858 2102 2861
rect 2106 2858 2134 2861
rect 2138 2858 2798 2861
rect 2886 2861 2889 2868
rect 3334 2862 3337 2868
rect 2886 2858 2918 2861
rect 2978 2858 2982 2861
rect 3042 2858 3110 2861
rect 3178 2858 3206 2861
rect 3346 2858 3390 2861
rect 3422 2861 3425 2868
rect 4006 2862 4009 2868
rect 3402 2858 3425 2861
rect 3506 2858 3510 2861
rect 3618 2858 3697 2861
rect 3754 2858 3766 2861
rect 3770 2858 3806 2861
rect 3810 2858 3846 2861
rect 3850 2858 3886 2861
rect 4058 2858 4102 2861
rect 4146 2858 4150 2861
rect 4170 2858 4206 2861
rect 4262 2861 4265 2868
rect 4430 2862 4433 2868
rect 4518 2862 4521 2868
rect 4734 2862 4737 2868
rect 4262 2858 4350 2861
rect 4450 2858 4454 2861
rect 4546 2858 4550 2861
rect 4618 2858 4622 2861
rect 4674 2858 4710 2861
rect 4714 2858 4726 2861
rect 4750 2861 4753 2868
rect 4814 2861 4817 2868
rect 4750 2858 4817 2861
rect 5070 2858 5142 2861
rect 3550 2852 3553 2858
rect 3694 2852 3697 2858
rect 226 2848 254 2851
rect 258 2848 430 2851
rect 498 2848 558 2851
rect 562 2848 710 2851
rect 762 2848 870 2851
rect 926 2848 934 2851
rect 938 2848 982 2851
rect 1274 2848 1342 2851
rect 1346 2848 1382 2851
rect 1394 2848 1470 2851
rect 1486 2848 1494 2851
rect 1498 2848 1510 2851
rect 1538 2848 1558 2851
rect 1594 2848 1598 2851
rect 1610 2848 1686 2851
rect 1738 2848 1750 2851
rect 1762 2848 1846 2851
rect 1882 2848 1902 2851
rect 2002 2848 2014 2851
rect 2050 2848 2054 2851
rect 2146 2848 2166 2851
rect 2306 2848 2310 2851
rect 2386 2848 2430 2851
rect 2466 2848 2470 2851
rect 2482 2848 2849 2851
rect 3018 2848 3022 2851
rect 3082 2848 3094 2851
rect 3122 2848 3206 2851
rect 3210 2848 3217 2851
rect 3258 2848 3446 2851
rect 3578 2848 3678 2851
rect 3718 2848 3758 2851
rect 3782 2848 3846 2851
rect 3874 2848 3910 2851
rect 3918 2851 3921 2858
rect 3918 2848 3942 2851
rect 4026 2848 4094 2851
rect 4254 2851 4257 2858
rect 4170 2848 4257 2851
rect 4458 2848 4462 2851
rect 4530 2848 4630 2851
rect 4634 2848 4710 2851
rect 4714 2848 4790 2851
rect 4822 2851 4825 2858
rect 5070 2852 5073 2858
rect 4822 2848 4958 2851
rect 5222 2851 5226 2852
rect 5182 2848 5226 2851
rect 146 2838 350 2841
rect 354 2838 374 2841
rect 378 2838 694 2841
rect 874 2838 934 2841
rect 1082 2838 1110 2841
rect 1142 2841 1145 2848
rect 1142 2838 1270 2841
rect 1282 2838 1334 2841
rect 1338 2838 1342 2841
rect 1354 2838 1502 2841
rect 1506 2838 1678 2841
rect 1710 2841 1713 2848
rect 1910 2841 1913 2848
rect 1710 2838 1753 2841
rect 1910 2838 2174 2841
rect 2178 2838 2382 2841
rect 2506 2838 2518 2841
rect 2522 2838 2606 2841
rect 2754 2838 2798 2841
rect 2834 2838 2838 2841
rect 2846 2841 2849 2848
rect 3718 2842 3721 2848
rect 3782 2842 3785 2848
rect 2846 2838 3278 2841
rect 3282 2838 3334 2841
rect 3346 2838 3366 2841
rect 3418 2838 3478 2841
rect 3514 2838 3566 2841
rect 3810 2838 3822 2841
rect 3826 2838 3894 2841
rect 4042 2838 4217 2841
rect 4626 2838 4790 2841
rect 5182 2841 5185 2848
rect 4794 2838 5185 2841
rect 1750 2832 1753 2838
rect 698 2828 718 2831
rect 722 2828 1230 2831
rect 1306 2828 1334 2831
rect 1362 2828 1518 2831
rect 1554 2828 1678 2831
rect 1690 2828 1718 2831
rect 1874 2828 1878 2831
rect 2122 2828 2678 2831
rect 2682 2828 2750 2831
rect 2818 2828 2878 2831
rect 2882 2828 2886 2831
rect 3170 2828 3246 2831
rect 3258 2828 3302 2831
rect 3314 2828 3390 2831
rect 3934 2831 3937 2838
rect 3402 2828 3937 2831
rect 4214 2832 4217 2838
rect 4338 2828 4422 2831
rect 4426 2828 4510 2831
rect 4570 2828 4654 2831
rect 4842 2828 4974 2831
rect 778 2818 2150 2821
rect 2154 2818 2206 2821
rect 2474 2818 3086 2821
rect 3330 2818 3574 2821
rect 3650 2818 3654 2821
rect 3658 2818 3998 2821
rect 4202 2818 4222 2821
rect 4354 2818 4606 2821
rect 4614 2818 4846 2821
rect 5018 2818 5158 2821
rect 762 2808 1441 2811
rect 1458 2808 1550 2811
rect 1682 2808 1990 2811
rect 2050 2808 2286 2811
rect 2338 2808 2414 2811
rect 2514 2808 2526 2811
rect 2794 2808 2894 2811
rect 3354 2808 3358 2811
rect 3366 2808 3526 2811
rect 3682 2808 3902 2811
rect 4090 2808 4182 2811
rect 4202 2808 4382 2811
rect 4614 2811 4617 2818
rect 4498 2808 4617 2811
rect 4674 2808 4910 2811
rect 536 2803 538 2807
rect 542 2803 545 2807
rect 550 2803 552 2807
rect 1438 2802 1441 2808
rect 1560 2803 1562 2807
rect 1566 2803 1569 2807
rect 1574 2803 1576 2807
rect 2584 2803 2586 2807
rect 2590 2803 2593 2807
rect 2598 2803 2600 2807
rect 610 2798 646 2801
rect 794 2798 838 2801
rect 842 2798 1190 2801
rect 1202 2798 1390 2801
rect 1482 2798 1502 2801
rect 1618 2798 1726 2801
rect 1786 2798 1966 2801
rect 2034 2798 2046 2801
rect 2058 2798 2102 2801
rect 3366 2801 3369 2808
rect 3608 2803 3610 2807
rect 3614 2803 3617 2807
rect 3622 2803 3624 2807
rect 4632 2803 4634 2807
rect 4638 2803 4641 2807
rect 4646 2803 4648 2807
rect 2626 2798 3369 2801
rect 3394 2798 3462 2801
rect 3770 2798 3910 2801
rect 3938 2798 3974 2801
rect 4090 2798 4166 2801
rect 4210 2798 4230 2801
rect 4250 2798 4534 2801
rect 4746 2798 4758 2801
rect 4930 2798 4966 2801
rect 410 2788 414 2791
rect 418 2788 974 2791
rect 1050 2788 1118 2791
rect 1138 2788 1166 2791
rect 1170 2788 1702 2791
rect 1738 2788 1798 2791
rect 1810 2788 1886 2791
rect 1890 2788 2406 2791
rect 2410 2788 2526 2791
rect 2818 2788 2822 2791
rect 2834 2788 2838 2791
rect 3034 2788 3174 2791
rect 3250 2788 3286 2791
rect 3314 2788 3342 2791
rect 3346 2788 3494 2791
rect 3506 2788 4945 2791
rect 4942 2782 4945 2788
rect 666 2778 870 2781
rect 962 2778 1782 2781
rect 1794 2778 1950 2781
rect 2138 2778 2190 2781
rect 2242 2778 2302 2781
rect 2306 2778 2350 2781
rect 2522 2778 2630 2781
rect 2858 2778 2902 2781
rect 3106 2778 3142 2781
rect 3146 2778 3166 2781
rect 3282 2778 4478 2781
rect 4570 2778 4646 2781
rect 4906 2778 4926 2781
rect 250 2768 262 2771
rect 266 2768 366 2771
rect 506 2768 582 2771
rect 746 2768 1126 2771
rect 1130 2768 1294 2771
rect 1298 2768 1494 2771
rect 1498 2768 1742 2771
rect 2034 2768 2134 2771
rect 2234 2768 2446 2771
rect 2458 2768 2606 2771
rect 2770 2768 2798 2771
rect 3050 2768 3086 2771
rect 3226 2768 3262 2771
rect 3378 2768 3478 2771
rect 3554 2768 3558 2771
rect 3574 2768 3582 2771
rect 3586 2768 3614 2771
rect 3622 2768 3638 2771
rect 3662 2768 3726 2771
rect 3730 2768 3830 2771
rect 3890 2768 3894 2771
rect 3914 2768 4350 2771
rect 4354 2768 4462 2771
rect 4498 2768 4758 2771
rect 4762 2768 5182 2771
rect 5222 2771 5226 2772
rect 5194 2768 5226 2771
rect 498 2758 550 2761
rect 810 2758 854 2761
rect 994 2758 1198 2761
rect 1262 2758 1270 2761
rect 1274 2758 1350 2761
rect 1426 2758 1470 2761
rect 1486 2758 1494 2761
rect 1498 2758 1590 2761
rect 1666 2758 1678 2761
rect 1790 2761 1793 2768
rect 1754 2758 1793 2761
rect 1854 2762 1857 2768
rect 1990 2762 1993 2768
rect 1874 2758 1990 2761
rect 2090 2758 2094 2761
rect 2130 2758 2158 2761
rect 2210 2758 2222 2761
rect 2434 2758 2486 2761
rect 2538 2758 2622 2761
rect 2714 2758 2782 2761
rect 2798 2761 2801 2768
rect 2830 2761 2833 2768
rect 2798 2758 2833 2761
rect 2842 2758 2846 2761
rect 2894 2761 2897 2768
rect 2890 2758 2897 2761
rect 3550 2761 3553 2768
rect 3042 2758 3553 2761
rect 3622 2762 3625 2768
rect 3662 2762 3665 2768
rect 3854 2762 3857 2768
rect 3878 2762 3881 2768
rect 3882 2758 3998 2761
rect 4178 2758 4182 2761
rect 4186 2758 4270 2761
rect 4282 2758 4574 2761
rect 4666 2758 4798 2761
rect 4898 2758 4902 2761
rect 5018 2758 5022 2761
rect 5034 2758 5110 2761
rect 382 2752 385 2758
rect 654 2752 657 2758
rect 1862 2752 1865 2758
rect 282 2748 302 2751
rect 6 2742 9 2748
rect 10 2738 70 2741
rect 158 2741 161 2748
rect 434 2748 510 2751
rect 514 2748 521 2751
rect 570 2748 582 2751
rect 586 2748 638 2751
rect 858 2748 878 2751
rect 954 2748 958 2751
rect 1010 2748 1062 2751
rect 1146 2748 1174 2751
rect 1178 2748 1206 2751
rect 1242 2748 1254 2751
rect 1346 2748 1542 2751
rect 1546 2748 1574 2751
rect 1642 2748 1670 2751
rect 1674 2748 1798 2751
rect 1834 2748 1838 2751
rect 1882 2748 1926 2751
rect 138 2738 161 2741
rect 186 2738 246 2741
rect 398 2741 401 2748
rect 814 2742 817 2748
rect 330 2738 646 2741
rect 826 2738 870 2741
rect 882 2738 974 2741
rect 1078 2741 1081 2748
rect 1946 2748 2030 2751
rect 2086 2748 2102 2751
rect 2206 2751 2209 2758
rect 2358 2752 2361 2758
rect 2202 2748 2209 2751
rect 2234 2748 2313 2751
rect 2086 2742 2089 2748
rect 2158 2742 2161 2748
rect 2310 2742 2313 2748
rect 2394 2748 2542 2751
rect 2554 2748 2558 2751
rect 2610 2748 2630 2751
rect 2634 2748 3246 2751
rect 3394 2748 3430 2751
rect 3474 2748 3486 2751
rect 3506 2748 3518 2751
rect 3554 2748 3782 2751
rect 1050 2738 1081 2741
rect 1106 2738 1185 2741
rect 1194 2738 1214 2741
rect 1410 2738 1454 2741
rect 1474 2738 1486 2741
rect 1490 2738 1622 2741
rect 1714 2738 1718 2741
rect 1738 2738 1750 2741
rect 1770 2738 1774 2741
rect 1794 2738 1822 2741
rect 1890 2738 1990 2741
rect 2114 2738 2142 2741
rect 2194 2738 2254 2741
rect 2334 2741 2337 2748
rect 3794 2748 3806 2751
rect 3834 2748 3854 2751
rect 3858 2748 3894 2751
rect 3914 2748 3934 2751
rect 3938 2748 3942 2751
rect 3954 2748 3974 2751
rect 3978 2748 4014 2751
rect 4066 2748 4070 2751
rect 4090 2748 4118 2751
rect 4146 2748 4526 2751
rect 4746 2748 4758 2751
rect 4834 2748 5070 2751
rect 5222 2751 5226 2752
rect 5122 2748 5226 2751
rect 2334 2738 2382 2741
rect 2386 2738 2393 2741
rect 2482 2738 2758 2741
rect 2762 2738 2857 2741
rect 2874 2738 2878 2741
rect 2890 2738 2942 2741
rect 2998 2738 3022 2741
rect 3026 2738 3054 2741
rect 3090 2738 3286 2741
rect 3290 2738 3369 2741
rect 3498 2738 3534 2741
rect 3538 2738 3694 2741
rect 3698 2738 3782 2741
rect 3794 2738 3798 2741
rect 3834 2738 3862 2741
rect 3906 2738 3958 2741
rect 3986 2738 4062 2741
rect 4234 2738 4398 2741
rect 4582 2741 4585 2748
rect 4678 2742 4681 2748
rect 4582 2738 4606 2741
rect 4690 2738 4734 2741
rect 4738 2738 4742 2741
rect 4822 2741 4825 2748
rect 4822 2738 4886 2741
rect 4890 2738 4958 2741
rect 4994 2738 5014 2741
rect 1182 2732 1185 2738
rect 2038 2732 2041 2738
rect 574 2728 798 2731
rect 818 2728 822 2731
rect 846 2728 862 2731
rect 1266 2728 1422 2731
rect 1506 2728 1630 2731
rect 1714 2728 1750 2731
rect 1762 2728 1774 2731
rect 1826 2728 1878 2731
rect 1882 2728 1921 2731
rect 1986 2728 2006 2731
rect 2182 2731 2185 2738
rect 2854 2732 2857 2738
rect 2998 2732 3001 2738
rect 3286 2732 3289 2738
rect 3366 2732 3369 2738
rect 2162 2728 2185 2731
rect 2226 2728 2246 2731
rect 2274 2728 2334 2731
rect 2354 2728 2430 2731
rect 2546 2728 2566 2731
rect 2706 2728 2718 2731
rect 2722 2728 2774 2731
rect 2878 2728 2966 2731
rect 3010 2728 3118 2731
rect 3130 2728 3214 2731
rect 3546 2728 3630 2731
rect 3650 2728 3678 2731
rect 3698 2728 3726 2731
rect 3810 2728 3870 2731
rect 3898 2728 3950 2731
rect 4010 2728 4022 2731
rect 4034 2728 4070 2731
rect 4074 2728 4177 2731
rect 4186 2728 4254 2731
rect 4258 2728 4414 2731
rect 4466 2728 4558 2731
rect 4578 2728 4582 2731
rect 4594 2728 4606 2731
rect 4682 2728 4806 2731
rect 4826 2728 4838 2731
rect 4906 2728 4910 2731
rect 4962 2728 5118 2731
rect 574 2722 577 2728
rect 314 2718 350 2721
rect 354 2718 502 2721
rect 838 2721 841 2728
rect 746 2718 841 2721
rect 846 2722 849 2728
rect 1918 2722 1921 2728
rect 2846 2722 2849 2728
rect 2878 2722 2881 2728
rect 954 2718 1046 2721
rect 1434 2718 1534 2721
rect 1714 2718 1814 2721
rect 1818 2718 1894 2721
rect 1938 2718 2118 2721
rect 2122 2718 2350 2721
rect 2354 2718 2558 2721
rect 2770 2718 2838 2721
rect 3074 2718 3518 2721
rect 3530 2718 3590 2721
rect 3594 2718 3662 2721
rect 3686 2721 3689 2728
rect 3686 2718 3838 2721
rect 3850 2718 3910 2721
rect 3922 2718 3926 2721
rect 4174 2721 4177 2728
rect 4174 2718 4254 2721
rect 4258 2718 4326 2721
rect 4422 2721 4425 2728
rect 4402 2718 4425 2721
rect 4458 2718 4598 2721
rect 4602 2718 4702 2721
rect 4866 2718 4926 2721
rect 586 2708 854 2711
rect 858 2708 998 2711
rect 1162 2708 1198 2711
rect 1258 2708 1278 2711
rect 1354 2708 1358 2711
rect 1362 2708 1406 2711
rect 1442 2708 1649 2711
rect 1858 2708 1942 2711
rect 2210 2708 2838 2711
rect 2850 2708 3006 2711
rect 3122 2708 3142 2711
rect 3202 2708 3406 2711
rect 3410 2708 3430 2711
rect 3562 2708 3758 2711
rect 3762 2708 3782 2711
rect 3890 2708 3894 2711
rect 4082 2708 4102 2711
rect 4162 2708 4542 2711
rect 4722 2708 4750 2711
rect 5066 2708 5086 2711
rect 1048 2703 1050 2707
rect 1054 2703 1057 2707
rect 1062 2703 1064 2707
rect 130 2698 214 2701
rect 450 2698 697 2701
rect 706 2698 1030 2701
rect 1074 2698 1166 2701
rect 1434 2698 1494 2701
rect 1498 2698 1582 2701
rect 1646 2701 1649 2708
rect 2072 2703 2074 2707
rect 2078 2703 2081 2707
rect 2086 2703 2088 2707
rect 3096 2703 3098 2707
rect 3102 2703 3105 2707
rect 3110 2703 3112 2707
rect 4112 2703 4114 2707
rect 4118 2703 4121 2707
rect 4126 2703 4128 2707
rect 1646 2698 2054 2701
rect 2210 2698 2262 2701
rect 2354 2698 2366 2701
rect 2378 2698 2422 2701
rect 2434 2698 2478 2701
rect 2530 2698 2542 2701
rect 2618 2698 2686 2701
rect 2826 2698 2870 2701
rect 3066 2698 3078 2701
rect 3122 2698 3182 2701
rect 3218 2698 3302 2701
rect 3562 2698 3582 2701
rect 3714 2698 3910 2701
rect 3930 2698 3998 2701
rect 4138 2698 4398 2701
rect 4402 2698 4958 2701
rect 186 2688 358 2691
rect 378 2688 470 2691
rect 578 2688 582 2691
rect 694 2691 697 2698
rect 694 2688 710 2691
rect 906 2688 1718 2691
rect 1722 2688 1838 2691
rect 1842 2688 2974 2691
rect 2978 2688 3662 2691
rect 3682 2688 3806 2691
rect 3914 2688 3942 2691
rect 4010 2688 4286 2691
rect 4298 2688 4318 2691
rect 4330 2688 4425 2691
rect 4594 2688 4622 2691
rect 4666 2688 4774 2691
rect 5002 2688 5110 2691
rect 5114 2688 5134 2691
rect 4422 2682 4425 2688
rect 194 2678 206 2681
rect 226 2678 702 2681
rect 722 2678 838 2681
rect 882 2678 982 2681
rect 1050 2678 1086 2681
rect 1506 2678 1550 2681
rect 1746 2678 1750 2681
rect 1810 2678 1822 2681
rect 1826 2678 1838 2681
rect 1898 2678 1934 2681
rect 1954 2678 2022 2681
rect 2082 2678 2110 2681
rect 2242 2678 2246 2681
rect 2258 2678 2374 2681
rect 2498 2678 2534 2681
rect 2562 2678 2766 2681
rect 3058 2678 3070 2681
rect 3102 2678 3126 2681
rect 3314 2678 3334 2681
rect 3338 2678 3534 2681
rect 3586 2678 3646 2681
rect 3674 2678 3718 2681
rect 3746 2678 3798 2681
rect 3810 2678 3894 2681
rect 3898 2678 3934 2681
rect 3938 2678 4062 2681
rect 4066 2678 4086 2681
rect 4230 2678 4366 2681
rect 4618 2678 4686 2681
rect 4946 2678 4966 2681
rect 4970 2678 4982 2681
rect 42 2668 118 2671
rect 154 2668 206 2671
rect 266 2668 270 2671
rect 338 2668 350 2671
rect 410 2668 510 2671
rect 682 2668 686 2671
rect 738 2668 1030 2671
rect 1118 2671 1121 2678
rect 1082 2668 1121 2671
rect 1366 2671 1369 2678
rect 1414 2672 1417 2678
rect 1446 2672 1449 2678
rect 1366 2668 1374 2671
rect 1402 2668 1406 2671
rect 1506 2668 1510 2671
rect 1658 2668 1678 2671
rect 1698 2668 1710 2671
rect 1730 2668 1750 2671
rect 1866 2668 1998 2671
rect 2026 2668 2046 2671
rect 2190 2671 2193 2678
rect 2854 2672 2857 2678
rect 2190 2668 2302 2671
rect 2810 2668 2830 2671
rect 2874 2668 2878 2671
rect 2882 2668 2894 2671
rect 3102 2671 3105 2678
rect 4230 2672 4233 2678
rect 2922 2668 3105 2671
rect 3114 2668 3358 2671
rect 3394 2668 3518 2671
rect 3522 2668 3598 2671
rect 3690 2668 3726 2671
rect 3778 2668 3886 2671
rect 3930 2668 4142 2671
rect 4338 2668 4350 2671
rect 4378 2668 4446 2671
rect 4490 2668 4518 2671
rect 4522 2668 4566 2671
rect 4594 2668 4646 2671
rect 4674 2668 4678 2671
rect 4774 2671 4777 2678
rect 4774 2668 4870 2671
rect 4874 2668 4878 2671
rect 5022 2671 5025 2678
rect 5022 2668 5054 2671
rect 5074 2668 5078 2671
rect 130 2658 142 2661
rect 242 2658 270 2661
rect 274 2658 294 2661
rect 366 2661 369 2668
rect 1030 2662 1033 2668
rect 366 2658 478 2661
rect 482 2658 814 2661
rect 834 2658 838 2661
rect 842 2658 982 2661
rect 986 2658 1014 2661
rect 1066 2658 1089 2661
rect 1106 2658 1166 2661
rect 1170 2658 1198 2661
rect 1238 2661 1241 2668
rect 1246 2661 1249 2668
rect 2102 2662 2105 2668
rect 2358 2662 2361 2668
rect 2374 2662 2377 2668
rect 2382 2662 2385 2668
rect 1238 2658 1249 2661
rect 1258 2658 1294 2661
rect 1386 2658 1406 2661
rect 1434 2658 1470 2661
rect 1474 2658 1774 2661
rect 1802 2658 1934 2661
rect 1938 2658 1950 2661
rect 1970 2658 2006 2661
rect 2042 2658 2078 2661
rect 2146 2658 2150 2661
rect 2170 2658 2222 2661
rect 2226 2658 2270 2661
rect 2282 2658 2334 2661
rect 2338 2658 2350 2661
rect 2414 2661 2417 2668
rect 2462 2661 2465 2668
rect 2414 2658 2465 2661
rect 2598 2661 2601 2668
rect 3678 2662 3681 2668
rect 2598 2658 2662 2661
rect 2698 2658 2702 2661
rect 2730 2658 2886 2661
rect 2906 2658 2926 2661
rect 3002 2658 3038 2661
rect 3090 2658 3382 2661
rect 3386 2658 3486 2661
rect 3490 2658 3566 2661
rect 3594 2658 3606 2661
rect 3610 2658 3670 2661
rect 3774 2658 3782 2661
rect 3786 2658 3846 2661
rect 3938 2658 3942 2661
rect 3946 2658 4006 2661
rect 4018 2658 4142 2661
rect 4194 2658 4206 2661
rect 4290 2658 4358 2661
rect 4386 2658 4510 2661
rect 4586 2658 4958 2661
rect 4962 2658 4974 2661
rect 4978 2658 4982 2661
rect 4986 2658 4998 2661
rect 5018 2658 5022 2661
rect 5170 2658 5182 2661
rect 190 2652 193 2658
rect 1086 2652 1089 2658
rect 3086 2652 3089 2658
rect 3694 2652 3697 2658
rect 5142 2652 5145 2658
rect -26 2651 -22 2652
rect -26 2648 158 2651
rect 234 2648 326 2651
rect 498 2648 526 2651
rect 530 2648 558 2651
rect 562 2648 582 2651
rect 650 2648 654 2651
rect 802 2648 849 2651
rect 874 2648 894 2651
rect 954 2648 993 2651
rect 1098 2648 1134 2651
rect 1154 2648 1270 2651
rect 1298 2648 1374 2651
rect 1378 2648 1385 2651
rect 1394 2648 1414 2651
rect 1434 2648 1462 2651
rect 1466 2648 1478 2651
rect 1530 2648 1726 2651
rect 1738 2648 1822 2651
rect 2002 2648 2041 2651
rect 2258 2648 2262 2651
rect 2298 2648 2302 2651
rect 2398 2648 2406 2651
rect 2410 2648 2526 2651
rect 2546 2648 2718 2651
rect 2786 2648 2790 2651
rect 2826 2648 2862 2651
rect 2898 2648 2910 2651
rect 3170 2648 3174 2651
rect 3298 2648 3318 2651
rect 3354 2648 3366 2651
rect 3390 2648 3430 2651
rect 3482 2648 3542 2651
rect 3906 2648 4014 2651
rect 4058 2648 4246 2651
rect 4402 2648 4518 2651
rect 4522 2648 4566 2651
rect 4650 2648 4670 2651
rect 4690 2648 5038 2651
rect 5058 2648 5062 2651
rect 5222 2651 5226 2652
rect 5194 2648 5226 2651
rect 846 2642 849 2648
rect 990 2642 993 2648
rect 578 2638 678 2641
rect 998 2638 2030 2641
rect 2038 2641 2041 2648
rect 3390 2642 3393 2648
rect 3566 2642 3569 2648
rect 2038 2638 2702 2641
rect 3162 2638 3318 2641
rect 3482 2638 3561 2641
rect 3682 2638 3790 2641
rect 3810 2638 4182 2641
rect 4330 2638 4438 2641
rect 4458 2638 4478 2641
rect 4566 2641 4569 2648
rect 5166 2642 5169 2648
rect 4566 2638 4790 2641
rect 4794 2638 5110 2641
rect 998 2632 1001 2638
rect 538 2628 670 2631
rect 810 2628 902 2631
rect 1474 2628 1766 2631
rect 1882 2628 1958 2631
rect 1962 2628 2054 2631
rect 2074 2628 2246 2631
rect 2394 2628 2406 2631
rect 2594 2628 2742 2631
rect 3134 2628 3142 2631
rect 3146 2628 3334 2631
rect 3466 2628 3550 2631
rect 3558 2631 3561 2638
rect 3558 2628 3574 2631
rect 3578 2628 3590 2631
rect 3642 2628 3694 2631
rect 3954 2628 4238 2631
rect 4806 2628 4942 2631
rect 274 2618 438 2621
rect 594 2618 606 2621
rect 610 2618 694 2621
rect 726 2621 729 2628
rect 726 2618 766 2621
rect 786 2618 918 2621
rect 934 2621 937 2628
rect 4806 2622 4809 2628
rect 934 2618 1070 2621
rect 1218 2618 1438 2621
rect 1570 2618 1574 2621
rect 1586 2618 1606 2621
rect 1610 2618 1830 2621
rect 1834 2618 2046 2621
rect 2066 2618 2374 2621
rect 2378 2618 2454 2621
rect 2458 2618 2534 2621
rect 2570 2618 2862 2621
rect 2882 2618 3110 2621
rect 3138 2618 3478 2621
rect 3554 2618 3654 2621
rect 3722 2618 3782 2621
rect 3794 2618 4094 2621
rect 4162 2618 4214 2621
rect 4450 2618 4686 2621
rect 4698 2618 4806 2621
rect 4834 2618 4838 2621
rect 4922 2618 4934 2621
rect 5082 2618 5142 2621
rect 754 2608 830 2611
rect 1002 2608 1006 2611
rect 1178 2608 1198 2611
rect 1234 2608 1390 2611
rect 1666 2608 1734 2611
rect 1742 2608 1990 2611
rect 2058 2608 2462 2611
rect 2962 2608 2966 2611
rect 2986 2608 3174 2611
rect 3178 2608 3198 2611
rect 3234 2608 3566 2611
rect 3674 2608 3742 2611
rect 3746 2608 3750 2611
rect 3978 2608 4046 2611
rect 4074 2608 4278 2611
rect 4450 2608 4574 2611
rect 4658 2608 4750 2611
rect 536 2603 538 2607
rect 542 2603 545 2607
rect 550 2603 552 2607
rect 1560 2603 1562 2607
rect 1566 2603 1569 2607
rect 1574 2603 1576 2607
rect 194 2598 342 2601
rect 730 2598 758 2601
rect 778 2598 782 2601
rect 794 2598 806 2601
rect 938 2598 1142 2601
rect 1186 2598 1286 2601
rect 1290 2598 1422 2601
rect 1450 2598 1542 2601
rect 1602 2598 1702 2601
rect 1742 2601 1745 2608
rect 2584 2603 2586 2607
rect 2590 2603 2593 2607
rect 2598 2603 2600 2607
rect 3608 2603 3610 2607
rect 3614 2603 3617 2607
rect 3622 2603 3624 2607
rect 3790 2602 3793 2608
rect 4632 2603 4634 2607
rect 4638 2603 4641 2607
rect 4646 2603 4648 2607
rect 1714 2598 1745 2601
rect 1938 2598 1950 2601
rect 1978 2598 2030 2601
rect 2074 2598 2241 2601
rect 2274 2598 2294 2601
rect 2658 2598 2862 2601
rect 3082 2598 3350 2601
rect 3362 2598 3598 2601
rect 3634 2598 3742 2601
rect 3794 2598 3814 2601
rect 4042 2598 4062 2601
rect 4070 2598 4622 2601
rect 4866 2598 5102 2601
rect 1862 2592 1865 2598
rect 258 2588 318 2591
rect 322 2588 622 2591
rect 722 2588 1022 2591
rect 1026 2588 1846 2591
rect 1898 2588 1918 2591
rect 1938 2588 2230 2591
rect 2238 2591 2241 2598
rect 2238 2588 2302 2591
rect 2338 2588 2366 2591
rect 2394 2588 2510 2591
rect 2538 2588 2622 2591
rect 2666 2588 2702 2591
rect 2794 2588 2870 2591
rect 2962 2588 3030 2591
rect 3322 2588 3534 2591
rect 3546 2588 3606 2591
rect 3682 2588 3806 2591
rect 4070 2591 4073 2598
rect 3814 2588 4073 2591
rect 4098 2588 4206 2591
rect 4226 2588 4310 2591
rect 4314 2588 5126 2591
rect 298 2578 390 2581
rect 394 2578 430 2581
rect 434 2578 790 2581
rect 794 2578 822 2581
rect 826 2578 862 2581
rect 866 2578 902 2581
rect 914 2578 1070 2581
rect 1162 2578 1166 2581
rect 1194 2578 1686 2581
rect 1802 2578 1838 2581
rect 1850 2578 2022 2581
rect 2058 2578 2238 2581
rect 2250 2578 2294 2581
rect 2298 2578 2398 2581
rect 2402 2578 2502 2581
rect 2506 2578 3014 2581
rect 3274 2578 3534 2581
rect 3594 2578 3678 2581
rect 3814 2581 3817 2588
rect 4766 2582 4769 2588
rect 3778 2578 3817 2581
rect 3866 2578 3918 2581
rect 3922 2578 4014 2581
rect 4026 2578 4382 2581
rect 4474 2578 4574 2581
rect 4578 2578 4742 2581
rect 5010 2578 5118 2581
rect 66 2568 166 2571
rect 170 2568 294 2571
rect 498 2568 502 2571
rect 538 2568 574 2571
rect 586 2568 742 2571
rect 786 2568 798 2571
rect 1082 2568 1094 2571
rect 1138 2568 1206 2571
rect 1354 2568 1486 2571
rect 1690 2568 2566 2571
rect 2650 2568 2686 2571
rect 2690 2568 2814 2571
rect 2850 2568 2854 2571
rect 2890 2568 2918 2571
rect 2922 2568 3014 2571
rect 3018 2568 3206 2571
rect 3394 2568 3526 2571
rect 3562 2568 3630 2571
rect 3634 2568 3950 2571
rect 3962 2568 4110 2571
rect 4202 2568 4294 2571
rect 4498 2568 4550 2571
rect 4586 2568 4638 2571
rect 4850 2568 4878 2571
rect 4930 2568 4934 2571
rect 4938 2568 5102 2571
rect 5122 2568 5174 2571
rect 130 2558 142 2561
rect 146 2558 382 2561
rect 486 2561 489 2568
rect 486 2558 574 2561
rect 610 2558 814 2561
rect 1038 2561 1041 2568
rect 1002 2558 1041 2561
rect 1054 2558 1142 2561
rect 1282 2558 1374 2561
rect 1386 2558 1406 2561
rect 1486 2558 1494 2561
rect 1498 2558 1510 2561
rect 1530 2558 1670 2561
rect 1674 2558 1702 2561
rect 1842 2558 2022 2561
rect 2026 2558 2318 2561
rect 2322 2558 2326 2561
rect 2386 2558 2414 2561
rect 2442 2558 2454 2561
rect 2562 2558 2598 2561
rect 2602 2558 2630 2561
rect 2778 2558 2814 2561
rect 2834 2558 2886 2561
rect 2930 2558 2934 2561
rect 2938 2558 3086 2561
rect 3362 2558 3382 2561
rect 3458 2558 3494 2561
rect 3510 2558 3518 2561
rect 3522 2558 3550 2561
rect 3570 2558 3686 2561
rect 3718 2558 3750 2561
rect 3842 2558 4150 2561
rect 4154 2558 4158 2561
rect 4394 2558 4430 2561
rect 4466 2558 4582 2561
rect 4602 2558 4702 2561
rect 4786 2558 4910 2561
rect 5114 2558 5126 2561
rect -26 2551 -22 2552
rect -26 2548 6 2551
rect 50 2548 102 2551
rect 210 2548 270 2551
rect 318 2548 401 2551
rect 426 2548 590 2551
rect 642 2548 646 2551
rect 774 2548 790 2551
rect 814 2551 817 2558
rect 810 2548 817 2551
rect 846 2552 849 2558
rect 1054 2552 1057 2558
rect 858 2548 918 2551
rect 1018 2548 1030 2551
rect 1162 2548 1166 2551
rect 1190 2551 1193 2558
rect 1190 2548 1214 2551
rect 1242 2548 1342 2551
rect 1414 2548 1422 2551
rect 1474 2548 1478 2551
rect 1490 2548 1494 2551
rect 1502 2548 1510 2551
rect 1822 2551 1825 2558
rect 2334 2552 2337 2558
rect 1674 2548 1830 2551
rect 1858 2548 1894 2551
rect 1930 2548 1934 2551
rect 1954 2548 1990 2551
rect 2010 2548 2014 2551
rect 2050 2548 2062 2551
rect 2090 2548 2102 2551
rect 2146 2548 2150 2551
rect 2162 2548 2294 2551
rect 2354 2548 2358 2551
rect 2402 2548 2558 2551
rect 2562 2548 2662 2551
rect 2694 2551 2697 2558
rect 2694 2548 2710 2551
rect 2746 2548 2750 2551
rect 2762 2548 2774 2551
rect 2826 2548 2846 2551
rect 2858 2548 2894 2551
rect 2898 2548 2950 2551
rect 2970 2548 2974 2551
rect 318 2542 321 2548
rect 398 2542 401 2548
rect 482 2538 486 2541
rect 514 2538 518 2541
rect 562 2538 582 2541
rect 742 2541 745 2548
rect 626 2538 745 2541
rect 774 2542 777 2548
rect 834 2538 870 2541
rect 890 2538 1014 2541
rect 1082 2538 1110 2541
rect 1154 2538 1158 2541
rect 1182 2541 1185 2548
rect 1414 2542 1417 2548
rect 1430 2542 1433 2548
rect 1502 2542 1505 2548
rect 1182 2538 1198 2541
rect 1202 2538 1230 2541
rect 1306 2538 1321 2541
rect 1450 2538 1454 2541
rect 1466 2538 1478 2541
rect 1574 2541 1577 2548
rect 1530 2538 1577 2541
rect 1662 2542 1665 2548
rect 1990 2542 1993 2548
rect 1746 2538 1782 2541
rect 1786 2538 1838 2541
rect 1890 2538 1894 2541
rect 1922 2538 1942 2541
rect 1998 2541 2001 2548
rect 3130 2548 3190 2551
rect 3334 2551 3337 2558
rect 3322 2548 3337 2551
rect 3490 2548 3502 2551
rect 3634 2548 3646 2551
rect 3710 2551 3713 2558
rect 3698 2548 3713 2551
rect 3718 2552 3721 2558
rect 3818 2548 3902 2551
rect 4074 2548 4121 2551
rect 4130 2548 4134 2551
rect 4166 2551 4169 2558
rect 4162 2548 4169 2551
rect 4246 2551 4249 2558
rect 4194 2548 4249 2551
rect 4354 2548 4406 2551
rect 4614 2548 4622 2551
rect 4710 2551 4713 2558
rect 5126 2552 5129 2558
rect 5158 2552 5161 2558
rect 4626 2548 4713 2551
rect 4762 2548 4766 2551
rect 4810 2548 5062 2551
rect 1998 2538 2057 2541
rect 2114 2538 2262 2541
rect 2282 2538 2622 2541
rect 2654 2538 2678 2541
rect 2706 2538 3006 2541
rect 3222 2541 3225 2548
rect 3454 2542 3457 2548
rect 3150 2538 3230 2541
rect 3330 2538 3358 2541
rect 3378 2538 3382 2541
rect 3466 2538 3486 2541
rect 3518 2541 3521 2548
rect 3518 2538 3646 2541
rect 3650 2538 3686 2541
rect 3746 2538 3774 2541
rect 3778 2538 3838 2541
rect 3850 2538 4102 2541
rect 4118 2541 4121 2548
rect 4526 2542 4529 2548
rect 4598 2542 4601 2548
rect 4118 2538 4142 2541
rect 4330 2538 4334 2541
rect 4362 2538 4390 2541
rect 4394 2538 4446 2541
rect 4578 2538 4590 2541
rect 4602 2538 4614 2541
rect 4618 2538 4798 2541
rect 4802 2538 4814 2541
rect 4978 2538 5102 2541
rect 5110 2541 5113 2548
rect 5106 2538 5113 2541
rect 5130 2538 5150 2541
rect 142 2531 145 2538
rect 1318 2532 1321 2538
rect 1494 2532 1497 2538
rect 2054 2532 2057 2538
rect 2654 2532 2657 2538
rect 114 2528 145 2531
rect 474 2528 494 2531
rect 506 2528 638 2531
rect 642 2528 686 2531
rect 874 2528 878 2531
rect 930 2528 1030 2531
rect 1042 2528 1134 2531
rect 1138 2528 1182 2531
rect 1234 2528 1238 2531
rect 1370 2528 1390 2531
rect 1394 2528 1470 2531
rect 1706 2528 1822 2531
rect 1962 2528 1990 2531
rect 2110 2528 2134 2531
rect 2218 2528 2273 2531
rect 2338 2528 2350 2531
rect 2370 2528 2574 2531
rect 2578 2528 2630 2531
rect 2698 2528 2750 2531
rect 2762 2528 2862 2531
rect 2914 2528 2966 2531
rect 3022 2531 3025 2538
rect 3150 2532 3153 2538
rect 3286 2532 3289 2538
rect 3022 2528 3086 2531
rect 3210 2528 3214 2531
rect 3298 2528 3334 2531
rect 3466 2528 3478 2531
rect 3586 2528 3670 2531
rect 3818 2528 3830 2531
rect 3834 2528 3950 2531
rect 3954 2528 4022 2531
rect 4058 2528 4086 2531
rect 4218 2528 4310 2531
rect 4370 2528 4494 2531
rect 4546 2528 4734 2531
rect 4778 2528 4782 2531
rect 4794 2528 4814 2531
rect 5098 2528 5134 2531
rect 5138 2528 5158 2531
rect 106 2518 150 2521
rect 386 2518 414 2521
rect 418 2518 478 2521
rect 522 2518 614 2521
rect 798 2521 801 2528
rect 2110 2522 2113 2528
rect 798 2518 902 2521
rect 922 2518 1862 2521
rect 1938 2518 1942 2521
rect 1946 2518 1950 2521
rect 2010 2518 2022 2521
rect 2042 2518 2046 2521
rect 2150 2521 2153 2528
rect 2150 2518 2158 2521
rect 2210 2518 2214 2521
rect 2242 2518 2262 2521
rect 2270 2521 2273 2528
rect 2270 2518 2278 2521
rect 2346 2518 2438 2521
rect 2514 2518 2574 2521
rect 2578 2518 2585 2521
rect 2594 2518 2686 2521
rect 2690 2518 2726 2521
rect 2730 2518 2822 2521
rect 2842 2518 2846 2521
rect 2906 2518 2918 2521
rect 3006 2521 3009 2528
rect 3334 2522 3337 2528
rect 3006 2518 3046 2521
rect 3050 2518 3166 2521
rect 3186 2518 3326 2521
rect 3342 2518 3430 2521
rect 3530 2518 4246 2521
rect 4250 2518 4342 2521
rect 4846 2521 4849 2528
rect 4586 2518 4849 2521
rect 4894 2521 4897 2528
rect 4894 2518 4966 2521
rect 5002 2518 5150 2521
rect -26 2511 -22 2512
rect -26 2508 14 2511
rect 138 2508 246 2511
rect 426 2508 454 2511
rect 570 2508 630 2511
rect 650 2508 758 2511
rect 762 2508 934 2511
rect 1122 2508 1262 2511
rect 1354 2508 1374 2511
rect 1402 2508 1574 2511
rect 1658 2508 1678 2511
rect 1690 2508 1726 2511
rect 1746 2508 1750 2511
rect 1834 2508 1990 2511
rect 1994 2508 2030 2511
rect 2034 2508 2062 2511
rect 2106 2508 2150 2511
rect 2170 2508 2198 2511
rect 2202 2508 2302 2511
rect 2386 2508 2534 2511
rect 2714 2508 2742 2511
rect 2786 2508 2806 2511
rect 2922 2508 3086 2511
rect 3342 2511 3345 2518
rect 3314 2508 3345 2511
rect 3354 2508 3390 2511
rect 3474 2508 3862 2511
rect 3922 2508 4006 2511
rect 4010 2508 4054 2511
rect 4162 2508 4174 2511
rect 4178 2508 4190 2511
rect 4194 2508 4198 2511
rect 4342 2511 4345 2518
rect 4342 2508 5038 2511
rect 5042 2508 5150 2511
rect 1048 2503 1050 2507
rect 1054 2503 1057 2507
rect 1062 2503 1064 2507
rect 2072 2503 2074 2507
rect 2078 2503 2081 2507
rect 2086 2503 2088 2507
rect 3096 2503 3098 2507
rect 3102 2503 3105 2507
rect 3110 2503 3112 2507
rect 4112 2503 4114 2507
rect 4118 2503 4121 2507
rect 4126 2503 4128 2507
rect 154 2498 622 2501
rect 666 2498 702 2501
rect 714 2498 918 2501
rect 1130 2498 1158 2501
rect 1186 2498 1358 2501
rect 1434 2498 1510 2501
rect 1690 2498 1710 2501
rect 1714 2498 1902 2501
rect 1938 2498 2046 2501
rect 2210 2498 2214 2501
rect 2242 2498 2446 2501
rect 2522 2498 2694 2501
rect 2706 2498 2742 2501
rect 2806 2498 2902 2501
rect 2938 2498 2950 2501
rect 2986 2498 3046 2501
rect 3138 2498 3158 2501
rect 3202 2498 3310 2501
rect 3338 2498 3366 2501
rect 3402 2498 3430 2501
rect 3546 2498 3609 2501
rect 1542 2492 1545 2498
rect -26 2491 -22 2492
rect -26 2488 6 2491
rect 26 2488 142 2491
rect 250 2488 270 2491
rect 274 2488 334 2491
rect 338 2488 446 2491
rect 450 2488 502 2491
rect 634 2488 798 2491
rect 810 2488 814 2491
rect 1018 2488 1054 2491
rect 1058 2488 1262 2491
rect 1306 2488 1358 2491
rect 1410 2488 1470 2491
rect 1482 2488 1526 2491
rect 1562 2488 1598 2491
rect 1602 2488 1670 2491
rect 1674 2488 1694 2491
rect 1746 2488 1758 2491
rect 1786 2488 1798 2491
rect 1810 2488 1814 2491
rect 1826 2488 1894 2491
rect 1914 2488 1966 2491
rect 1970 2488 2014 2491
rect 2018 2488 2118 2491
rect 2122 2488 2193 2491
rect 2226 2488 2494 2491
rect 2538 2488 2654 2491
rect 2806 2491 2809 2498
rect 2682 2488 2809 2491
rect 2970 2488 3006 2491
rect 3066 2488 3070 2491
rect 3082 2488 3206 2491
rect 3218 2488 3262 2491
rect 3266 2488 3273 2491
rect 3282 2488 3294 2491
rect 3362 2488 3366 2491
rect 3386 2488 3462 2491
rect 3466 2488 3473 2491
rect 3482 2488 3486 2491
rect 3490 2488 3582 2491
rect 3586 2488 3590 2491
rect 3606 2491 3609 2498
rect 3646 2498 3662 2501
rect 3674 2498 3742 2501
rect 3754 2498 3958 2501
rect 3978 2498 4078 2501
rect 4138 2498 4214 2501
rect 4218 2498 4342 2501
rect 4434 2498 4486 2501
rect 4530 2498 4534 2501
rect 4538 2498 4558 2501
rect 4570 2498 4750 2501
rect 4986 2498 5009 2501
rect 5050 2498 5174 2501
rect 3646 2491 3649 2498
rect 4102 2492 4105 2498
rect 3606 2488 3649 2491
rect 3706 2488 3766 2491
rect 3802 2488 3934 2491
rect 3938 2488 4086 2491
rect 4266 2488 4342 2491
rect 4426 2488 4454 2491
rect 4482 2488 4550 2491
rect 4558 2488 4630 2491
rect 4650 2488 4734 2491
rect 4746 2488 4782 2491
rect 4842 2488 4998 2491
rect 5006 2491 5009 2498
rect 5182 2492 5185 2498
rect 5006 2488 5142 2491
rect 374 2482 377 2488
rect 426 2478 534 2481
rect 546 2478 550 2481
rect 594 2478 846 2481
rect 858 2478 870 2481
rect 890 2478 1158 2481
rect 1186 2478 1550 2481
rect 1554 2478 1582 2481
rect 1658 2478 1702 2481
rect 1706 2478 1726 2481
rect 1762 2478 1830 2481
rect 1842 2478 1854 2481
rect 1882 2478 1886 2481
rect 1930 2478 1950 2481
rect 2010 2478 2062 2481
rect 2098 2478 2182 2481
rect 2190 2481 2193 2488
rect 2190 2478 2246 2481
rect 2306 2478 2342 2481
rect 2346 2478 2393 2481
rect 2390 2472 2393 2478
rect 2434 2478 2510 2481
rect 2530 2478 2582 2481
rect 2642 2478 2646 2481
rect 2738 2478 2798 2481
rect 2826 2478 3446 2481
rect 3466 2478 4166 2481
rect 4274 2478 4470 2481
rect 4558 2481 4561 2488
rect 4482 2478 4561 2481
rect 4570 2478 4638 2481
rect 4642 2478 4830 2481
rect 4834 2478 4838 2481
rect 4866 2478 4878 2481
rect 4890 2478 4910 2481
rect 4978 2478 5118 2481
rect 2422 2472 2425 2478
rect -26 2471 -22 2472
rect -26 2468 14 2471
rect 474 2468 649 2471
rect 114 2459 118 2461
rect 110 2458 118 2459
rect 182 2461 185 2468
rect 138 2458 185 2461
rect 310 2461 313 2468
rect 266 2458 313 2461
rect 382 2461 385 2468
rect 646 2462 649 2468
rect 762 2468 766 2471
rect 834 2468 862 2471
rect 906 2468 950 2471
rect 954 2468 958 2471
rect 970 2468 1182 2471
rect 1234 2468 1278 2471
rect 1298 2468 1318 2471
rect 1402 2468 1662 2471
rect 1682 2468 1758 2471
rect 1770 2468 2246 2471
rect 2282 2468 2366 2471
rect 2402 2468 2406 2471
rect 2466 2468 2542 2471
rect 2566 2468 2582 2471
rect 2642 2468 2646 2471
rect 2706 2468 2710 2471
rect 2746 2468 2785 2471
rect 2818 2468 2846 2471
rect 3058 2468 3062 2471
rect 3130 2468 3134 2471
rect 3142 2468 3150 2471
rect 3154 2468 3174 2471
rect 3186 2468 3190 2471
rect 3242 2468 3246 2471
rect 3322 2468 3846 2471
rect 3858 2468 3910 2471
rect 3938 2468 3950 2471
rect 3978 2468 3982 2471
rect 4034 2468 4038 2471
rect 4098 2468 4113 2471
rect 4266 2468 4350 2471
rect 4362 2468 4374 2471
rect 4378 2468 4398 2471
rect 4418 2468 4430 2471
rect 4434 2468 4446 2471
rect 4450 2468 4662 2471
rect 4754 2468 4846 2471
rect 4850 2468 4854 2471
rect 5114 2468 5174 2471
rect 382 2458 406 2461
rect 410 2458 430 2461
rect 538 2458 590 2461
rect 602 2458 606 2461
rect 702 2461 705 2468
rect 666 2458 705 2461
rect 806 2462 809 2468
rect 898 2458 905 2461
rect 914 2458 1038 2461
rect 1042 2458 1246 2461
rect 1258 2458 1502 2461
rect 1506 2458 1550 2461
rect 1554 2458 1614 2461
rect 1626 2458 1710 2461
rect 1738 2458 1750 2461
rect 1794 2458 1798 2461
rect 1866 2458 1870 2461
rect 1906 2458 1910 2461
rect 2010 2458 2118 2461
rect 2130 2458 2166 2461
rect 2202 2458 2230 2461
rect 2254 2461 2257 2468
rect 2566 2462 2569 2468
rect 2254 2458 2270 2461
rect 2362 2458 2382 2461
rect 2386 2458 2430 2461
rect 2454 2458 2462 2461
rect 2482 2458 2486 2461
rect 2598 2461 2601 2468
rect 2598 2458 2614 2461
rect 2686 2461 2689 2468
rect 2686 2458 2694 2461
rect 2714 2458 2742 2461
rect 2770 2458 2777 2461
rect 830 2452 833 2458
rect 838 2452 841 2458
rect -26 2451 -22 2452
rect -26 2448 30 2451
rect 234 2448 302 2451
rect 306 2448 398 2451
rect 578 2448 606 2451
rect 642 2448 662 2451
rect 706 2448 782 2451
rect 866 2448 886 2451
rect 902 2451 905 2458
rect 1878 2452 1881 2458
rect 1942 2452 1945 2458
rect 2318 2452 2321 2458
rect 2334 2452 2337 2458
rect 902 2448 982 2451
rect 1162 2448 1230 2451
rect 1266 2448 1286 2451
rect 1346 2448 1454 2451
rect 1474 2448 1806 2451
rect 1814 2448 1830 2451
rect 1846 2448 1870 2451
rect 1970 2448 2030 2451
rect 2074 2448 2206 2451
rect 2210 2448 2222 2451
rect 2298 2448 2310 2451
rect 2430 2448 2438 2451
rect 2454 2451 2457 2458
rect 2442 2448 2457 2451
rect 2510 2451 2513 2458
rect 2774 2452 2777 2458
rect 2782 2452 2785 2468
rect 2802 2458 2934 2461
rect 2954 2458 3014 2461
rect 3042 2458 3078 2461
rect 3082 2458 3150 2461
rect 3154 2458 3198 2461
rect 3202 2458 3254 2461
rect 3266 2458 3270 2461
rect 3306 2458 3310 2461
rect 3346 2458 3390 2461
rect 3410 2458 3414 2461
rect 3442 2458 3462 2461
rect 3514 2458 3526 2461
rect 3538 2458 3550 2461
rect 3626 2458 3630 2461
rect 3674 2458 3702 2461
rect 3762 2458 3782 2461
rect 3814 2458 3982 2461
rect 3990 2461 3993 2468
rect 4110 2462 4113 2468
rect 4862 2462 4865 2468
rect 3990 2458 4006 2461
rect 4010 2458 4014 2461
rect 4018 2458 4046 2461
rect 4050 2458 4089 2461
rect 3022 2452 3025 2458
rect 3814 2452 3817 2458
rect 4086 2452 4089 2458
rect 4202 2458 4206 2461
rect 4314 2458 4326 2461
rect 4346 2458 4366 2461
rect 4370 2458 4438 2461
rect 4462 2458 4497 2461
rect 4514 2458 4518 2461
rect 4522 2458 4534 2461
rect 4550 2458 4598 2461
rect 4690 2458 4734 2461
rect 4874 2458 4894 2461
rect 4898 2458 4945 2461
rect 5122 2458 5142 2461
rect 4094 2452 4097 2458
rect 4462 2452 4465 2458
rect 4494 2452 4497 2458
rect 4550 2452 4553 2458
rect 4942 2452 4945 2458
rect 2466 2448 2513 2451
rect 2578 2448 2606 2451
rect 2618 2448 2694 2451
rect 2834 2448 2838 2451
rect 3066 2448 3102 2451
rect 3106 2448 3222 2451
rect 3258 2448 3310 2451
rect 3426 2448 3438 2451
rect 3586 2448 3598 2451
rect 3618 2448 3726 2451
rect 3866 2448 3902 2451
rect 3914 2448 3926 2451
rect 3954 2448 3958 2451
rect 4038 2448 4062 2451
rect 4162 2448 4337 2451
rect 4346 2448 4377 2451
rect 4546 2448 4550 2451
rect 4606 2448 4678 2451
rect 4706 2448 4750 2451
rect 4786 2448 4846 2451
rect 5026 2448 5126 2451
rect 5146 2448 5158 2451
rect 5162 2448 5174 2451
rect 1238 2442 1241 2448
rect 1814 2442 1817 2448
rect 1846 2442 1849 2448
rect 506 2438 1078 2441
rect 1098 2438 1214 2441
rect 1266 2438 1558 2441
rect 1594 2438 1702 2441
rect 1858 2438 1878 2441
rect 1906 2438 1926 2441
rect 1994 2438 2070 2441
rect 2154 2438 2166 2441
rect 2242 2438 2294 2441
rect 2306 2438 2326 2441
rect 2358 2438 2366 2441
rect 2370 2438 2398 2441
rect 2410 2438 2758 2441
rect 2762 2438 3142 2441
rect 3186 2438 3206 2441
rect 3238 2441 3241 2448
rect 3238 2438 3270 2441
rect 3290 2438 3302 2441
rect 3322 2438 3350 2441
rect 3386 2438 3390 2441
rect 3418 2438 3422 2441
rect 3562 2438 3614 2441
rect 3642 2438 3654 2441
rect 3734 2441 3737 2448
rect 3722 2438 3737 2441
rect 3766 2442 3769 2448
rect 4038 2442 4041 2448
rect 3794 2438 3822 2441
rect 3914 2438 3934 2441
rect 3938 2438 3945 2441
rect 3974 2438 3998 2441
rect 4086 2441 4089 2448
rect 4334 2442 4337 2448
rect 4374 2442 4377 2448
rect 4606 2442 4609 2448
rect 4086 2438 4150 2441
rect 4490 2438 4574 2441
rect 4794 2438 4878 2441
rect 4882 2438 5110 2441
rect 5114 2438 5126 2441
rect 218 2428 630 2431
rect 850 2428 1166 2431
rect 1170 2428 1302 2431
rect 1378 2428 1390 2431
rect 1426 2428 1750 2431
rect 1786 2428 1942 2431
rect 1970 2428 2110 2431
rect 2114 2428 2174 2431
rect 2186 2428 2294 2431
rect 2326 2431 2329 2438
rect 3974 2432 3977 2438
rect 2326 2428 2382 2431
rect 2434 2428 2614 2431
rect 2634 2428 2902 2431
rect 2906 2428 3382 2431
rect 3386 2428 3950 2431
rect 3994 2428 4510 2431
rect 4542 2428 4550 2431
rect 4554 2428 4590 2431
rect 4762 2428 4942 2431
rect 5098 2428 5150 2431
rect 346 2418 654 2421
rect 658 2418 718 2421
rect 782 2421 785 2428
rect 782 2418 1206 2421
rect 1226 2418 1374 2421
rect 1530 2418 1646 2421
rect 1806 2418 1854 2421
rect 1874 2418 2158 2421
rect 2186 2418 2678 2421
rect 2810 2418 3126 2421
rect 3146 2418 3414 2421
rect 3426 2418 3486 2421
rect 3490 2418 3590 2421
rect 3610 2418 3638 2421
rect 3666 2418 3694 2421
rect 3794 2418 3886 2421
rect 3890 2418 3982 2421
rect 3986 2418 4030 2421
rect 4162 2418 4222 2421
rect 4474 2418 4798 2421
rect 4802 2418 4822 2421
rect 4826 2418 4902 2421
rect 4906 2418 5166 2421
rect 5170 2418 5182 2421
rect 802 2408 886 2411
rect 1002 2408 1110 2411
rect 1178 2408 1254 2411
rect 1290 2408 1310 2411
rect 1322 2408 1414 2411
rect 1626 2408 1686 2411
rect 1806 2411 1809 2418
rect 1690 2408 1809 2411
rect 1842 2408 2150 2411
rect 2282 2408 2382 2411
rect 2506 2408 2550 2411
rect 2658 2408 2782 2411
rect 2802 2408 2838 2411
rect 3018 2408 3030 2411
rect 3034 2408 3110 2411
rect 3162 2408 3190 2411
rect 3210 2408 3278 2411
rect 3294 2408 3430 2411
rect 3450 2408 3582 2411
rect 3786 2408 3966 2411
rect 3970 2408 4070 2411
rect 4074 2408 4118 2411
rect 4122 2408 4166 2411
rect 4186 2408 4366 2411
rect 4658 2408 4854 2411
rect 536 2403 538 2407
rect 542 2403 545 2407
rect 550 2403 552 2407
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1574 2403 1576 2407
rect 2584 2403 2586 2407
rect 2590 2403 2593 2407
rect 2598 2403 2600 2407
rect 3294 2402 3297 2408
rect 3608 2403 3610 2407
rect 3614 2403 3617 2407
rect 3622 2403 3624 2407
rect 4632 2403 4634 2407
rect 4638 2403 4641 2407
rect 4646 2403 4648 2407
rect 602 2398 622 2401
rect 634 2398 1417 2401
rect 1810 2398 2158 2401
rect 2162 2398 2262 2401
rect 2290 2398 2446 2401
rect 2658 2398 3086 2401
rect 3090 2398 3182 2401
rect 3194 2398 3198 2401
rect 3258 2398 3294 2401
rect 3306 2398 3334 2401
rect 3370 2398 3569 2401
rect 3810 2398 3846 2401
rect 4074 2398 4382 2401
rect 4386 2398 4518 2401
rect 4986 2398 5030 2401
rect 130 2388 206 2391
rect 210 2388 470 2391
rect 482 2388 825 2391
rect 850 2388 854 2391
rect 946 2388 1174 2391
rect 1186 2388 1278 2391
rect 1290 2388 1406 2391
rect 1414 2391 1417 2398
rect 1414 2388 1606 2391
rect 1706 2388 1750 2391
rect 1834 2388 1902 2391
rect 1922 2388 1990 2391
rect 2138 2388 2142 2391
rect 2178 2388 2182 2391
rect 2474 2388 2926 2391
rect 2930 2388 2990 2391
rect 2994 2388 3022 2391
rect 3026 2388 3366 2391
rect 3402 2388 3422 2391
rect 3498 2388 3510 2391
rect 3566 2391 3569 2398
rect 3566 2388 3742 2391
rect 3746 2388 3758 2391
rect 3762 2388 3790 2391
rect 3802 2388 3806 2391
rect 3954 2388 4446 2391
rect 4450 2388 4470 2391
rect 4770 2388 4886 2391
rect 546 2378 558 2381
rect 570 2378 742 2381
rect 822 2381 825 2388
rect 822 2378 1254 2381
rect 1314 2378 1318 2381
rect 1354 2378 1366 2381
rect 1386 2378 1502 2381
rect 1546 2378 1702 2381
rect 1722 2378 2174 2381
rect 2178 2378 2214 2381
rect 2218 2378 2286 2381
rect 2290 2378 2470 2381
rect 2610 2378 2646 2381
rect 2738 2378 2822 2381
rect 3014 2378 3270 2381
rect 3274 2378 3406 2381
rect 3410 2378 3742 2381
rect 3746 2378 3790 2381
rect 3798 2378 3878 2381
rect 4018 2378 4238 2381
rect 4386 2378 4774 2381
rect 4798 2378 4854 2381
rect -26 2371 -22 2372
rect 6 2371 9 2378
rect 1278 2372 1281 2378
rect -26 2368 9 2371
rect 182 2368 270 2371
rect 274 2368 318 2371
rect 362 2368 382 2371
rect 434 2368 478 2371
rect 498 2368 526 2371
rect 530 2368 574 2371
rect 818 2368 846 2371
rect 906 2368 1198 2371
rect 1218 2368 1262 2371
rect 1290 2368 1358 2371
rect 1370 2368 1398 2371
rect 1458 2368 1558 2371
rect 1586 2368 1606 2371
rect 1638 2368 1646 2371
rect 1650 2368 1670 2371
rect 1826 2368 1862 2371
rect 1882 2368 1910 2371
rect 1930 2368 1934 2371
rect 2010 2368 2014 2371
rect 2018 2368 2046 2371
rect 2090 2368 2118 2371
rect 2146 2368 2166 2371
rect 2170 2368 2193 2371
rect 2250 2368 2334 2371
rect 2338 2368 2358 2371
rect 2362 2368 2502 2371
rect 2534 2371 2537 2378
rect 3014 2372 3017 2378
rect 2534 2368 2550 2371
rect 2570 2368 2614 2371
rect 2634 2368 2694 2371
rect 2714 2368 2998 2371
rect 3098 2368 3118 2371
rect 3234 2368 3374 2371
rect 3378 2368 3462 2371
rect 3466 2368 3542 2371
rect 3546 2368 3678 2371
rect 3798 2371 3801 2378
rect 3786 2368 3801 2371
rect 3898 2368 4182 2371
rect 4222 2368 4230 2371
rect 4234 2368 4278 2371
rect 4798 2371 4801 2378
rect 4522 2368 4801 2371
rect 4938 2368 5038 2371
rect 5050 2368 5086 2371
rect 166 2361 169 2368
rect 162 2358 169 2361
rect 182 2362 185 2368
rect 330 2358 598 2361
rect 610 2358 646 2361
rect 650 2358 766 2361
rect 826 2358 846 2361
rect 882 2358 894 2361
rect 962 2358 1102 2361
rect 1170 2358 1206 2361
rect 1234 2358 1710 2361
rect 1714 2358 1926 2361
rect 1962 2358 2046 2361
rect 2066 2358 2142 2361
rect 2190 2361 2193 2368
rect 2190 2358 2278 2361
rect 2346 2358 2382 2361
rect 2394 2358 2478 2361
rect 2482 2358 2489 2361
rect 2514 2358 2814 2361
rect 2938 2358 3166 2361
rect 3170 2358 3190 2361
rect 3202 2358 3230 2361
rect 3250 2358 3254 2361
rect 3266 2358 3310 2361
rect 3314 2358 3326 2361
rect 3338 2358 3358 2361
rect 3474 2358 3638 2361
rect 3754 2358 3766 2361
rect 3810 2358 3814 2361
rect 3870 2361 3873 2368
rect 3870 2358 3910 2361
rect 4002 2358 4025 2361
rect 4034 2358 4198 2361
rect 4218 2358 4342 2361
rect 4514 2358 4526 2361
rect 4538 2358 4542 2361
rect 4806 2361 4809 2368
rect 4786 2358 4809 2361
rect 4834 2358 4886 2361
rect 4906 2358 4942 2361
rect 4994 2358 5070 2361
rect 5094 2361 5097 2368
rect 5094 2358 5134 2361
rect 94 2352 97 2358
rect -26 2351 -22 2352
rect -26 2348 6 2351
rect 214 2351 217 2358
rect 1126 2352 1129 2358
rect 2822 2352 2825 2358
rect 4022 2352 4025 2358
rect 162 2348 217 2351
rect 354 2348 366 2351
rect 370 2348 526 2351
rect 530 2348 622 2351
rect 626 2348 646 2351
rect 650 2348 934 2351
rect 1018 2348 1110 2351
rect 1218 2348 1222 2351
rect 1302 2348 1326 2351
rect 1346 2348 1350 2351
rect 1358 2348 1446 2351
rect 1514 2348 1622 2351
rect 1650 2348 1670 2351
rect 1722 2348 1726 2351
rect 1754 2348 1790 2351
rect 1794 2348 1838 2351
rect 1890 2348 1934 2351
rect 1946 2348 1950 2351
rect 2018 2348 2070 2351
rect 2266 2348 2302 2351
rect 2322 2348 2326 2351
rect 2362 2348 2414 2351
rect 2458 2348 2518 2351
rect 2526 2348 2590 2351
rect 2594 2348 2614 2351
rect 2618 2348 2673 2351
rect 2746 2348 2777 2351
rect 2890 2348 2942 2351
rect 2962 2348 2974 2351
rect 3298 2348 3302 2351
rect 3362 2348 3382 2351
rect 3386 2348 3398 2351
rect 3418 2348 3494 2351
rect 3586 2348 3598 2351
rect 3602 2348 3630 2351
rect 3850 2348 3862 2351
rect 4042 2348 4054 2351
rect 4130 2348 4134 2351
rect 4186 2348 4190 2351
rect 4202 2348 4206 2351
rect 4210 2348 4238 2351
rect 4370 2348 4374 2351
rect 4478 2351 4481 2358
rect 4474 2348 4481 2351
rect 4770 2348 4798 2351
rect 4858 2348 4894 2351
rect 4898 2348 4902 2351
rect 5058 2348 5118 2351
rect 1302 2342 1305 2348
rect 474 2338 486 2341
rect 514 2338 526 2341
rect 586 2338 638 2341
rect 794 2338 814 2341
rect 874 2338 878 2341
rect 922 2338 934 2341
rect 1106 2338 1118 2341
rect 1154 2338 1238 2341
rect 1266 2338 1294 2341
rect 1358 2341 1361 2348
rect 1354 2338 1361 2341
rect 1394 2338 1486 2341
rect 1522 2338 1598 2341
rect 1634 2338 1798 2341
rect 1850 2338 2006 2341
rect 2010 2338 2038 2341
rect 2098 2338 2110 2341
rect 2174 2341 2177 2348
rect 2230 2341 2233 2348
rect 2138 2338 2177 2341
rect 2206 2338 2233 2341
rect 2314 2338 2318 2341
rect 2370 2338 2374 2341
rect 2442 2338 2494 2341
rect 2526 2341 2529 2348
rect 2670 2342 2673 2348
rect 2774 2342 2777 2348
rect 3174 2342 3177 2348
rect 2506 2338 2529 2341
rect 2578 2338 2582 2341
rect 2618 2338 2622 2341
rect 2882 2338 2886 2341
rect 2986 2338 3054 2341
rect 3234 2338 3249 2341
rect 3314 2338 3318 2341
rect 3370 2338 3502 2341
rect 3522 2338 3542 2341
rect 3730 2338 3822 2341
rect 3830 2341 3833 2348
rect 4926 2342 4929 2348
rect 5054 2342 5057 2348
rect 3826 2338 3833 2341
rect 3954 2338 3982 2341
rect 4034 2338 4049 2341
rect 4058 2338 4414 2341
rect 4466 2338 4598 2341
rect 4706 2338 4710 2341
rect 4734 2338 4750 2341
rect 4874 2338 4910 2341
rect 5058 2338 5086 2341
rect 5106 2338 5110 2341
rect 502 2332 505 2338
rect 2206 2332 2209 2338
rect -26 2331 -22 2332
rect -26 2328 6 2331
rect 770 2328 846 2331
rect 938 2328 1150 2331
rect 1162 2328 1382 2331
rect 1410 2328 1430 2331
rect 1578 2328 1638 2331
rect 1690 2328 1694 2331
rect 1842 2328 1870 2331
rect 1874 2328 1902 2331
rect 1922 2328 1974 2331
rect 2034 2328 2054 2331
rect 2082 2328 2094 2331
rect 2106 2328 2182 2331
rect 2186 2328 2198 2331
rect 2242 2328 2286 2331
rect 2290 2328 2297 2331
rect 2326 2328 2497 2331
rect 2506 2328 2534 2331
rect 2546 2328 2790 2331
rect 2826 2328 3030 2331
rect 3070 2331 3073 2338
rect 3246 2332 3249 2338
rect 4046 2332 4049 2338
rect 4734 2332 4737 2338
rect 5126 2332 5129 2338
rect 3070 2328 3134 2331
rect 3138 2328 3238 2331
rect 3366 2328 3374 2331
rect 3378 2328 3414 2331
rect 3458 2328 3526 2331
rect 3530 2328 3550 2331
rect 3610 2328 3646 2331
rect 3762 2328 3766 2331
rect 3842 2328 4022 2331
rect 4082 2328 4262 2331
rect 4306 2328 4398 2331
rect 4626 2328 4734 2331
rect 5050 2328 5086 2331
rect 306 2318 382 2321
rect 410 2318 662 2321
rect 802 2318 806 2321
rect 818 2318 1694 2321
rect 1822 2321 1825 2328
rect 1918 2322 1921 2328
rect 1698 2318 1825 2321
rect 1842 2318 1870 2321
rect 1898 2318 1910 2321
rect 1938 2318 1942 2321
rect 2010 2318 2022 2321
rect 2326 2321 2329 2328
rect 2194 2318 2329 2321
rect 2338 2318 2486 2321
rect 2494 2321 2497 2328
rect 3278 2322 3281 2328
rect 3422 2322 3425 2328
rect 2494 2318 2510 2321
rect 2818 2318 3054 2321
rect 3526 2318 4174 2321
rect 4202 2318 4222 2321
rect 4242 2318 4246 2321
rect 4250 2318 4310 2321
rect 4314 2318 4326 2321
rect 4362 2318 4366 2321
rect 4414 2321 4417 2328
rect 4386 2318 4417 2321
rect 4434 2318 4534 2321
rect 4642 2318 4646 2321
rect 4738 2318 4822 2321
rect 4946 2318 5030 2321
rect 5034 2318 5134 2321
rect 782 2312 785 2318
rect 3526 2312 3529 2318
rect 138 2308 510 2311
rect 802 2308 910 2311
rect 1170 2308 1174 2311
rect 1266 2308 1374 2311
rect 1434 2308 1494 2311
rect 1498 2308 1526 2311
rect 1594 2308 1598 2311
rect 1626 2308 1638 2311
rect 1658 2308 1662 2311
rect 1802 2308 1854 2311
rect 1890 2308 1926 2311
rect 1994 2308 2006 2311
rect 2170 2308 2286 2311
rect 2290 2308 2302 2311
rect 2306 2308 2358 2311
rect 2634 2308 2678 2311
rect 2762 2308 2782 2311
rect 2786 2308 2854 2311
rect 2866 2308 2910 2311
rect 2946 2308 3030 2311
rect 3050 2308 3070 2311
rect 3122 2308 3262 2311
rect 3266 2308 3318 2311
rect 3330 2308 3478 2311
rect 3502 2308 3526 2311
rect 3542 2308 3614 2311
rect 3626 2308 3702 2311
rect 3914 2308 3974 2311
rect 4194 2308 4238 2311
rect 4322 2308 4390 2311
rect 4426 2308 4694 2311
rect 4802 2308 5030 2311
rect 5034 2308 5070 2311
rect 1048 2303 1050 2307
rect 1054 2303 1057 2307
rect 1062 2303 1064 2307
rect 1878 2302 1881 2308
rect 2072 2303 2074 2307
rect 2078 2303 2081 2307
rect 2086 2303 2088 2307
rect 2134 2302 2137 2308
rect 3096 2303 3098 2307
rect 3102 2303 3105 2307
rect 3110 2303 3112 2307
rect 3502 2302 3505 2308
rect 3542 2302 3545 2308
rect 4112 2303 4114 2307
rect 4118 2303 4121 2307
rect 4126 2303 4128 2307
rect 362 2298 382 2301
rect 394 2298 446 2301
rect 450 2298 470 2301
rect 506 2298 550 2301
rect 554 2298 630 2301
rect 634 2298 710 2301
rect 714 2298 830 2301
rect 834 2298 854 2301
rect 906 2298 958 2301
rect 1234 2298 1350 2301
rect 1410 2298 1670 2301
rect 1738 2298 1758 2301
rect 1762 2298 1806 2301
rect 1850 2298 1854 2301
rect 1890 2298 1950 2301
rect 1954 2298 2065 2301
rect 2162 2298 2198 2301
rect 2210 2298 2382 2301
rect 2450 2298 2694 2301
rect 2754 2298 2814 2301
rect 2826 2298 3070 2301
rect 3154 2298 3206 2301
rect 3242 2298 3326 2301
rect 3330 2298 3334 2301
rect 3346 2298 3350 2301
rect 3386 2298 3398 2301
rect 3498 2298 3502 2301
rect 3530 2298 3542 2301
rect 3562 2298 3566 2301
rect 3578 2298 3630 2301
rect 3682 2298 3686 2301
rect 3818 2298 3878 2301
rect 3882 2298 3902 2301
rect 4002 2298 4078 2301
rect 4178 2298 4342 2301
rect 4346 2298 4366 2301
rect 4370 2298 4662 2301
rect 4666 2298 4790 2301
rect 5066 2298 5078 2301
rect 5098 2298 5110 2301
rect 18 2288 134 2291
rect 298 2288 326 2291
rect 330 2288 454 2291
rect 594 2288 630 2291
rect 986 2288 1494 2291
rect 1506 2288 1654 2291
rect 1746 2288 1881 2291
rect 1890 2288 1950 2291
rect 1954 2288 1998 2291
rect 2002 2288 2054 2291
rect 2062 2291 2065 2298
rect 2062 2288 2102 2291
rect 2106 2288 2270 2291
rect 2290 2288 2310 2291
rect 2386 2288 2718 2291
rect 2722 2288 2934 2291
rect 2962 2288 3758 2291
rect 3786 2288 3798 2291
rect 3810 2288 3830 2291
rect 3866 2288 3886 2291
rect 3890 2288 4158 2291
rect 4202 2288 4206 2291
rect 4290 2288 4334 2291
rect 4354 2288 4494 2291
rect 4538 2288 4574 2291
rect 5026 2288 5054 2291
rect 5082 2288 5102 2291
rect 5130 2288 5142 2291
rect 5146 2288 5150 2291
rect 74 2278 118 2281
rect 218 2278 350 2281
rect 478 2281 481 2288
rect 478 2278 582 2281
rect 618 2278 774 2281
rect 874 2278 1046 2281
rect 1050 2278 1105 2281
rect 1114 2278 1118 2281
rect 1202 2278 1254 2281
rect 1266 2278 1329 2281
rect 1338 2278 1342 2281
rect 1506 2278 1582 2281
rect 1698 2278 1750 2281
rect 1842 2278 1862 2281
rect 1878 2281 1881 2288
rect 1878 2278 1918 2281
rect 2002 2278 2014 2281
rect 2202 2278 2230 2281
rect 2266 2278 2326 2281
rect 2546 2278 2550 2281
rect 2570 2278 2702 2281
rect 2746 2278 2854 2281
rect 2914 2278 2958 2281
rect 3002 2278 3006 2281
rect 3014 2278 3062 2281
rect 3066 2278 3222 2281
rect 3234 2278 3238 2281
rect 3314 2278 3334 2281
rect 3338 2278 3574 2281
rect 3634 2278 3926 2281
rect 3930 2278 4598 2281
rect 4650 2278 4686 2281
rect 4834 2278 4838 2281
rect 4890 2278 4934 2281
rect 5010 2278 5086 2281
rect 5106 2278 5134 2281
rect 1102 2272 1105 2278
rect 114 2268 294 2271
rect 306 2268 342 2271
rect 474 2268 510 2271
rect 682 2268 790 2271
rect 794 2268 806 2271
rect 874 2268 894 2271
rect 1110 2268 1174 2271
rect 1250 2268 1286 2271
rect 1290 2268 1302 2271
rect 1326 2271 1329 2278
rect 1678 2272 1681 2278
rect 2238 2272 2241 2278
rect 3014 2272 3017 2278
rect 1326 2268 1478 2271
rect 1486 2268 1510 2271
rect 1538 2268 1542 2271
rect 1618 2268 1622 2271
rect 1666 2268 1670 2271
rect 1722 2268 1726 2271
rect 1794 2268 1942 2271
rect 1946 2268 1958 2271
rect 1970 2268 1998 2271
rect 2042 2268 2126 2271
rect 2154 2268 2174 2271
rect 2274 2268 2278 2271
rect 2306 2268 2374 2271
rect 2378 2268 2406 2271
rect 2426 2268 2654 2271
rect 2682 2268 2726 2271
rect 2778 2268 2806 2271
rect 2810 2268 2950 2271
rect 2970 2268 2974 2271
rect 3050 2268 3070 2271
rect 3194 2268 3302 2271
rect 3330 2268 3334 2271
rect 3378 2268 4374 2271
rect 4378 2268 4774 2271
rect 4778 2268 4926 2271
rect 4930 2268 4950 2271
rect 4954 2268 5110 2271
rect 5114 2268 5150 2271
rect 114 2258 126 2261
rect 170 2258 270 2261
rect 274 2258 350 2261
rect 354 2258 366 2261
rect 570 2258 590 2261
rect 618 2258 622 2261
rect 650 2258 654 2261
rect 730 2258 742 2261
rect 794 2258 814 2261
rect 918 2261 921 2268
rect 1110 2262 1113 2268
rect 1486 2262 1489 2268
rect 1750 2262 1753 2268
rect 866 2258 921 2261
rect 946 2258 950 2261
rect 1194 2258 1198 2261
rect 1218 2258 1222 2261
rect 1234 2258 1310 2261
rect 1314 2258 1374 2261
rect 1506 2258 1726 2261
rect 1730 2258 1734 2261
rect 1782 2261 1785 2268
rect 1782 2258 1886 2261
rect 1898 2258 2046 2261
rect 2066 2258 2142 2261
rect 2450 2258 2454 2261
rect 2538 2258 2694 2261
rect 2706 2258 2766 2261
rect 2922 2258 2990 2261
rect 2994 2258 3046 2261
rect 3094 2261 3097 2268
rect 3082 2258 3097 2261
rect 3106 2258 3313 2261
rect 3330 2258 3342 2261
rect 3354 2258 3406 2261
rect 3418 2258 3550 2261
rect 3554 2258 3590 2261
rect 3642 2258 3742 2261
rect 3754 2258 3838 2261
rect 3842 2258 4030 2261
rect 4034 2258 4102 2261
rect 4194 2258 4246 2261
rect 4298 2258 4358 2261
rect 4466 2258 4470 2261
rect 4482 2258 4510 2261
rect 4562 2258 4630 2261
rect 4698 2258 4702 2261
rect 4826 2258 4846 2261
rect 4858 2258 4886 2261
rect 4938 2258 5158 2261
rect 5162 2258 5190 2261
rect 234 2248 305 2251
rect 566 2251 569 2258
rect 2150 2252 2153 2258
rect 450 2248 569 2251
rect 574 2248 606 2251
rect 690 2248 718 2251
rect 894 2248 902 2251
rect 906 2248 982 2251
rect 1154 2248 1161 2251
rect 1282 2248 1406 2251
rect 1554 2248 1598 2251
rect 1674 2248 1710 2251
rect 1714 2248 1782 2251
rect 1818 2248 2014 2251
rect 2018 2248 2054 2251
rect 2066 2248 2070 2251
rect 2106 2248 2118 2251
rect 2214 2251 2217 2258
rect 2162 2248 2217 2251
rect 2234 2248 2318 2251
rect 2354 2248 2646 2251
rect 2650 2248 2750 2251
rect 2754 2248 2838 2251
rect 2842 2248 3102 2251
rect 3146 2248 3174 2251
rect 3310 2251 3313 2258
rect 4286 2252 4289 2258
rect 3266 2248 3305 2251
rect 3310 2248 3358 2251
rect 3402 2248 3494 2251
rect 3634 2248 3646 2251
rect 3714 2248 3758 2251
rect 3762 2248 3782 2251
rect 3822 2248 3846 2251
rect 3850 2248 3918 2251
rect 3978 2248 3982 2251
rect 4050 2248 4070 2251
rect 4074 2248 4118 2251
rect 4198 2248 4214 2251
rect 4330 2248 4430 2251
rect 4442 2248 4462 2251
rect 4698 2248 4702 2251
rect 4706 2248 4726 2251
rect 4754 2248 4966 2251
rect 5010 2248 5142 2251
rect 302 2242 305 2248
rect 574 2242 577 2248
rect 3302 2242 3305 2248
rect 3366 2242 3369 2248
rect 706 2238 846 2241
rect 850 2238 1081 2241
rect 1122 2238 1294 2241
rect 1306 2238 1334 2241
rect 1354 2238 1462 2241
rect 1466 2238 1606 2241
rect 1706 2238 1742 2241
rect 1754 2238 2094 2241
rect 2122 2238 2137 2241
rect 2170 2238 2254 2241
rect 2258 2238 2606 2241
rect 2886 2238 2942 2241
rect 2946 2238 3046 2241
rect 3090 2238 3158 2241
rect 3502 2241 3505 2248
rect 3806 2242 3809 2248
rect 3822 2242 3825 2248
rect 3466 2238 3505 2241
rect 3514 2238 3702 2241
rect 3730 2238 3737 2241
rect 3762 2238 3766 2241
rect 3898 2238 3902 2241
rect 4198 2241 4201 2248
rect 4066 2238 4201 2241
rect 4266 2238 4294 2241
rect 4462 2238 4582 2241
rect 4726 2241 4729 2248
rect 4726 2238 4790 2241
rect 4802 2238 4886 2241
rect 1078 2232 1081 2238
rect 2134 2232 2137 2238
rect 2846 2232 2849 2238
rect 2886 2232 2889 2238
rect 3734 2232 3737 2238
rect 3862 2232 3865 2238
rect 3870 2232 3873 2238
rect 202 2228 486 2231
rect 546 2228 622 2231
rect 682 2228 870 2231
rect 914 2228 958 2231
rect 1170 2228 1238 2231
rect 1298 2228 1662 2231
rect 1714 2228 2078 2231
rect 2210 2228 2302 2231
rect 2498 2228 2798 2231
rect 2962 2228 3006 2231
rect 3010 2228 3017 2231
rect 3066 2228 3102 2231
rect 3122 2228 3286 2231
rect 3298 2228 3326 2231
rect 3330 2228 3566 2231
rect 3570 2228 3721 2231
rect 3882 2228 3942 2231
rect 4214 2231 4217 2238
rect 4462 2232 4465 2238
rect 4214 2228 4230 2231
rect 4258 2228 4414 2231
rect 4506 2228 4614 2231
rect 4650 2228 4798 2231
rect 5034 2228 5134 2231
rect 678 2221 681 2228
rect 442 2218 681 2221
rect 834 2218 846 2221
rect 850 2218 886 2221
rect 890 2218 926 2221
rect 1210 2218 1214 2221
rect 1310 2218 1318 2221
rect 1322 2218 1638 2221
rect 1810 2218 1822 2221
rect 1834 2218 1838 2221
rect 1874 2218 1886 2221
rect 1930 2218 1934 2221
rect 1994 2218 2006 2221
rect 2018 2218 2049 2221
rect 2058 2218 2110 2221
rect 2122 2218 2142 2221
rect 2154 2218 2350 2221
rect 2362 2218 2534 2221
rect 2594 2218 2654 2221
rect 2746 2218 2790 2221
rect 2794 2218 2902 2221
rect 3018 2218 3126 2221
rect 3138 2218 3470 2221
rect 3718 2221 3721 2228
rect 3718 2218 3766 2221
rect 3810 2218 4390 2221
rect 4602 2218 4974 2221
rect 298 2208 446 2211
rect 698 2208 1542 2211
rect 1690 2208 1718 2211
rect 1870 2211 1873 2218
rect 1966 2212 1969 2218
rect 1746 2208 1873 2211
rect 1914 2208 1934 2211
rect 2046 2211 2049 2218
rect 2046 2208 2230 2211
rect 2234 2208 2486 2211
rect 2506 2208 2518 2211
rect 2610 2208 3126 2211
rect 3162 2208 3446 2211
rect 3450 2208 3462 2211
rect 3474 2208 3534 2211
rect 3578 2208 3582 2211
rect 3890 2208 4134 2211
rect 4138 2208 4174 2211
rect 4210 2208 4422 2211
rect 4730 2208 4766 2211
rect 4842 2208 5182 2211
rect 536 2203 538 2207
rect 542 2203 545 2207
rect 550 2203 552 2207
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1574 2203 1576 2207
rect 1950 2202 1953 2208
rect 2584 2203 2586 2207
rect 2590 2203 2593 2207
rect 2598 2203 2600 2207
rect 3608 2203 3610 2207
rect 3614 2203 3617 2207
rect 3622 2203 3624 2207
rect 4632 2203 4634 2207
rect 4638 2203 4641 2207
rect 4646 2203 4648 2207
rect 602 2198 814 2201
rect 834 2198 918 2201
rect 1250 2198 1422 2201
rect 1442 2198 1526 2201
rect 1586 2198 1814 2201
rect 1866 2198 1878 2201
rect 1922 2198 1926 2201
rect 1994 2198 2070 2201
rect 2074 2198 2102 2201
rect 2210 2198 2486 2201
rect 2794 2198 3310 2201
rect 3330 2198 3414 2201
rect 3474 2198 3478 2201
rect 3778 2198 4030 2201
rect 4042 2198 4278 2201
rect 4298 2198 4350 2201
rect 4690 2198 4830 2201
rect 154 2188 366 2191
rect 426 2188 582 2191
rect 682 2188 838 2191
rect 866 2188 870 2191
rect 938 2188 1169 2191
rect 1178 2188 1246 2191
rect 1354 2188 1958 2191
rect 1994 2188 2062 2191
rect 2066 2188 2070 2191
rect 2082 2188 2185 2191
rect 2274 2188 2478 2191
rect 2482 2188 2510 2191
rect 2514 2188 2582 2191
rect 3050 2188 3214 2191
rect 3226 2188 3393 2191
rect 3514 2188 3654 2191
rect 3674 2188 3745 2191
rect 3826 2188 3838 2191
rect 3930 2188 4022 2191
rect 4082 2188 4334 2191
rect 4730 2188 4774 2191
rect 4778 2188 4830 2191
rect 162 2178 278 2181
rect 282 2178 462 2181
rect 466 2178 702 2181
rect 722 2178 814 2181
rect 918 2181 921 2188
rect 818 2178 982 2181
rect 986 2178 1118 2181
rect 1138 2178 1150 2181
rect 1166 2181 1169 2188
rect 2182 2182 2185 2188
rect 1166 2178 1286 2181
rect 1370 2178 1814 2181
rect 1842 2178 1910 2181
rect 1938 2178 1958 2181
rect 1962 2178 2014 2181
rect 2034 2178 2046 2181
rect 2058 2178 2158 2181
rect 2234 2178 2430 2181
rect 2590 2181 2593 2188
rect 2450 2178 2758 2181
rect 2970 2178 3382 2181
rect 3390 2181 3393 2188
rect 3742 2182 3745 2188
rect 3390 2178 3633 2181
rect 3730 2178 3734 2181
rect 3778 2178 4694 2181
rect 4746 2178 5158 2181
rect 3630 2172 3633 2178
rect 226 2168 246 2171
rect 250 2168 382 2171
rect 482 2168 614 2171
rect 650 2168 1350 2171
rect 1362 2168 1398 2171
rect 1418 2168 1430 2171
rect 1458 2168 1598 2171
rect 1602 2168 1630 2171
rect 1698 2168 1726 2171
rect 1738 2168 1790 2171
rect 1938 2168 1990 2171
rect 2050 2168 2118 2171
rect 2202 2168 2286 2171
rect 2298 2168 2342 2171
rect 2466 2168 2470 2171
rect 2530 2168 2734 2171
rect 2810 2168 2926 2171
rect 2994 2168 2998 2171
rect 3018 2168 3030 2171
rect 3082 2168 3398 2171
rect 3442 2168 3582 2171
rect 3698 2168 3806 2171
rect 3810 2168 3822 2171
rect 3826 2168 4054 2171
rect 4154 2168 4246 2171
rect 4250 2168 4286 2171
rect 4290 2168 4318 2171
rect 4342 2168 4438 2171
rect 4490 2168 4550 2171
rect 4554 2168 4734 2171
rect 4738 2168 4758 2171
rect 4858 2168 5014 2171
rect 510 2162 513 2168
rect 1662 2162 1665 2168
rect 114 2158 230 2161
rect 234 2158 438 2161
rect 802 2158 846 2161
rect 858 2158 942 2161
rect 962 2158 1086 2161
rect 1090 2158 1118 2161
rect 1130 2158 1134 2161
rect 1394 2158 1398 2161
rect 1418 2158 1430 2161
rect 1434 2158 1542 2161
rect 1778 2158 1790 2161
rect 1902 2161 1905 2168
rect 1866 2158 1905 2161
rect 1922 2158 1958 2161
rect 2026 2158 2062 2161
rect 2146 2158 2150 2161
rect 2178 2158 2182 2161
rect 2202 2158 2302 2161
rect 2306 2158 2350 2161
rect 2378 2158 2446 2161
rect 2474 2158 2526 2161
rect 2622 2158 2774 2161
rect 2842 2158 2894 2161
rect 3006 2161 3009 2168
rect 2986 2158 3009 2161
rect 3042 2158 3054 2161
rect 3114 2158 3246 2161
rect 3266 2158 3270 2161
rect 3274 2158 3342 2161
rect 3514 2158 3558 2161
rect 3570 2158 3590 2161
rect 3594 2158 3630 2161
rect 3658 2158 3758 2161
rect 3770 2158 3782 2161
rect 3834 2158 3902 2161
rect 3922 2158 3974 2161
rect 4150 2158 4158 2161
rect 4162 2158 4190 2161
rect 4342 2161 4345 2168
rect 4258 2158 4345 2161
rect 4450 2158 4494 2161
rect 4530 2158 4742 2161
rect 4794 2158 4798 2161
rect 4858 2158 4862 2161
rect 4906 2158 4918 2161
rect 606 2152 609 2158
rect 630 2152 633 2158
rect 646 2152 649 2158
rect -26 2151 -22 2152
rect -26 2148 6 2151
rect 90 2148 94 2151
rect 170 2148 246 2151
rect 290 2148 313 2151
rect 410 2148 502 2151
rect 690 2148 694 2151
rect 702 2151 705 2158
rect 702 2148 710 2151
rect 754 2148 825 2151
rect 914 2148 958 2151
rect 974 2148 1025 2151
rect 1182 2151 1185 2158
rect 1130 2148 1185 2151
rect 1278 2151 1281 2158
rect 1318 2152 1321 2158
rect 1366 2152 1369 2158
rect 1990 2152 1993 2158
rect 1278 2148 1286 2151
rect 1370 2148 1406 2151
rect 1458 2148 1502 2151
rect 1506 2148 1526 2151
rect 1722 2148 1974 2151
rect 2066 2148 2078 2151
rect 2090 2148 2174 2151
rect 2178 2148 2182 2151
rect 2206 2148 2270 2151
rect 2282 2148 2286 2151
rect 2350 2151 2353 2158
rect 2290 2148 2305 2151
rect 2350 2148 2414 2151
rect 2438 2148 2502 2151
rect 2622 2151 2625 2158
rect 2546 2148 2625 2151
rect 2634 2148 2646 2151
rect 2794 2148 2894 2151
rect 2914 2148 2926 2151
rect 2954 2148 3078 2151
rect 3114 2148 3118 2151
rect 3274 2148 3310 2151
rect 3354 2148 3358 2151
rect 3410 2148 3422 2151
rect 3478 2151 3481 2158
rect 3478 2148 3494 2151
rect 3538 2148 3598 2151
rect 3602 2148 3606 2151
rect 3646 2151 3649 2158
rect 3646 2148 3678 2151
rect 3690 2148 3694 2151
rect 3746 2148 3750 2151
rect 3794 2148 3862 2151
rect 3866 2148 3894 2151
rect 3898 2148 3990 2151
rect 4026 2148 4030 2151
rect 4110 2151 4113 2158
rect 4222 2152 4225 2158
rect 4082 2148 4113 2151
rect 4154 2148 4182 2151
rect 4354 2148 4358 2151
rect 4490 2148 4518 2151
rect 4674 2148 4726 2151
rect 4750 2148 4790 2151
rect 4802 2148 4822 2151
rect 4826 2148 4934 2151
rect 4970 2148 5078 2151
rect 310 2142 313 2148
rect 822 2142 825 2148
rect 974 2142 977 2148
rect 1022 2142 1025 2148
rect 2206 2142 2209 2148
rect 2302 2142 2305 2148
rect 2438 2142 2441 2148
rect 186 2138 297 2141
rect 338 2138 494 2141
rect 570 2138 662 2141
rect 882 2138 894 2141
rect 906 2138 910 2141
rect 938 2138 942 2141
rect 1138 2138 1294 2141
rect 1370 2138 1382 2141
rect 1410 2138 1446 2141
rect 1522 2138 1622 2141
rect 1666 2138 1710 2141
rect 1802 2138 1830 2141
rect 1850 2138 1918 2141
rect 1938 2138 1942 2141
rect 1954 2138 1966 2141
rect 2002 2138 2054 2141
rect 2106 2138 2110 2141
rect 2126 2138 2142 2141
rect 2450 2138 2486 2141
rect 2890 2138 2926 2141
rect 2942 2141 2945 2148
rect 2942 2138 3038 2141
rect 3050 2138 3350 2141
rect 3418 2138 3446 2141
rect 3530 2138 3622 2141
rect 3642 2138 3654 2141
rect 3738 2138 3758 2141
rect 3858 2138 3862 2141
rect 3946 2138 4017 2141
rect 4042 2138 4142 2141
rect 4170 2138 4174 2141
rect 4306 2138 4366 2141
rect 4462 2141 4465 2148
rect 4750 2142 4753 2148
rect 4462 2138 4590 2141
rect 4650 2138 4654 2141
rect 4770 2138 4790 2141
rect 4794 2138 4846 2141
rect 4858 2138 4966 2141
rect 294 2132 297 2138
rect 370 2128 590 2131
rect 642 2128 646 2131
rect 650 2128 782 2131
rect 826 2128 830 2131
rect 934 2131 937 2138
rect 1126 2132 1129 2138
rect 1742 2132 1745 2138
rect 2126 2132 2129 2138
rect 866 2128 937 2131
rect 978 2128 990 2131
rect 1274 2128 1718 2131
rect 1786 2128 1814 2131
rect 1818 2128 1926 2131
rect 1946 2128 1958 2131
rect 1962 2128 1969 2131
rect 1978 2128 2014 2131
rect 2098 2128 2102 2131
rect 2530 2128 2534 2131
rect 2838 2131 2841 2138
rect 4014 2132 4017 2138
rect 2838 2128 2862 2131
rect 2954 2128 2974 2131
rect 3082 2128 3118 2131
rect 3170 2128 3302 2131
rect 3414 2128 3550 2131
rect 3554 2128 3574 2131
rect 3650 2128 3774 2131
rect 3858 2128 3958 2131
rect 4042 2128 4046 2131
rect 4170 2128 4230 2131
rect 4370 2128 4374 2131
rect 4414 2131 4417 2138
rect 4414 2128 4502 2131
rect 4530 2128 4534 2131
rect 4570 2128 4718 2131
rect 4794 2128 4862 2131
rect 4954 2128 4998 2131
rect 5074 2128 5134 2131
rect 2670 2122 2673 2128
rect 3054 2122 3057 2128
rect 3134 2122 3137 2128
rect 122 2118 286 2121
rect 298 2118 526 2121
rect 562 2118 566 2121
rect 762 2118 766 2121
rect 818 2118 870 2121
rect 982 2118 1302 2121
rect 1330 2118 1470 2121
rect 1490 2118 1550 2121
rect 1562 2118 1702 2121
rect 1730 2118 1790 2121
rect 1794 2118 1809 2121
rect 1818 2118 1878 2121
rect 1882 2118 1886 2121
rect 1914 2118 2062 2121
rect 2146 2118 2294 2121
rect 2882 2118 2982 2121
rect 2986 2118 3014 2121
rect 3082 2118 3134 2121
rect 3226 2118 3270 2121
rect 3278 2118 3302 2121
rect 3414 2121 3417 2128
rect 4950 2122 4953 2128
rect 3322 2118 3417 2121
rect 3426 2118 3558 2121
rect 3586 2118 3822 2121
rect 3962 2118 4006 2121
rect 4114 2118 4382 2121
rect 4706 2118 4718 2121
rect 5058 2118 5150 2121
rect 982 2112 985 2118
rect 218 2108 222 2111
rect 234 2108 246 2111
rect 450 2108 478 2111
rect 490 2108 502 2111
rect 506 2108 694 2111
rect 698 2108 806 2111
rect 810 2108 886 2111
rect 890 2108 982 2111
rect 1098 2108 1126 2111
rect 1178 2108 1334 2111
rect 1338 2108 1398 2111
rect 1634 2108 1662 2111
rect 1674 2108 1678 2111
rect 1706 2108 1798 2111
rect 1806 2111 1809 2118
rect 3278 2112 3281 2118
rect 1806 2108 1894 2111
rect 1930 2108 1990 2111
rect 2114 2108 2254 2111
rect 2506 2108 2534 2111
rect 2538 2108 2590 2111
rect 2594 2108 2734 2111
rect 2938 2108 2990 2111
rect 2998 2108 3006 2111
rect 3130 2108 3142 2111
rect 3146 2108 3150 2111
rect 3194 2108 3198 2111
rect 3290 2108 3326 2111
rect 3466 2108 3486 2111
rect 3506 2108 3526 2111
rect 3706 2108 3710 2111
rect 3818 2108 3886 2111
rect 4346 2108 4518 2111
rect 4994 2108 5022 2111
rect 1048 2103 1050 2107
rect 1054 2103 1057 2107
rect 1062 2103 1064 2107
rect 2072 2103 2074 2107
rect 2078 2103 2081 2107
rect 2086 2103 2088 2107
rect 170 2098 302 2101
rect 650 2098 718 2101
rect 722 2098 886 2101
rect 890 2098 1006 2101
rect 1082 2098 1345 2101
rect 1354 2098 1374 2101
rect 1378 2098 1494 2101
rect 1498 2098 1574 2101
rect 1578 2098 1758 2101
rect 1770 2098 1846 2101
rect 1874 2098 1902 2101
rect 1906 2098 1934 2101
rect 1946 2098 2046 2101
rect 2186 2098 2246 2101
rect 2266 2098 2278 2101
rect 2310 2101 2313 2108
rect 2998 2102 3001 2108
rect 3096 2103 3098 2107
rect 3102 2103 3105 2107
rect 3110 2103 3112 2107
rect 4112 2103 4114 2107
rect 4118 2103 4121 2107
rect 4126 2103 4128 2107
rect 2282 2098 2313 2101
rect 2322 2098 2921 2101
rect 3178 2098 3646 2101
rect 3914 2098 3966 2101
rect 4178 2098 4262 2101
rect 4346 2098 4358 2101
rect 4434 2098 4494 2101
rect 4938 2098 5062 2101
rect 5170 2098 5174 2101
rect 18 2088 70 2091
rect 218 2088 222 2091
rect 230 2088 238 2091
rect 242 2088 774 2091
rect 854 2088 974 2091
rect 1006 2091 1009 2098
rect 1006 2088 1166 2091
rect 1222 2088 1230 2091
rect 1234 2088 1238 2091
rect 1250 2088 1270 2091
rect 1342 2091 1345 2098
rect 1342 2088 1465 2091
rect 1474 2088 1518 2091
rect 1522 2088 1598 2091
rect 1602 2088 1678 2091
rect 1682 2088 1718 2091
rect 1874 2088 1894 2091
rect 1930 2088 2038 2091
rect 2042 2088 2318 2091
rect 2394 2088 2398 2091
rect 2426 2088 2542 2091
rect 2710 2088 2766 2091
rect 2770 2088 2822 2091
rect 2918 2091 2921 2098
rect 3174 2091 3177 2098
rect 2918 2088 3177 2091
rect 3298 2088 3366 2091
rect 3370 2088 3382 2091
rect 3418 2088 3534 2091
rect 3554 2088 4390 2091
rect 4394 2088 4414 2091
rect 4458 2088 4710 2091
rect 4738 2088 4878 2091
rect 4906 2088 5121 2091
rect 158 2081 161 2088
rect 854 2082 857 2088
rect 1190 2082 1193 2088
rect 1462 2082 1465 2088
rect 2710 2082 2713 2088
rect 74 2078 161 2081
rect 170 2078 190 2081
rect 194 2078 230 2081
rect 330 2078 486 2081
rect 490 2078 518 2081
rect 538 2078 582 2081
rect 626 2078 702 2081
rect 746 2078 838 2081
rect 1042 2078 1094 2081
rect 1098 2078 1102 2081
rect 1154 2078 1166 2081
rect 1218 2078 1310 2081
rect 1458 2078 1462 2081
rect 1554 2078 1625 2081
rect 1630 2078 1638 2081
rect 1730 2078 1790 2081
rect 1794 2078 1910 2081
rect 1930 2078 2110 2081
rect 2162 2078 2233 2081
rect 2258 2078 2342 2081
rect 2362 2078 2430 2081
rect 2434 2078 2510 2081
rect 2514 2078 2550 2081
rect 2738 2078 2790 2081
rect 2794 2078 2934 2081
rect 3026 2078 3126 2081
rect 3254 2081 3257 2088
rect 5118 2082 5121 2088
rect 5174 2082 5177 2088
rect 3146 2078 3462 2081
rect 3506 2078 3686 2081
rect 3786 2078 3870 2081
rect 3906 2078 3910 2081
rect 3946 2078 4086 2081
rect 4090 2078 4110 2081
rect 4122 2078 4134 2081
rect 4170 2078 4254 2081
rect 4386 2078 4438 2081
rect 4474 2078 4478 2081
rect 4626 2078 4814 2081
rect 4922 2078 4982 2081
rect 4986 2078 5030 2081
rect 122 2068 134 2071
rect 178 2068 438 2071
rect 442 2068 686 2071
rect 762 2068 1030 2071
rect 1034 2068 1230 2071
rect 1310 2071 1313 2078
rect 1306 2068 1313 2071
rect 1342 2072 1345 2078
rect 1502 2072 1505 2078
rect 1586 2068 1590 2071
rect 1598 2068 1614 2071
rect 1622 2071 1625 2078
rect 1926 2071 1929 2078
rect 2118 2072 2121 2078
rect 2230 2072 2233 2078
rect 2350 2072 2353 2078
rect 5094 2072 5097 2078
rect 5110 2072 5113 2078
rect 1622 2068 1929 2071
rect 1978 2068 2006 2071
rect 2058 2068 2102 2071
rect 2154 2068 2222 2071
rect 2282 2068 2310 2071
rect 2314 2068 2318 2071
rect 2378 2068 2462 2071
rect 2586 2068 2622 2071
rect 2794 2068 2830 2071
rect 2834 2068 2894 2071
rect 3122 2068 3182 2071
rect 3402 2068 3414 2071
rect 3442 2068 3446 2071
rect 3490 2068 3518 2071
rect 3674 2068 3718 2071
rect 3722 2068 3729 2071
rect 3850 2068 3862 2071
rect 3930 2068 3942 2071
rect 3946 2068 4046 2071
rect 4066 2068 4070 2071
rect 4114 2068 4198 2071
rect 4202 2068 4486 2071
rect 4490 2068 4526 2071
rect 4570 2068 4582 2071
rect 4666 2068 4742 2071
rect 4746 2068 4774 2071
rect 4978 2068 4990 2071
rect 5010 2068 5014 2071
rect 5066 2068 5070 2071
rect 5154 2068 5182 2071
rect 134 2062 137 2068
rect 138 2058 422 2061
rect 442 2058 446 2061
rect 578 2058 750 2061
rect 810 2058 982 2061
rect 994 2058 998 2061
rect 1002 2058 1110 2061
rect 1122 2058 1126 2061
rect 1154 2058 1174 2061
rect 1274 2058 1286 2061
rect 1294 2061 1297 2068
rect 1294 2059 1390 2061
rect 1486 2062 1489 2068
rect 1294 2058 1393 2059
rect 1598 2061 1601 2068
rect 2710 2062 2713 2068
rect 1570 2058 1601 2061
rect 1606 2058 1614 2061
rect 1690 2058 1694 2061
rect 1738 2058 1758 2061
rect 1834 2058 1878 2061
rect 1898 2058 2614 2061
rect 2738 2058 2766 2061
rect 2770 2058 2814 2061
rect 2818 2058 2862 2061
rect 2930 2058 2934 2061
rect 3070 2061 3073 2068
rect 3042 2058 3073 2061
rect 3098 2058 3142 2061
rect 3206 2061 3209 2068
rect 3398 2062 3401 2068
rect 4798 2062 4801 2068
rect 5038 2062 5041 2068
rect 3206 2058 3334 2061
rect 3434 2058 3446 2061
rect 3474 2058 3478 2061
rect 3522 2058 3654 2061
rect 3730 2058 3910 2061
rect 3938 2058 4014 2061
rect 4130 2058 4238 2061
rect 4314 2058 4401 2061
rect 4410 2058 4438 2061
rect 4482 2058 4590 2061
rect 4594 2058 4782 2061
rect 5050 2058 5062 2061
rect 5090 2058 5110 2061
rect 5222 2061 5226 2062
rect 5194 2058 5226 2061
rect 1606 2052 1609 2058
rect 3174 2052 3177 2058
rect 106 2048 182 2051
rect 370 2048 374 2051
rect 466 2048 473 2051
rect 490 2048 510 2051
rect 578 2048 598 2051
rect 682 2048 718 2051
rect 722 2048 742 2051
rect 770 2048 790 2051
rect 938 2048 974 2051
rect 1026 2048 1238 2051
rect 1274 2048 1446 2051
rect 1450 2048 1526 2051
rect 1706 2048 1742 2051
rect 1834 2048 1838 2051
rect 1846 2048 1854 2051
rect 1858 2048 2078 2051
rect 2090 2048 2270 2051
rect 2378 2048 2449 2051
rect 2490 2048 2662 2051
rect 2706 2048 2830 2051
rect 2842 2048 2862 2051
rect 2870 2048 2878 2051
rect 2882 2048 2910 2051
rect 3034 2048 3118 2051
rect 3266 2048 3278 2051
rect 3298 2048 3462 2051
rect 3490 2048 3502 2051
rect 3506 2048 3542 2051
rect 3586 2048 3646 2051
rect 4082 2048 4382 2051
rect 4386 2048 4390 2051
rect 4398 2051 4401 2058
rect 4398 2048 4406 2051
rect 4466 2048 4574 2051
rect 4578 2048 4606 2051
rect 4662 2048 4702 2051
rect 4806 2048 4814 2051
rect 4818 2048 4894 2051
rect 4954 2048 5070 2051
rect 5074 2048 5166 2051
rect 5170 2048 5174 2051
rect 206 2041 209 2048
rect 162 2038 209 2041
rect 438 2041 441 2048
rect 274 2038 441 2041
rect 470 2042 473 2048
rect 530 2038 670 2041
rect 690 2038 958 2041
rect 1006 2041 1009 2048
rect 978 2038 1038 2041
rect 1058 2038 1078 2041
rect 1098 2038 1102 2041
rect 1114 2038 1166 2041
rect 1194 2038 1206 2041
rect 1282 2038 1310 2041
rect 1322 2038 1366 2041
rect 1546 2038 1630 2041
rect 1674 2038 1726 2041
rect 1762 2038 2174 2041
rect 2250 2038 2438 2041
rect 2446 2041 2449 2048
rect 2446 2038 2606 2041
rect 2730 2038 2734 2041
rect 2754 2038 2854 2041
rect 3018 2038 3318 2041
rect 3354 2038 3414 2041
rect 3426 2038 3446 2041
rect 3482 2038 3854 2041
rect 3986 2038 4110 2041
rect 4446 2041 4449 2048
rect 4662 2042 4665 2048
rect 4122 2038 4449 2041
rect 4498 2038 4518 2041
rect 4942 2041 4945 2048
rect 4942 2038 5150 2041
rect 5170 2038 5182 2041
rect 458 2028 494 2031
rect 818 2028 902 2031
rect 914 2028 985 2031
rect 1042 2028 1070 2031
rect 1186 2028 1190 2031
rect 1210 2028 1230 2031
rect 1274 2028 1774 2031
rect 1810 2028 2030 2031
rect 2106 2028 2406 2031
rect 2490 2028 3198 2031
rect 3434 2028 3494 2031
rect 3498 2028 3678 2031
rect 3682 2028 3998 2031
rect 4010 2028 4190 2031
rect 4194 2028 4206 2031
rect 4242 2028 4390 2031
rect 4418 2028 4638 2031
rect 4642 2028 4662 2031
rect 4666 2028 4670 2031
rect 4682 2028 4950 2031
rect 982 2022 985 2028
rect 5086 2022 5089 2028
rect 658 2018 734 2021
rect 738 2018 830 2021
rect 834 2018 846 2021
rect 1034 2018 1094 2021
rect 1274 2018 1334 2021
rect 1342 2018 1350 2021
rect 1354 2018 1670 2021
rect 1690 2018 1862 2021
rect 1914 2018 1974 2021
rect 1978 2018 2038 2021
rect 2042 2018 2158 2021
rect 2186 2018 2310 2021
rect 2362 2018 2382 2021
rect 2402 2018 2822 2021
rect 2866 2018 3286 2021
rect 3290 2018 3558 2021
rect 3562 2018 3766 2021
rect 3770 2018 3798 2021
rect 3810 2018 4062 2021
rect 4066 2018 4086 2021
rect 4170 2018 4934 2021
rect 4954 2018 5006 2021
rect 1110 2012 1113 2018
rect 4134 2012 4137 2018
rect 5102 2012 5105 2018
rect 90 2008 134 2011
rect 138 2008 262 2011
rect 266 2008 342 2011
rect 346 2008 518 2011
rect 666 2008 758 2011
rect 842 2008 966 2011
rect 994 2008 1054 2011
rect 1186 2008 1550 2011
rect 1650 2008 1790 2011
rect 1802 2008 2022 2011
rect 2122 2008 2134 2011
rect 2146 2008 2334 2011
rect 2338 2008 2494 2011
rect 2546 2008 2550 2011
rect 2658 2008 2758 2011
rect 2786 2008 2790 2011
rect 2834 2008 3038 2011
rect 3066 2008 3102 2011
rect 3346 2008 3478 2011
rect 3482 2008 3598 2011
rect 3658 2008 4078 2011
rect 4090 2008 4094 2011
rect 4218 2008 4406 2011
rect 4426 2008 4478 2011
rect 536 2003 538 2007
rect 542 2003 545 2007
rect 550 2003 552 2007
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1574 2003 1576 2007
rect 2584 2003 2586 2007
rect 2590 2003 2593 2007
rect 2598 2003 2600 2007
rect 3608 2003 3610 2007
rect 3614 2003 3617 2007
rect 3622 2003 3624 2007
rect 4632 2003 4634 2007
rect 4638 2003 4641 2007
rect 4646 2003 4648 2007
rect 5022 2002 5025 2008
rect 826 1998 998 2001
rect 1018 1998 1118 2001
rect 1418 1998 1510 2001
rect 1682 1998 1758 2001
rect 1786 1998 1950 2001
rect 1970 1998 1974 2001
rect 2018 1998 2110 2001
rect 2162 1998 2230 2001
rect 2234 1998 2286 2001
rect 2314 1998 2390 2001
rect 2394 1998 2574 2001
rect 2626 1998 2646 2001
rect 2650 1998 3454 2001
rect 3466 1998 3582 2001
rect 4026 1998 4134 2001
rect 4138 1998 4158 2001
rect 4306 1998 4454 2001
rect 4506 1998 4534 2001
rect 4538 1998 4542 2001
rect 1990 1992 1993 1998
rect 2118 1992 2121 1998
rect 570 1988 1342 1991
rect 1382 1988 1606 1991
rect 1714 1988 1750 1991
rect 2214 1988 2262 1991
rect 2298 1988 2406 1991
rect 2434 1988 2462 1991
rect 2466 1988 2662 1991
rect 2666 1988 2694 1991
rect 2802 1988 2998 1991
rect 3050 1988 3846 1991
rect 3850 1988 4030 1991
rect 4034 1988 4326 1991
rect 4330 1988 4374 1991
rect 4378 1988 4566 1991
rect 4570 1988 5046 1991
rect 5050 1988 5126 1991
rect 5130 1988 5150 1991
rect 254 1981 257 1988
rect 1382 1982 1385 1988
rect 186 1978 257 1981
rect 282 1978 302 1981
rect 638 1978 1334 1981
rect 1506 1978 1550 1981
rect 1554 1978 1742 1981
rect 1778 1978 1894 1981
rect 1906 1978 2006 1981
rect 2014 1981 2017 1988
rect 2214 1982 2217 1988
rect 2014 1978 2054 1981
rect 2242 1978 2246 1981
rect 2282 1978 2622 1981
rect 2650 1978 2870 1981
rect 2882 1978 3030 1981
rect 3054 1978 3086 1981
rect 3170 1978 3486 1981
rect 3594 1978 3710 1981
rect 3714 1978 3774 1981
rect 3794 1978 3982 1981
rect 4106 1978 4286 1981
rect 4586 1978 4894 1981
rect 5178 1978 5182 1981
rect 238 1968 281 1971
rect 638 1971 641 1978
rect 610 1968 641 1971
rect 706 1968 801 1971
rect 238 1962 241 1968
rect 278 1962 281 1968
rect 638 1962 641 1968
rect 798 1962 801 1968
rect 898 1968 1502 1971
rect 1538 1968 1542 1971
rect 1554 1968 1910 1971
rect 1922 1968 2006 1971
rect 2066 1968 2502 1971
rect 2538 1968 2622 1971
rect 2634 1968 2638 1971
rect 2642 1968 2718 1971
rect 2818 1968 2961 1971
rect 2986 1968 2998 1971
rect 3054 1971 3057 1978
rect 3018 1968 3057 1971
rect 3158 1971 3161 1978
rect 3158 1968 3198 1971
rect 3358 1968 3862 1971
rect 3866 1968 3918 1971
rect 3922 1968 4166 1971
rect 4186 1968 4254 1971
rect 4258 1968 4318 1971
rect 4470 1971 4473 1978
rect 4458 1968 4473 1971
rect 4498 1968 4590 1971
rect 4738 1968 4790 1971
rect 5022 1971 5025 1978
rect 4826 1968 5025 1971
rect 5090 1968 5190 1971
rect 878 1962 881 1968
rect 2958 1962 2961 1968
rect 3222 1962 3225 1968
rect 3358 1962 3361 1968
rect 282 1958 294 1961
rect 306 1958 462 1961
rect 466 1958 470 1961
rect 546 1958 622 1961
rect 714 1958 758 1961
rect 762 1958 790 1961
rect 890 1958 894 1961
rect 918 1958 926 1961
rect 930 1958 942 1961
rect 954 1958 966 1961
rect 1018 1958 1102 1961
rect 1154 1958 1158 1961
rect 1298 1958 1302 1961
rect 1354 1958 1358 1961
rect 1434 1958 1454 1961
rect 1842 1958 1862 1961
rect 1866 1958 1902 1961
rect 2210 1958 2478 1961
rect 2498 1958 2502 1961
rect 2546 1958 2558 1961
rect 2674 1958 2761 1961
rect 2778 1958 2870 1961
rect 2962 1958 2990 1961
rect 2994 1958 3142 1961
rect 3330 1958 3358 1961
rect 3458 1958 3462 1961
rect 3514 1958 3574 1961
rect 3626 1958 3718 1961
rect 3762 1958 3766 1961
rect 3794 1958 3822 1961
rect 3906 1958 3950 1961
rect 4002 1958 4038 1961
rect 4042 1958 4078 1961
rect 4114 1958 4150 1961
rect 4194 1958 4222 1961
rect 4238 1958 4246 1961
rect 4250 1958 4350 1961
rect 4458 1958 4470 1961
rect 4602 1958 4646 1961
rect 4650 1958 4657 1961
rect 4754 1958 4774 1961
rect 4778 1958 4854 1961
rect 4870 1958 4878 1961
rect 4882 1958 4958 1961
rect 5082 1958 5166 1961
rect 122 1948 246 1951
rect 426 1948 446 1951
rect 482 1948 486 1951
rect 506 1948 614 1951
rect 626 1948 694 1951
rect 794 1948 822 1951
rect 826 1948 966 1951
rect 970 1948 974 1951
rect 986 1948 1030 1951
rect 1050 1948 1070 1951
rect 1090 1948 1094 1951
rect 1146 1948 1206 1951
rect 1286 1951 1289 1958
rect 1310 1952 1313 1958
rect 1286 1948 1302 1951
rect 1338 1948 1382 1951
rect 1458 1948 1558 1951
rect 1594 1948 1662 1951
rect 1686 1951 1689 1958
rect 1734 1951 1737 1958
rect 1686 1948 1737 1951
rect 1778 1948 1785 1951
rect 1950 1951 1953 1958
rect 1898 1948 1953 1951
rect 2022 1952 2025 1958
rect 2494 1952 2497 1958
rect 2758 1952 2761 1958
rect 3430 1952 3433 1958
rect 3854 1952 3857 1958
rect 4494 1952 4497 1958
rect 2026 1948 2062 1951
rect 2082 1948 2086 1951
rect 2242 1948 2310 1951
rect 774 1942 777 1948
rect 1782 1942 1785 1948
rect 2198 1942 2201 1948
rect 2354 1948 2414 1951
rect 2438 1948 2470 1951
rect 2570 1948 2582 1951
rect 2838 1948 2894 1951
rect 2914 1948 2950 1951
rect 2954 1948 2966 1951
rect 3042 1948 3110 1951
rect 2438 1942 2441 1948
rect 2702 1942 2705 1948
rect 2838 1942 2841 1948
rect 2982 1942 2985 1948
rect 3314 1948 3358 1951
rect 3378 1948 3406 1951
rect 3462 1948 3505 1951
rect 3570 1948 3593 1951
rect 3658 1948 3662 1951
rect 3762 1948 3782 1951
rect 3874 1948 3878 1951
rect 3914 1948 4022 1951
rect 4026 1948 4030 1951
rect 4050 1948 4078 1951
rect 4090 1948 4198 1951
rect 4266 1948 4270 1951
rect 4426 1948 4438 1951
rect 4522 1948 4638 1951
rect 4650 1948 4694 1951
rect 4710 1951 4713 1958
rect 4706 1948 4713 1951
rect 4746 1948 4774 1951
rect 4810 1948 4814 1951
rect 4854 1951 4857 1958
rect 4854 1948 4862 1951
rect 18 1938 70 1941
rect 202 1938 254 1941
rect 258 1938 558 1941
rect 570 1938 681 1941
rect 802 1938 926 1941
rect 1066 1938 1086 1941
rect 1138 1938 1142 1941
rect 1162 1938 1166 1941
rect 1178 1938 1190 1941
rect 1282 1938 1294 1941
rect 1346 1938 1358 1941
rect 1362 1938 1398 1941
rect 1762 1938 1766 1941
rect 1866 1938 1886 1941
rect 1898 1938 2094 1941
rect 2298 1938 2334 1941
rect 2338 1938 2390 1941
rect 2410 1938 2422 1941
rect 2474 1938 2526 1941
rect 2570 1938 2614 1941
rect 2890 1938 2910 1941
rect 3162 1938 3230 1941
rect 3234 1938 3302 1941
rect 3366 1941 3369 1948
rect 3362 1938 3369 1941
rect 3374 1942 3377 1948
rect 3422 1942 3425 1948
rect 3462 1942 3465 1948
rect 3502 1942 3505 1948
rect 3590 1942 3593 1948
rect 3670 1942 3673 1948
rect 3386 1938 3390 1941
rect 3538 1938 3574 1941
rect 3682 1938 3838 1941
rect 3842 1938 4590 1941
rect 4594 1938 4654 1941
rect 4658 1938 4678 1941
rect 4698 1938 4822 1941
rect 5170 1938 5174 1941
rect 678 1932 681 1938
rect 250 1928 342 1931
rect 490 1928 654 1931
rect 762 1928 814 1931
rect 1486 1931 1489 1938
rect 818 1928 1489 1931
rect 1618 1928 1646 1931
rect 1850 1928 1902 1931
rect 1914 1928 2030 1931
rect 2162 1928 2422 1931
rect 2434 1928 2454 1931
rect 2618 1928 2710 1931
rect 2958 1931 2961 1938
rect 3534 1932 3537 1938
rect 2730 1928 2961 1931
rect 3058 1928 3350 1931
rect 3362 1928 3390 1931
rect 3490 1928 3526 1931
rect 3546 1928 3558 1931
rect 3682 1928 3758 1931
rect 3794 1928 3798 1931
rect 3834 1928 3838 1931
rect 3866 1928 3894 1931
rect 3962 1928 3982 1931
rect 4018 1928 4102 1931
rect 4130 1928 4182 1931
rect 4322 1928 4350 1931
rect 4386 1928 4390 1931
rect 4434 1928 4462 1931
rect 4618 1928 4702 1931
rect 4754 1928 4878 1931
rect 4882 1928 5062 1931
rect 5154 1928 5174 1931
rect 226 1918 294 1921
rect 438 1921 441 1928
rect 4574 1922 4577 1928
rect 314 1918 441 1921
rect 450 1918 486 1921
rect 550 1918 798 1921
rect 810 1918 814 1921
rect 946 1918 958 1921
rect 962 1918 1094 1921
rect 1106 1918 1414 1921
rect 1490 1918 1606 1921
rect 1626 1918 1990 1921
rect 1994 1918 2217 1921
rect 2418 1918 2422 1921
rect 2538 1918 2710 1921
rect 2794 1918 3174 1921
rect 3178 1918 4038 1921
rect 4298 1918 4342 1921
rect 4386 1918 4526 1921
rect 4618 1918 4726 1921
rect 4962 1918 4998 1921
rect 550 1911 553 1918
rect 418 1908 553 1911
rect 562 1908 606 1911
rect 738 1908 758 1911
rect 786 1908 854 1911
rect 1226 1908 1230 1911
rect 1282 1908 1526 1911
rect 1770 1908 1862 1911
rect 1882 1908 2022 1911
rect 2214 1911 2217 1918
rect 2214 1908 2286 1911
rect 2486 1908 2646 1911
rect 2810 1908 3006 1911
rect 3066 1908 3078 1911
rect 3154 1908 3262 1911
rect 3338 1908 3358 1911
rect 3482 1908 3574 1911
rect 3610 1908 3630 1911
rect 3938 1908 4054 1911
rect 4394 1908 4398 1911
rect 4410 1908 4542 1911
rect 4674 1908 4710 1911
rect 4714 1908 4782 1911
rect 4970 1908 5078 1911
rect 5146 1908 5174 1911
rect 1048 1903 1050 1907
rect 1054 1903 1057 1907
rect 1062 1903 1064 1907
rect 2072 1903 2074 1907
rect 2078 1903 2081 1907
rect 2086 1903 2088 1907
rect 162 1898 302 1901
rect 386 1898 462 1901
rect 690 1898 1030 1901
rect 1218 1898 1366 1901
rect 1530 1898 1734 1901
rect 1738 1898 1894 1901
rect 1906 1898 2054 1901
rect 2098 1898 2110 1901
rect 2114 1898 2190 1901
rect 2274 1898 2318 1901
rect 2486 1901 2489 1908
rect 3096 1903 3098 1907
rect 3102 1903 3105 1907
rect 3110 1903 3112 1907
rect 4112 1903 4114 1907
rect 4118 1903 4121 1907
rect 4126 1903 4128 1907
rect 2322 1898 2489 1901
rect 2498 1898 2638 1901
rect 2810 1898 3030 1901
rect 3082 1898 3086 1901
rect 3138 1898 3142 1901
rect 3234 1898 3262 1901
rect 3442 1898 3486 1901
rect 3498 1898 3542 1901
rect 3826 1898 3838 1901
rect 3874 1898 3886 1901
rect 3890 1898 4070 1901
rect 4098 1898 4102 1901
rect 4282 1898 4366 1901
rect 4394 1898 4438 1901
rect 4442 1898 4462 1901
rect 4490 1898 4798 1901
rect 4802 1898 4854 1901
rect 378 1888 406 1891
rect 410 1888 422 1891
rect 754 1888 790 1891
rect 1066 1888 1182 1891
rect 1186 1888 1430 1891
rect 1498 1888 1598 1891
rect 1602 1888 1718 1891
rect 1738 1888 1966 1891
rect 2010 1888 2350 1891
rect 2378 1888 2382 1891
rect 2434 1888 2438 1891
rect 2450 1888 2750 1891
rect 2794 1888 2926 1891
rect 3082 1888 3134 1891
rect 3266 1888 3366 1891
rect 3418 1888 4062 1891
rect 4082 1888 4342 1891
rect 4442 1888 4478 1891
rect 4658 1888 4822 1891
rect 4978 1888 5006 1891
rect 10 1878 134 1881
rect 174 1881 177 1888
rect 138 1878 169 1881
rect 174 1878 390 1881
rect 498 1878 662 1881
rect 842 1878 993 1881
rect 166 1872 169 1878
rect 242 1868 374 1871
rect 378 1868 398 1871
rect 450 1868 574 1871
rect 602 1868 654 1871
rect 658 1868 702 1871
rect 762 1868 766 1871
rect 794 1868 798 1871
rect 990 1871 993 1878
rect 1154 1878 1158 1881
rect 1378 1878 1502 1881
rect 1586 1878 1590 1881
rect 1594 1878 2038 1881
rect 2098 1878 2142 1881
rect 2298 1878 2358 1881
rect 2362 1878 2590 1881
rect 2706 1878 2806 1881
rect 2922 1878 3022 1881
rect 3034 1878 3054 1881
rect 3058 1878 3214 1881
rect 3538 1878 3550 1881
rect 3554 1878 3598 1881
rect 3642 1878 3678 1881
rect 3802 1878 3806 1881
rect 3818 1878 3822 1881
rect 3826 1878 3870 1881
rect 4062 1881 4065 1888
rect 5142 1882 5145 1888
rect 3906 1878 4001 1881
rect 4062 1878 4238 1881
rect 4242 1878 4270 1881
rect 4410 1878 4526 1881
rect 4626 1878 4742 1881
rect 4842 1878 4854 1881
rect 1022 1871 1025 1878
rect 990 1868 1174 1871
rect 1210 1868 1214 1871
rect 1226 1868 1230 1871
rect 1326 1868 1345 1871
rect 1426 1868 1446 1871
rect 1474 1868 1478 1871
rect 1602 1868 1614 1871
rect 1642 1868 1742 1871
rect 1810 1868 1814 1871
rect 1834 1868 1846 1871
rect 1866 1868 2086 1871
rect 2230 1871 2233 1878
rect 2138 1868 2233 1871
rect 2354 1868 2409 1871
rect 2426 1868 2566 1871
rect 2590 1871 2593 1878
rect 2590 1868 2630 1871
rect 2634 1868 2678 1871
rect 2702 1871 2705 1878
rect 3998 1872 4001 1878
rect 4326 1872 4329 1878
rect 5014 1872 5017 1878
rect 2682 1868 2705 1871
rect 2802 1868 2806 1871
rect 2874 1868 2886 1871
rect 2914 1868 3006 1871
rect 3034 1868 3134 1871
rect 3178 1868 3182 1871
rect 3186 1868 3254 1871
rect 3498 1868 3550 1871
rect 3562 1868 3574 1871
rect 3578 1868 3582 1871
rect 3594 1868 3878 1871
rect 3898 1868 3974 1871
rect 4066 1868 4094 1871
rect 4170 1868 4174 1871
rect 4210 1868 4286 1871
rect 4370 1868 4454 1871
rect 4482 1868 4486 1871
rect 4554 1868 4678 1871
rect 4714 1868 4718 1871
rect 4722 1868 4782 1871
rect 5102 1871 5105 1878
rect 5058 1868 5118 1871
rect 70 1858 102 1861
rect 162 1858 190 1861
rect 222 1861 225 1868
rect 194 1858 225 1861
rect 402 1858 406 1861
rect 466 1858 470 1861
rect 570 1858 646 1861
rect 666 1859 718 1861
rect 662 1858 718 1859
rect 982 1861 985 1868
rect 1326 1862 1329 1868
rect 1342 1862 1345 1868
rect 890 1858 985 1861
rect 1010 1858 1014 1861
rect 1090 1858 1198 1861
rect 1234 1858 1321 1861
rect 1534 1861 1537 1868
rect 1854 1862 1857 1868
rect 2406 1862 2409 1868
rect 1514 1858 1537 1861
rect 1570 1858 1654 1861
rect 1738 1858 1750 1861
rect 1770 1858 1774 1861
rect 1818 1858 1830 1861
rect 1842 1858 1846 1861
rect 1922 1858 1926 1861
rect 1946 1858 2022 1861
rect 2026 1858 2062 1861
rect 2066 1858 2102 1861
rect 2210 1858 2214 1861
rect 2282 1858 2326 1861
rect 2354 1858 2366 1861
rect 2370 1858 2382 1861
rect 2458 1858 2486 1861
rect 2618 1858 3118 1861
rect 3154 1858 3158 1861
rect 3170 1858 3198 1861
rect 3250 1858 3337 1861
rect 3394 1858 3494 1861
rect 3658 1858 3734 1861
rect 3786 1858 4510 1861
rect 4514 1858 4534 1861
rect 4538 1858 4814 1861
rect 4850 1858 5118 1861
rect 5122 1858 5166 1861
rect 70 1852 73 1858
rect 114 1848 142 1851
rect 274 1848 446 1851
rect 450 1848 478 1851
rect 698 1848 710 1851
rect 738 1848 766 1851
rect 774 1851 777 1858
rect 774 1848 814 1851
rect 1002 1848 1038 1851
rect 1082 1848 1126 1851
rect 1234 1848 1241 1851
rect 1238 1842 1241 1848
rect 1318 1851 1321 1858
rect 2142 1852 2145 1858
rect 3334 1852 3337 1858
rect 4846 1852 4849 1858
rect 1318 1848 1358 1851
rect 1522 1848 1526 1851
rect 1778 1848 1782 1851
rect 1842 1848 1902 1851
rect 1914 1848 1918 1851
rect 2122 1848 2126 1851
rect 2170 1848 2334 1851
rect 2386 1848 2430 1851
rect 2478 1848 2566 1851
rect 2858 1848 2862 1851
rect 2866 1848 2918 1851
rect 2978 1848 3022 1851
rect 3042 1848 3086 1851
rect 3106 1848 3134 1851
rect 3146 1848 3150 1851
rect 3154 1848 3326 1851
rect 3450 1848 3470 1851
rect 3498 1848 3502 1851
rect 3674 1848 3830 1851
rect 3858 1848 3862 1851
rect 3970 1848 4094 1851
rect 4146 1848 4158 1851
rect 4178 1848 4182 1851
rect 4210 1848 4214 1851
rect 4218 1848 4310 1851
rect 4434 1848 4454 1851
rect 4482 1848 4486 1851
rect 4562 1848 4574 1851
rect 4746 1848 4750 1851
rect 4810 1848 4814 1851
rect 4818 1848 4838 1851
rect 4866 1848 4870 1851
rect 4914 1848 4950 1851
rect 4970 1848 5102 1851
rect 130 1838 422 1841
rect 426 1838 454 1841
rect 778 1838 782 1841
rect 922 1838 1214 1841
rect 1254 1841 1257 1848
rect 1254 1838 1414 1841
rect 1482 1838 1937 1841
rect 2118 1841 2121 1848
rect 2478 1842 2481 1848
rect 2090 1838 2121 1841
rect 2130 1838 2246 1841
rect 2426 1838 2430 1841
rect 2490 1838 2721 1841
rect 3038 1841 3041 1848
rect 2906 1838 3041 1841
rect 3046 1838 3110 1841
rect 3378 1838 3638 1841
rect 3642 1838 3678 1841
rect 3722 1838 3902 1841
rect 4122 1838 4150 1841
rect 4170 1838 4454 1841
rect 4522 1838 4577 1841
rect 4714 1838 4753 1841
rect 10 1828 502 1831
rect 802 1828 1038 1831
rect 1130 1828 1134 1831
rect 1438 1831 1441 1838
rect 1934 1832 1937 1838
rect 2718 1832 2721 1838
rect 1438 1828 1894 1831
rect 1914 1828 1926 1831
rect 1938 1828 2038 1831
rect 2074 1828 2614 1831
rect 2722 1828 2750 1831
rect 2754 1828 3014 1831
rect 3046 1831 3049 1838
rect 4574 1832 4577 1838
rect 4750 1832 4753 1838
rect 4822 1838 4910 1841
rect 4822 1832 4825 1838
rect 3026 1828 3049 1831
rect 3082 1828 3182 1831
rect 3194 1828 3582 1831
rect 3594 1828 4094 1831
rect 4282 1828 4374 1831
rect 4410 1828 4438 1831
rect 4842 1828 4958 1831
rect 266 1818 278 1821
rect 282 1818 326 1821
rect 330 1818 446 1821
rect 450 1818 750 1821
rect 754 1818 958 1821
rect 962 1818 1078 1821
rect 1082 1818 1086 1821
rect 1106 1818 1278 1821
rect 1282 1818 1414 1821
rect 1474 1818 1478 1821
rect 1490 1818 3174 1821
rect 3426 1818 3614 1821
rect 3618 1818 3646 1821
rect 3938 1818 3958 1821
rect 4038 1818 4046 1821
rect 4050 1818 4542 1821
rect 4562 1818 4582 1821
rect 4706 1818 4806 1821
rect 210 1808 470 1811
rect 1122 1808 1190 1811
rect 1218 1808 1246 1811
rect 1506 1808 1526 1811
rect 1898 1808 2182 1811
rect 2226 1808 2502 1811
rect 3034 1808 3542 1811
rect 3698 1808 4318 1811
rect 4386 1808 4566 1811
rect 4778 1808 5062 1811
rect 536 1803 538 1807
rect 542 1803 545 1807
rect 550 1803 552 1807
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1574 1803 1576 1807
rect 2584 1803 2586 1807
rect 2590 1803 2593 1807
rect 2598 1803 2600 1807
rect 3608 1803 3610 1807
rect 3614 1803 3617 1807
rect 3622 1803 3624 1807
rect 4632 1803 4634 1807
rect 4638 1803 4641 1807
rect 4646 1803 4648 1807
rect 170 1798 446 1801
rect 818 1798 838 1801
rect 1242 1798 1494 1801
rect 1890 1798 1934 1801
rect 1962 1798 1990 1801
rect 2066 1798 2526 1801
rect 2842 1798 2854 1801
rect 2938 1798 3558 1801
rect 3682 1798 3790 1801
rect 3962 1798 3974 1801
rect 4098 1798 4222 1801
rect 4370 1798 4582 1801
rect 4666 1798 5078 1801
rect 474 1788 1118 1791
rect 1218 1788 1294 1791
rect 1322 1788 1510 1791
rect 1546 1788 1758 1791
rect 1762 1788 2654 1791
rect 2934 1788 3102 1791
rect 3202 1788 3270 1791
rect 3274 1788 3406 1791
rect 3602 1788 3646 1791
rect 3650 1788 3750 1791
rect 3986 1788 4014 1791
rect 4058 1788 4070 1791
rect 4226 1788 4246 1791
rect 4298 1788 4326 1791
rect 4338 1788 4502 1791
rect 4578 1788 4742 1791
rect 4746 1788 4886 1791
rect 318 1781 321 1788
rect 2934 1782 2937 1788
rect 318 1778 358 1781
rect 874 1778 1190 1781
rect 1258 1778 1262 1781
rect 1298 1778 1366 1781
rect 1546 1778 1678 1781
rect 1714 1778 1718 1781
rect 1730 1778 1870 1781
rect 1906 1778 1958 1781
rect 2082 1778 2206 1781
rect 2434 1778 2518 1781
rect 2522 1778 2550 1781
rect 2554 1778 2622 1781
rect 2642 1778 2734 1781
rect 3018 1778 3046 1781
rect 3066 1778 3126 1781
rect 3386 1778 3422 1781
rect 3522 1778 3574 1781
rect 3610 1778 3662 1781
rect 3666 1778 3782 1781
rect 3810 1778 4022 1781
rect 4026 1778 4062 1781
rect 4066 1778 4086 1781
rect 4090 1778 4206 1781
rect 4210 1778 4350 1781
rect 4378 1778 4630 1781
rect 4834 1778 4918 1781
rect 490 1768 542 1771
rect 882 1768 1350 1771
rect 1370 1768 1526 1771
rect 1666 1768 1878 1771
rect 1882 1768 1982 1771
rect 2050 1768 2310 1771
rect 2434 1768 2462 1771
rect 2626 1768 2782 1771
rect 2938 1768 2990 1771
rect 2994 1768 2998 1771
rect 3058 1768 3758 1771
rect 3834 1768 3982 1771
rect 3986 1768 4062 1771
rect 4078 1768 4470 1771
rect 4602 1768 4758 1771
rect 4774 1771 4777 1778
rect 4774 1768 4862 1771
rect 4922 1768 4950 1771
rect 266 1758 342 1761
rect 658 1758 702 1761
rect 714 1758 734 1761
rect 1422 1758 1550 1761
rect 1754 1758 1774 1761
rect 1778 1758 1790 1761
rect 2414 1761 2417 1768
rect 4078 1762 4081 1768
rect 4438 1762 4441 1768
rect 4590 1762 4593 1768
rect 2266 1758 2417 1761
rect 2562 1758 2662 1761
rect 2914 1758 2942 1761
rect 2986 1758 2990 1761
rect 3530 1758 3553 1761
rect 3562 1758 3574 1761
rect 3586 1758 3630 1761
rect 3634 1758 4006 1761
rect 4018 1758 4038 1761
rect 4146 1758 4206 1761
rect 4218 1758 4222 1761
rect 4266 1758 4286 1761
rect 4462 1758 4470 1761
rect 4474 1758 4534 1761
rect 4594 1758 4614 1761
rect 4806 1758 4814 1761
rect 4818 1758 4889 1761
rect 4898 1758 4926 1761
rect 5082 1758 5102 1761
rect 218 1748 382 1751
rect 430 1751 433 1758
rect 430 1748 510 1751
rect 706 1748 710 1751
rect 714 1748 718 1751
rect 774 1751 777 1758
rect 1158 1751 1161 1758
rect 1422 1752 1425 1758
rect 762 1748 777 1751
rect 958 1748 1161 1751
rect 1178 1748 1182 1751
rect 1258 1748 1286 1751
rect 1290 1748 1406 1751
rect 1578 1748 1662 1751
rect 1686 1751 1689 1758
rect 1686 1748 1737 1751
rect 86 1741 89 1748
rect 574 1742 577 1748
rect 734 1742 737 1748
rect 958 1742 961 1748
rect 1206 1742 1209 1748
rect 66 1738 158 1741
rect 162 1738 182 1741
rect 378 1738 382 1741
rect 482 1738 486 1741
rect 498 1738 518 1741
rect 642 1738 686 1741
rect 690 1738 721 1741
rect 746 1738 902 1741
rect 1026 1738 1102 1741
rect 1114 1738 1118 1741
rect 1218 1738 1262 1741
rect 1282 1738 1286 1741
rect 1322 1738 1382 1741
rect 1386 1738 1398 1741
rect 1410 1738 1430 1741
rect 1478 1741 1481 1748
rect 1734 1742 1737 1748
rect 1862 1751 1865 1758
rect 1778 1748 1865 1751
rect 1870 1752 1873 1758
rect 1918 1751 1921 1758
rect 1890 1748 2198 1751
rect 2234 1748 2238 1751
rect 2410 1748 2414 1751
rect 2438 1751 2441 1758
rect 2434 1748 2441 1751
rect 2462 1751 2465 1758
rect 2958 1752 2961 1758
rect 3070 1752 3073 1758
rect 3270 1752 3273 1758
rect 2462 1748 2478 1751
rect 2490 1748 2494 1751
rect 2506 1748 2542 1751
rect 2546 1748 2566 1751
rect 2658 1748 2718 1751
rect 2738 1748 2742 1751
rect 2866 1748 2918 1751
rect 2986 1748 2990 1751
rect 3002 1748 3062 1751
rect 3138 1748 3166 1751
rect 3194 1748 3222 1751
rect 3342 1751 3345 1758
rect 3342 1748 3374 1751
rect 3398 1751 3401 1758
rect 3454 1752 3457 1758
rect 3502 1752 3505 1758
rect 3398 1748 3406 1751
rect 3514 1748 3542 1751
rect 3550 1751 3553 1758
rect 4302 1752 4305 1758
rect 4382 1752 4385 1758
rect 3550 1748 3646 1751
rect 3658 1748 3662 1751
rect 3706 1748 3774 1751
rect 3810 1748 3814 1751
rect 3826 1748 3838 1751
rect 3994 1748 4030 1751
rect 4106 1748 4230 1751
rect 4418 1748 4430 1751
rect 4474 1748 4478 1751
rect 4498 1748 4590 1751
rect 4610 1748 4790 1751
rect 4886 1751 4889 1758
rect 5182 1752 5185 1758
rect 4886 1748 5014 1751
rect 1750 1742 1753 1748
rect 1478 1738 1614 1741
rect 1618 1738 1718 1741
rect 1922 1738 2022 1741
rect 2034 1738 2102 1741
rect 2106 1738 2134 1741
rect 2138 1738 2166 1741
rect 2226 1738 2230 1741
rect 2234 1738 2278 1741
rect 2390 1741 2393 1748
rect 2390 1738 2646 1741
rect 2706 1738 2710 1741
rect 2818 1738 2958 1741
rect 2966 1741 2969 1748
rect 2966 1738 3238 1741
rect 3242 1738 3270 1741
rect 3274 1738 3534 1741
rect 3538 1738 4806 1741
rect 4826 1738 4910 1741
rect 4918 1738 4934 1741
rect 4970 1738 5078 1741
rect 5082 1738 5110 1741
rect 5138 1738 5150 1741
rect 186 1728 214 1731
rect 222 1731 225 1738
rect 718 1732 721 1738
rect 222 1728 694 1731
rect 898 1728 982 1731
rect 1034 1728 1086 1731
rect 1098 1728 1118 1731
rect 1282 1728 1286 1731
rect 1446 1731 1449 1738
rect 4918 1732 4921 1738
rect 1446 1728 1486 1731
rect 1498 1728 1502 1731
rect 1618 1728 1702 1731
rect 1810 1728 1926 1731
rect 2002 1728 2078 1731
rect 2082 1728 2089 1731
rect 2114 1728 2190 1731
rect 2202 1728 2214 1731
rect 2218 1728 2278 1731
rect 2426 1728 2430 1731
rect 2434 1728 2510 1731
rect 2890 1728 2982 1731
rect 2986 1728 3014 1731
rect 3026 1728 3062 1731
rect 3210 1728 3214 1731
rect 3234 1728 3310 1731
rect 3402 1728 3430 1731
rect 3458 1728 3462 1731
rect 3498 1728 3662 1731
rect 3666 1728 3686 1731
rect 3754 1728 3798 1731
rect 3802 1728 3833 1731
rect 3914 1728 4118 1731
rect 4298 1728 4422 1731
rect 4578 1728 4582 1731
rect 4610 1728 4718 1731
rect 4730 1728 4846 1731
rect 4978 1728 5110 1731
rect 2374 1722 2377 1728
rect 3830 1722 3833 1728
rect 130 1718 169 1721
rect 362 1718 518 1721
rect 682 1718 686 1721
rect 706 1718 910 1721
rect 962 1718 1102 1721
rect 1274 1718 1358 1721
rect 1378 1718 1726 1721
rect 1746 1718 2214 1721
rect 2418 1718 2422 1721
rect 2810 1718 3182 1721
rect 3194 1718 3222 1721
rect 3274 1718 3278 1721
rect 3386 1718 3390 1721
rect 3394 1718 3422 1721
rect 3754 1718 3758 1721
rect 3834 1718 4078 1721
rect 4106 1718 4118 1721
rect 4290 1718 4414 1721
rect 4570 1718 4582 1721
rect 4714 1718 4782 1721
rect 4786 1718 4830 1721
rect 4922 1718 4958 1721
rect 166 1712 169 1718
rect 3790 1712 3793 1718
rect 3814 1712 3817 1718
rect 578 1708 758 1711
rect 770 1708 886 1711
rect 954 1708 982 1711
rect 1114 1708 1262 1711
rect 1306 1708 1470 1711
rect 1482 1708 1745 1711
rect 1794 1708 1798 1711
rect 1890 1708 1950 1711
rect 2138 1708 2614 1711
rect 2618 1708 2774 1711
rect 2786 1708 2870 1711
rect 2946 1708 2998 1711
rect 3034 1708 3038 1711
rect 3146 1708 3518 1711
rect 3530 1708 3758 1711
rect 3922 1708 3998 1711
rect 4226 1708 4286 1711
rect 4306 1708 4310 1711
rect 4762 1708 4798 1711
rect 4802 1708 4806 1711
rect 5026 1708 5150 1711
rect 1048 1703 1050 1707
rect 1054 1703 1057 1707
rect 1062 1703 1064 1707
rect 1742 1702 1745 1708
rect 2072 1703 2074 1707
rect 2078 1703 2081 1707
rect 2086 1703 2088 1707
rect 3096 1703 3098 1707
rect 3102 1703 3105 1707
rect 3110 1703 3112 1707
rect 4112 1703 4114 1707
rect 4118 1703 4121 1707
rect 4126 1703 4128 1707
rect 82 1698 270 1701
rect 330 1698 422 1701
rect 498 1698 670 1701
rect 818 1698 982 1701
rect 986 1698 1030 1701
rect 1202 1698 1326 1701
rect 1610 1698 1662 1701
rect 1746 1698 1798 1701
rect 1970 1698 1974 1701
rect 2826 1698 2846 1701
rect 2858 1698 2966 1701
rect 3178 1698 3230 1701
rect 3290 1698 3454 1701
rect 3514 1698 3686 1701
rect 3770 1698 3966 1701
rect 3986 1698 3990 1701
rect 4002 1698 4070 1701
rect 4230 1698 4294 1701
rect 4386 1698 4462 1701
rect 4514 1698 4782 1701
rect 4802 1698 4814 1701
rect 5026 1698 5030 1701
rect 1862 1692 1865 1698
rect 4230 1692 4233 1698
rect 194 1688 494 1691
rect 750 1688 758 1691
rect 762 1688 838 1691
rect 946 1688 950 1691
rect 1058 1688 1190 1691
rect 1202 1688 1206 1691
rect 1250 1688 1302 1691
rect 1314 1688 1422 1691
rect 1442 1688 1454 1691
rect 1522 1688 1822 1691
rect 1874 1688 2009 1691
rect 2014 1688 2022 1691
rect 2026 1688 2086 1691
rect 2106 1688 2166 1691
rect 2178 1688 2190 1691
rect 2214 1688 2222 1691
rect 2226 1688 2318 1691
rect 2442 1688 2478 1691
rect 2554 1688 2670 1691
rect 2738 1688 2766 1691
rect 2970 1688 2974 1691
rect 2978 1688 3086 1691
rect 3114 1688 3126 1691
rect 3170 1688 3174 1691
rect 3178 1688 3262 1691
rect 3418 1688 3486 1691
rect 3490 1688 3606 1691
rect 3650 1688 3654 1691
rect 3730 1688 3742 1691
rect 3858 1688 3926 1691
rect 4010 1688 4022 1691
rect 4114 1688 4150 1691
rect 4210 1688 4214 1691
rect 4226 1688 4230 1691
rect 4282 1688 4318 1691
rect 4418 1688 4478 1691
rect 4538 1688 4614 1691
rect 4690 1688 4702 1691
rect 4706 1688 4854 1691
rect 4866 1688 4950 1691
rect 4954 1688 5081 1691
rect 162 1678 262 1681
rect 266 1678 374 1681
rect 378 1678 398 1681
rect 442 1678 446 1681
rect 474 1678 494 1681
rect 510 1678 766 1681
rect 826 1678 926 1681
rect 930 1678 966 1681
rect 1106 1678 1134 1681
rect 1138 1678 1166 1681
rect 1210 1678 1462 1681
rect 1466 1678 1894 1681
rect 1906 1678 1998 1681
rect 2006 1681 2009 1688
rect 2006 1678 2038 1681
rect 2042 1678 2126 1681
rect 2138 1678 2150 1681
rect 2186 1678 2190 1681
rect 2250 1678 2262 1681
rect 2266 1678 2350 1681
rect 2394 1678 2406 1681
rect 2410 1678 2502 1681
rect 2634 1678 2646 1681
rect 2650 1678 2750 1681
rect 2770 1678 2870 1681
rect 3026 1678 3046 1681
rect 3074 1678 3126 1681
rect 3158 1681 3161 1688
rect 3798 1682 3801 1688
rect 3990 1682 3993 1688
rect 5078 1682 5081 1688
rect 3138 1678 3206 1681
rect 3650 1678 3758 1681
rect 3858 1678 3990 1681
rect 4002 1678 4086 1681
rect 4090 1678 4118 1681
rect 4194 1678 4334 1681
rect 4426 1678 4502 1681
rect 4514 1678 4638 1681
rect 4682 1678 4729 1681
rect 4738 1678 4806 1681
rect 510 1672 513 1678
rect 782 1672 785 1678
rect 98 1668 110 1671
rect 338 1668 358 1671
rect 386 1668 486 1671
rect 578 1668 582 1671
rect 610 1668 686 1671
rect 1026 1668 1046 1671
rect 1098 1668 1102 1671
rect 1118 1668 1230 1671
rect 1242 1668 1286 1671
rect 1306 1668 1334 1671
rect 1682 1668 1750 1671
rect 1778 1668 2094 1671
rect 2130 1668 2254 1671
rect 2394 1668 2398 1671
rect 2450 1668 2454 1671
rect 2578 1668 2777 1671
rect 2786 1668 2790 1671
rect 2958 1671 2961 1678
rect 2958 1668 3062 1671
rect 3090 1668 3118 1671
rect 3122 1668 3326 1671
rect 3386 1668 3494 1671
rect 3498 1668 3510 1671
rect 3706 1668 3718 1671
rect 3770 1668 3806 1671
rect 3814 1671 3817 1678
rect 3814 1668 3846 1671
rect 3874 1668 4270 1671
rect 4274 1668 4294 1671
rect 4394 1668 4406 1671
rect 4554 1668 4558 1671
rect 4610 1668 4622 1671
rect 4634 1668 4638 1671
rect 4726 1671 4729 1678
rect 4726 1668 4766 1671
rect 4786 1668 4958 1671
rect 5054 1671 5057 1678
rect 5054 1668 5062 1671
rect 926 1662 929 1668
rect 274 1658 286 1661
rect 338 1658 382 1661
rect 434 1658 470 1661
rect 650 1658 657 1661
rect 674 1658 702 1661
rect 706 1658 766 1661
rect 810 1658 865 1661
rect 914 1658 918 1661
rect 986 1658 1006 1661
rect 1118 1661 1121 1668
rect 1042 1658 1121 1661
rect 1250 1658 1262 1661
rect 1266 1658 1278 1661
rect 1334 1658 1366 1661
rect 1374 1661 1377 1668
rect 1374 1658 1446 1661
rect 1478 1661 1481 1668
rect 1478 1658 1486 1661
rect 1506 1658 1526 1661
rect 1682 1658 1726 1661
rect 1750 1658 1766 1661
rect 1810 1658 1814 1661
rect 1818 1658 1870 1661
rect 1890 1658 1894 1661
rect 1898 1658 1926 1661
rect 1986 1658 2030 1661
rect 2090 1658 2150 1661
rect 2178 1658 2222 1661
rect 2258 1658 2430 1661
rect 2690 1658 2734 1661
rect 2774 1661 2777 1668
rect 2774 1658 2910 1661
rect 2954 1658 2966 1661
rect 2994 1658 3006 1661
rect 3010 1658 3374 1661
rect 3386 1658 3446 1661
rect 3450 1658 3838 1661
rect 3854 1661 3857 1668
rect 3854 1659 3910 1661
rect 4446 1662 4449 1668
rect 3854 1658 3913 1659
rect 3970 1658 3990 1661
rect 4058 1658 4366 1661
rect 4454 1661 4457 1668
rect 4670 1662 4673 1668
rect 4718 1662 4721 1668
rect 4454 1658 4470 1661
rect 4498 1658 4566 1661
rect 4578 1658 4582 1661
rect 4738 1658 4750 1661
rect 4782 1658 4838 1661
rect 614 1652 617 1658
rect 654 1652 657 1658
rect 862 1652 865 1658
rect 378 1648 454 1651
rect 586 1648 598 1651
rect 666 1648 710 1651
rect 938 1648 950 1651
rect 1002 1648 1006 1651
rect 1050 1648 1070 1651
rect 1114 1648 1174 1651
rect 1182 1651 1185 1658
rect 1178 1648 1185 1651
rect 1334 1652 1337 1658
rect 1750 1652 1753 1658
rect 4438 1652 4441 1658
rect 1450 1648 1462 1651
rect 1602 1648 1702 1651
rect 1730 1648 1734 1651
rect 1882 1648 1934 1651
rect 2026 1648 2046 1651
rect 2158 1648 2294 1651
rect 2354 1648 2374 1651
rect 2474 1648 2566 1651
rect 2722 1648 2726 1651
rect 2882 1648 3030 1651
rect 3034 1648 3038 1651
rect 3066 1648 3222 1651
rect 3226 1648 3233 1651
rect 3282 1648 3302 1651
rect 3434 1648 3438 1651
rect 3546 1648 3585 1651
rect 2150 1642 2153 1648
rect 2158 1642 2161 1648
rect 2422 1642 2425 1648
rect 3582 1642 3585 1648
rect 3642 1648 3673 1651
rect 3770 1648 3774 1651
rect 3794 1648 3806 1651
rect 3810 1648 4142 1651
rect 4154 1648 4198 1651
rect 4354 1648 4358 1651
rect 4586 1648 4598 1651
rect 4658 1648 4678 1651
rect 4758 1648 4766 1651
rect 4782 1651 4785 1658
rect 5070 1652 5073 1658
rect 4770 1648 4785 1651
rect 4794 1648 4846 1651
rect 5058 1648 5070 1651
rect 3630 1642 3633 1648
rect 3670 1642 3673 1648
rect 362 1638 374 1641
rect 378 1638 486 1641
rect 618 1638 662 1641
rect 698 1638 710 1641
rect 738 1638 950 1641
rect 1178 1638 1214 1641
rect 1442 1638 1510 1641
rect 1666 1638 2094 1641
rect 2098 1638 2142 1641
rect 2322 1638 2366 1641
rect 2434 1638 3174 1641
rect 3274 1638 3278 1641
rect 3302 1638 3310 1641
rect 3314 1638 3558 1641
rect 3838 1638 3846 1641
rect 3850 1638 3974 1641
rect 4018 1638 4166 1641
rect 4290 1638 4382 1641
rect 4650 1638 4726 1641
rect 4842 1638 4926 1641
rect 4942 1641 4945 1648
rect 4942 1638 5150 1641
rect 670 1632 673 1638
rect 258 1628 518 1631
rect 610 1628 622 1631
rect 706 1628 790 1631
rect 794 1628 814 1631
rect 818 1628 1110 1631
rect 1178 1628 1262 1631
rect 1698 1628 1718 1631
rect 1722 1628 1790 1631
rect 1794 1628 1878 1631
rect 1882 1628 1894 1631
rect 1898 1628 2270 1631
rect 2418 1628 3782 1631
rect 3842 1628 3910 1631
rect 4066 1628 4070 1631
rect 4422 1631 4425 1638
rect 4082 1628 4425 1631
rect 4466 1628 4654 1631
rect 4690 1628 4774 1631
rect 250 1618 758 1621
rect 786 1618 1017 1621
rect 1170 1618 2110 1621
rect 2162 1618 2590 1621
rect 2594 1618 2742 1621
rect 2946 1618 2982 1621
rect 3074 1618 3134 1621
rect 3418 1618 3814 1621
rect 3946 1618 3950 1621
rect 3954 1618 4278 1621
rect 4434 1618 4534 1621
rect 4538 1618 4734 1621
rect 4810 1618 5150 1621
rect 370 1608 422 1611
rect 594 1608 622 1611
rect 690 1608 774 1611
rect 1014 1611 1017 1618
rect 1014 1608 1318 1611
rect 1738 1608 2318 1611
rect 2402 1608 2422 1611
rect 2698 1608 2838 1611
rect 3026 1608 3070 1611
rect 3122 1608 3182 1611
rect 3218 1608 3414 1611
rect 3794 1608 3822 1611
rect 3866 1608 3910 1611
rect 4026 1608 4390 1611
rect 4658 1608 4910 1611
rect 536 1603 538 1607
rect 542 1603 545 1607
rect 550 1603 552 1607
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1574 1603 1576 1607
rect 2584 1603 2586 1607
rect 2590 1603 2593 1607
rect 2598 1603 2600 1607
rect 3608 1603 3610 1607
rect 3614 1603 3617 1607
rect 3622 1603 3624 1607
rect 4632 1603 4634 1607
rect 4638 1603 4641 1607
rect 4646 1603 4648 1607
rect 650 1598 726 1601
rect 738 1598 782 1601
rect 1074 1598 1206 1601
rect 1426 1598 1505 1601
rect 1698 1598 1702 1601
rect 1730 1598 1758 1601
rect 1778 1598 1974 1601
rect 2154 1598 2342 1601
rect 2742 1598 2998 1601
rect 3010 1598 3206 1601
rect 3314 1598 3382 1601
rect 3634 1598 4022 1601
rect 4186 1598 4246 1601
rect 4378 1598 4606 1601
rect 4874 1598 4894 1601
rect 1502 1592 1505 1598
rect 674 1588 1014 1591
rect 1018 1588 1046 1591
rect 1202 1588 1318 1591
rect 1326 1588 1334 1591
rect 1338 1588 1478 1591
rect 1506 1588 1774 1591
rect 1834 1588 1926 1591
rect 2034 1588 2078 1591
rect 2394 1588 2414 1591
rect 2742 1591 2745 1598
rect 2570 1588 2745 1591
rect 2754 1588 2982 1591
rect 3122 1588 3406 1591
rect 3410 1588 4006 1591
rect 4010 1588 4030 1591
rect 4042 1588 4054 1591
rect 4106 1588 4166 1591
rect 4250 1588 4270 1591
rect 4346 1588 4350 1591
rect 4610 1588 4654 1591
rect 4810 1588 4854 1591
rect 4878 1588 4902 1591
rect 2230 1582 2233 1588
rect 426 1578 734 1581
rect 766 1578 774 1581
rect 778 1578 1022 1581
rect 1074 1578 1078 1581
rect 1194 1578 1198 1581
rect 1322 1578 1334 1581
rect 1430 1578 1438 1581
rect 1442 1578 1534 1581
rect 1546 1578 1790 1581
rect 1794 1578 1910 1581
rect 1922 1578 1926 1581
rect 2082 1578 2102 1581
rect 2154 1578 2206 1581
rect 2286 1581 2289 1588
rect 4878 1582 4881 1588
rect 2242 1578 2289 1581
rect 2298 1578 2302 1581
rect 2314 1578 2790 1581
rect 2914 1578 2926 1581
rect 2930 1578 3118 1581
rect 3130 1578 3166 1581
rect 3178 1578 3326 1581
rect 3330 1578 3337 1581
rect 3346 1578 3350 1581
rect 3410 1578 3414 1581
rect 3498 1578 3566 1581
rect 3570 1578 3577 1581
rect 3586 1578 3622 1581
rect 3626 1578 3750 1581
rect 3754 1578 3878 1581
rect 3882 1578 4286 1581
rect 4322 1578 4414 1581
rect 106 1568 150 1571
rect 154 1568 614 1571
rect 738 1568 870 1571
rect 874 1568 942 1571
rect 1018 1568 1038 1571
rect 1050 1568 3166 1571
rect 3178 1568 4390 1571
rect 4394 1568 4550 1571
rect 4554 1568 4614 1571
rect 4802 1568 5046 1571
rect 370 1558 462 1561
rect 554 1558 614 1561
rect 618 1558 662 1561
rect 666 1558 686 1561
rect 778 1558 926 1561
rect 1002 1558 1006 1561
rect 1130 1558 1142 1561
rect 1358 1558 1366 1561
rect 1490 1558 1566 1561
rect 1602 1558 1678 1561
rect 1786 1558 1798 1561
rect 1930 1558 1950 1561
rect 1970 1558 2054 1561
rect 2106 1558 2110 1561
rect 2146 1558 2174 1561
rect 2186 1558 2190 1561
rect 2202 1558 2518 1561
rect 2530 1558 2630 1561
rect 2642 1558 2782 1561
rect 2874 1558 2886 1561
rect 3034 1558 3142 1561
rect 3146 1558 3206 1561
rect 3258 1558 3366 1561
rect 3434 1558 3470 1561
rect 3474 1558 3526 1561
rect 3626 1558 3798 1561
rect 3962 1558 3977 1561
rect 1022 1552 1025 1558
rect 50 1548 126 1551
rect 326 1548 358 1551
rect 442 1548 510 1551
rect 326 1542 329 1548
rect 406 1542 409 1548
rect 602 1548 606 1551
rect 778 1548 782 1551
rect 882 1548 894 1551
rect 922 1548 950 1551
rect 994 1548 998 1551
rect 1034 1548 1046 1551
rect 1082 1548 1086 1551
rect 1142 1548 1150 1551
rect 1162 1548 1174 1551
rect 1190 1551 1193 1558
rect 1318 1552 1321 1558
rect 1590 1552 1593 1558
rect 1702 1552 1705 1558
rect 2198 1552 2201 1558
rect 2846 1552 2849 1558
rect 1190 1548 1214 1551
rect 1410 1548 1414 1551
rect 1554 1548 1558 1551
rect 1570 1548 1574 1551
rect 1674 1548 1686 1551
rect 1738 1548 1742 1551
rect 1782 1548 1798 1551
rect 1842 1548 1846 1551
rect 1946 1548 1950 1551
rect 1978 1548 1982 1551
rect 2050 1548 2054 1551
rect 2098 1548 2150 1551
rect 2210 1548 2222 1551
rect 2234 1548 2238 1551
rect 2282 1548 2286 1551
rect 2306 1548 2310 1551
rect 2334 1548 2358 1551
rect 2366 1548 2726 1551
rect 2730 1548 2734 1551
rect 2866 1548 2870 1551
rect 2882 1548 2910 1551
rect 2914 1548 2958 1551
rect 3050 1548 3054 1551
rect 3162 1548 3246 1551
rect 3322 1548 3366 1551
rect 3538 1548 3542 1551
rect 3614 1551 3617 1558
rect 3614 1548 3646 1551
rect 3650 1548 3814 1551
rect 3854 1551 3857 1558
rect 3974 1552 3977 1558
rect 4082 1558 4230 1561
rect 4314 1558 4462 1561
rect 4642 1558 4662 1561
rect 4670 1558 4678 1561
rect 4682 1558 4710 1561
rect 4846 1558 4934 1561
rect 4938 1558 5046 1561
rect 5066 1558 5070 1561
rect 5222 1561 5226 1562
rect 5170 1558 5226 1561
rect 4054 1552 4057 1558
rect 4078 1552 4081 1558
rect 4830 1552 4833 1558
rect 4846 1552 4849 1558
rect 3850 1548 3857 1551
rect 3958 1548 3966 1551
rect 4130 1548 4142 1551
rect 4346 1548 4374 1551
rect 4530 1548 4566 1551
rect 4682 1548 4782 1551
rect 4858 1548 4894 1551
rect 4898 1548 4982 1551
rect 4986 1548 4998 1551
rect 5074 1548 5142 1551
rect 1142 1542 1145 1548
rect 106 1538 222 1541
rect 226 1538 278 1541
rect 450 1538 526 1541
rect 570 1538 582 1541
rect 642 1538 790 1541
rect 842 1538 886 1541
rect 954 1538 958 1541
rect 978 1538 1030 1541
rect 1230 1541 1233 1548
rect 1390 1542 1393 1548
rect 1470 1542 1473 1548
rect 1494 1542 1497 1548
rect 1782 1542 1785 1548
rect 2334 1542 2337 1548
rect 1154 1538 1233 1541
rect 1266 1538 1374 1541
rect 1554 1538 1598 1541
rect 1666 1538 1766 1541
rect 1882 1538 1902 1541
rect 1922 1538 2238 1541
rect 2266 1538 2286 1541
rect 2366 1541 2369 1548
rect 3958 1542 3961 1548
rect 3990 1542 3993 1548
rect 2346 1538 2369 1541
rect 2378 1538 2390 1541
rect 2626 1538 2638 1541
rect 2642 1538 2649 1541
rect 2854 1538 2870 1541
rect 2914 1538 2998 1541
rect 3010 1538 3014 1541
rect 3026 1538 3030 1541
rect 3034 1538 3062 1541
rect 3074 1538 3158 1541
rect 3194 1538 3246 1541
rect 3546 1538 3566 1541
rect 3570 1538 3590 1541
rect 3722 1538 3862 1541
rect 3906 1538 3918 1541
rect 4090 1538 4238 1541
rect 4290 1538 4398 1541
rect 4746 1538 4974 1541
rect 5018 1538 5062 1541
rect 5066 1538 5086 1541
rect 66 1528 166 1531
rect 330 1528 334 1531
rect 794 1528 1118 1531
rect 1122 1528 1126 1531
rect 1202 1528 1366 1531
rect 1370 1528 1502 1531
rect 1522 1528 1526 1531
rect 1538 1528 1566 1531
rect 1698 1528 1710 1531
rect 1922 1528 1942 1531
rect 1962 1528 2006 1531
rect 2034 1528 2094 1531
rect 2130 1528 2158 1531
rect 2210 1528 2222 1531
rect 2258 1528 2270 1531
rect 2670 1531 2673 1538
rect 2854 1532 2857 1538
rect 3342 1532 3345 1538
rect 3350 1532 3353 1538
rect 2290 1528 2750 1531
rect 2786 1528 2822 1531
rect 2898 1528 2926 1531
rect 2930 1528 2942 1531
rect 2962 1528 3022 1531
rect 3026 1528 3214 1531
rect 3242 1528 3310 1531
rect 3418 1528 3478 1531
rect 3666 1528 3686 1531
rect 3762 1528 3894 1531
rect 4106 1528 4150 1531
rect 4162 1528 4286 1531
rect 4394 1528 4814 1531
rect 4858 1528 5038 1531
rect 5042 1528 5046 1531
rect 5074 1528 5102 1531
rect 282 1518 286 1521
rect 426 1518 454 1521
rect 566 1521 569 1528
rect 670 1522 673 1528
rect 3534 1522 3537 1528
rect 474 1518 569 1521
rect 722 1518 1014 1521
rect 1018 1518 1022 1521
rect 1038 1518 1158 1521
rect 1322 1518 1782 1521
rect 1922 1518 1974 1521
rect 1994 1518 2110 1521
rect 2146 1518 2158 1521
rect 2194 1518 2214 1521
rect 2362 1518 2398 1521
rect 2402 1518 2414 1521
rect 2418 1518 2454 1521
rect 2458 1518 2486 1521
rect 2490 1518 2550 1521
rect 2698 1518 2814 1521
rect 2850 1518 2886 1521
rect 2954 1518 2998 1521
rect 3002 1518 3070 1521
rect 3086 1518 3278 1521
rect 3650 1518 3710 1521
rect 3726 1521 3729 1528
rect 3726 1518 3766 1521
rect 3810 1518 3846 1521
rect 3858 1518 3862 1521
rect 4098 1518 4150 1521
rect 4178 1518 4502 1521
rect 4626 1518 4694 1521
rect 4826 1518 5038 1521
rect 654 1512 657 1518
rect 114 1508 134 1511
rect 138 1508 174 1511
rect 178 1508 270 1511
rect 274 1508 422 1511
rect 738 1508 766 1511
rect 1038 1511 1041 1518
rect 970 1508 1041 1511
rect 1346 1508 1422 1511
rect 1522 1508 1638 1511
rect 1674 1508 1846 1511
rect 1962 1508 1990 1511
rect 2098 1508 2214 1511
rect 2266 1508 2406 1511
rect 2434 1508 2510 1511
rect 2738 1508 2790 1511
rect 2906 1508 2958 1511
rect 2962 1508 3006 1511
rect 3086 1511 3089 1518
rect 3034 1508 3089 1511
rect 3146 1508 3190 1511
rect 3674 1508 3734 1511
rect 3970 1508 4102 1511
rect 4170 1508 4766 1511
rect 4890 1508 4934 1511
rect 5002 1508 5134 1511
rect 1048 1503 1050 1507
rect 1054 1503 1057 1507
rect 1062 1503 1064 1507
rect 1166 1502 1169 1508
rect 2072 1503 2074 1507
rect 2078 1503 2081 1507
rect 2086 1503 2088 1507
rect 3096 1503 3098 1507
rect 3102 1503 3105 1507
rect 3110 1503 3112 1507
rect 4112 1503 4114 1507
rect 4118 1503 4121 1507
rect 4126 1503 4128 1507
rect 134 1498 342 1501
rect 394 1498 462 1501
rect 522 1498 622 1501
rect 938 1498 942 1501
rect 1178 1498 1390 1501
rect 1434 1498 1806 1501
rect 2122 1498 2126 1501
rect 2154 1498 2206 1501
rect 2322 1498 2342 1501
rect 2426 1498 2454 1501
rect 2466 1498 2638 1501
rect 2674 1498 2790 1501
rect 2818 1498 2854 1501
rect 2874 1498 2934 1501
rect 2938 1498 2982 1501
rect 3122 1498 3134 1501
rect 3578 1498 3670 1501
rect 4074 1498 4094 1501
rect 4138 1498 4158 1501
rect 4242 1498 4318 1501
rect 4402 1498 4742 1501
rect 4850 1498 4870 1501
rect 134 1492 137 1498
rect 94 1488 134 1491
rect 194 1488 262 1491
rect 294 1488 486 1491
rect 490 1488 494 1491
rect 578 1488 630 1491
rect 674 1488 934 1491
rect 938 1488 1150 1491
rect 1154 1488 1230 1491
rect 1234 1488 1254 1491
rect 1306 1488 1406 1491
rect 1414 1491 1417 1498
rect 5086 1492 5089 1498
rect 1414 1488 1422 1491
rect 1482 1488 1486 1491
rect 1506 1488 1510 1491
rect 1538 1488 1550 1491
rect 1682 1488 1702 1491
rect 1738 1488 1814 1491
rect 2042 1488 2126 1491
rect 2394 1488 2422 1491
rect 2442 1488 2446 1491
rect 2462 1488 2702 1491
rect 2706 1488 2750 1491
rect 2786 1488 2798 1491
rect 2874 1488 2974 1491
rect 3010 1488 3046 1491
rect 3050 1488 3094 1491
rect 3106 1488 3142 1491
rect 3162 1488 3198 1491
rect 3202 1488 3222 1491
rect 3226 1488 3270 1491
rect 3322 1488 3350 1491
rect 3394 1488 3398 1491
rect 3402 1488 3510 1491
rect 3514 1488 3542 1491
rect 3586 1488 3590 1491
rect 3594 1488 3654 1491
rect 3690 1488 3734 1491
rect 3786 1488 3918 1491
rect 3922 1488 3926 1491
rect 3938 1488 3985 1491
rect 3994 1488 3998 1491
rect 4130 1488 4334 1491
rect 4382 1488 4390 1491
rect 4394 1488 4462 1491
rect 4570 1488 4694 1491
rect 4866 1488 4878 1491
rect 5026 1488 5046 1491
rect 94 1482 97 1488
rect 294 1482 297 1488
rect 170 1478 294 1481
rect 426 1478 878 1481
rect 882 1478 1598 1481
rect 1602 1478 2166 1481
rect 2170 1478 2182 1481
rect 2250 1478 2286 1481
rect 2330 1478 2342 1481
rect 2462 1481 2465 1488
rect 2346 1478 2465 1481
rect 2506 1478 3854 1481
rect 3962 1478 3974 1481
rect 3982 1481 3985 1488
rect 3982 1478 4102 1481
rect 4194 1478 4246 1481
rect 4250 1478 4257 1481
rect 4266 1478 4486 1481
rect 4726 1481 4729 1488
rect 4942 1482 4945 1488
rect 4618 1478 4729 1481
rect 4746 1478 4750 1481
rect 4770 1478 4926 1481
rect 186 1468 270 1471
rect 398 1471 401 1478
rect 2198 1472 2201 1478
rect 398 1468 414 1471
rect 434 1468 446 1471
rect 610 1468 630 1471
rect 666 1468 670 1471
rect 706 1468 718 1471
rect 722 1468 742 1471
rect 754 1468 758 1471
rect 770 1468 774 1471
rect 930 1468 945 1471
rect 50 1458 126 1461
rect 178 1458 246 1461
rect 282 1458 318 1461
rect 322 1458 446 1461
rect 562 1458 598 1461
rect 602 1458 694 1461
rect 698 1458 790 1461
rect 810 1459 854 1461
rect 942 1462 945 1468
rect 1042 1468 1262 1471
rect 1266 1468 1646 1471
rect 1682 1468 1686 1471
rect 1794 1468 1798 1471
rect 1938 1468 1942 1471
rect 2090 1468 2102 1471
rect 2114 1468 2126 1471
rect 2162 1468 2166 1471
rect 2410 1468 2430 1471
rect 2618 1468 2638 1471
rect 2666 1468 2686 1471
rect 2778 1468 2846 1471
rect 2938 1468 3014 1471
rect 3042 1468 3046 1471
rect 3058 1468 3078 1471
rect 3082 1468 3126 1471
rect 3162 1468 3182 1471
rect 3194 1468 3206 1471
rect 3322 1468 3406 1471
rect 3442 1468 3446 1471
rect 3458 1468 3462 1471
rect 3530 1468 3718 1471
rect 3722 1468 3870 1471
rect 3874 1468 3902 1471
rect 3978 1468 4054 1471
rect 4066 1468 4158 1471
rect 4250 1468 4254 1471
rect 4322 1468 4326 1471
rect 4362 1468 4366 1471
rect 4370 1468 4406 1471
rect 4486 1471 4489 1478
rect 4486 1468 4574 1471
rect 4682 1468 4830 1471
rect 4858 1468 4862 1471
rect 4906 1468 4910 1471
rect 4934 1471 4937 1478
rect 4934 1468 5054 1471
rect 5058 1468 5065 1471
rect 958 1462 961 1468
rect 2462 1462 2465 1468
rect 3902 1462 3905 1468
rect 810 1458 857 1459
rect 1018 1458 1118 1461
rect 1138 1458 1142 1461
rect 1202 1458 1209 1461
rect 1282 1458 1302 1461
rect 1346 1458 1350 1461
rect 1418 1458 1438 1461
rect 1474 1458 1766 1461
rect 1770 1458 1774 1461
rect 1970 1458 1974 1461
rect 2042 1458 2454 1461
rect 2554 1458 2614 1461
rect 2618 1458 2646 1461
rect 2650 1458 2678 1461
rect 2762 1458 2822 1461
rect 2826 1458 2934 1461
rect 2938 1458 2958 1461
rect 2962 1458 2974 1461
rect 2978 1458 3150 1461
rect 3210 1458 3230 1461
rect 3258 1458 3374 1461
rect 3402 1458 3518 1461
rect 3554 1458 3566 1461
rect 3570 1458 3574 1461
rect 3610 1458 3630 1461
rect 3682 1458 3710 1461
rect 3714 1458 3862 1461
rect 3866 1458 3886 1461
rect 3914 1458 3934 1461
rect 3994 1458 4542 1461
rect 4690 1458 5062 1461
rect 5090 1458 5134 1461
rect 1206 1452 1209 1458
rect 218 1448 366 1451
rect 434 1448 438 1451
rect 466 1448 638 1451
rect 642 1448 646 1451
rect 882 1448 982 1451
rect 1018 1448 1030 1451
rect 1058 1448 1070 1451
rect 1110 1448 1142 1451
rect 1326 1451 1329 1458
rect 1290 1448 1329 1451
rect 1370 1448 1462 1451
rect 1466 1448 1510 1451
rect 1530 1448 1750 1451
rect 1754 1448 1758 1451
rect 1818 1448 1846 1451
rect 1874 1448 2014 1451
rect 2118 1448 2145 1451
rect 2194 1448 2198 1451
rect 2206 1448 2238 1451
rect 2250 1448 2254 1451
rect 2266 1448 2334 1451
rect 2658 1448 2686 1451
rect 2986 1448 3350 1451
rect 3362 1448 3422 1451
rect 3426 1448 3470 1451
rect 3474 1448 3646 1451
rect 3690 1448 3734 1451
rect 3866 1448 3870 1451
rect 3922 1448 3966 1451
rect 3970 1448 3990 1451
rect 4130 1448 4254 1451
rect 4306 1448 4329 1451
rect 4354 1448 4390 1451
rect 4714 1448 4734 1451
rect 4762 1448 4814 1451
rect 4822 1448 4846 1451
rect 4922 1448 4953 1451
rect 5098 1448 5110 1451
rect 1110 1442 1113 1448
rect 2094 1442 2097 1448
rect 2102 1442 2105 1448
rect 2118 1442 2121 1448
rect 2142 1442 2145 1448
rect 2206 1442 2209 1448
rect 2798 1442 2801 1448
rect 4326 1442 4329 1448
rect 4710 1442 4713 1448
rect 4822 1442 4825 1448
rect 4950 1442 4953 1448
rect 114 1438 606 1441
rect 618 1438 798 1441
rect 938 1438 966 1441
rect 1074 1438 1110 1441
rect 1394 1438 1446 1441
rect 1498 1438 1590 1441
rect 1626 1438 1678 1441
rect 1694 1438 1758 1441
rect 1826 1438 1862 1441
rect 2186 1438 2190 1441
rect 2234 1438 2294 1441
rect 2426 1438 2686 1441
rect 2970 1438 3014 1441
rect 3034 1438 3918 1441
rect 3938 1438 4134 1441
rect 4666 1438 4686 1441
rect 5026 1438 5126 1441
rect 1198 1432 1201 1438
rect 242 1428 254 1431
rect 370 1428 374 1431
rect 442 1428 702 1431
rect 786 1428 798 1431
rect 994 1428 1198 1431
rect 1226 1428 1238 1431
rect 1370 1428 1406 1431
rect 1410 1428 1521 1431
rect 1694 1431 1697 1438
rect 1554 1428 1697 1431
rect 1706 1428 1742 1431
rect 1754 1428 1790 1431
rect 1794 1428 2134 1431
rect 2186 1428 2574 1431
rect 2610 1428 2654 1431
rect 2706 1428 2918 1431
rect 2994 1428 3198 1431
rect 3338 1428 3382 1431
rect 3482 1428 3550 1431
rect 3858 1428 3886 1431
rect 3890 1428 3910 1431
rect 4050 1428 4310 1431
rect 4546 1428 4750 1431
rect 4754 1428 4814 1431
rect 4818 1428 4830 1431
rect 4962 1428 5086 1431
rect 222 1421 225 1428
rect 222 1418 310 1421
rect 378 1418 406 1421
rect 530 1418 742 1421
rect 834 1418 902 1421
rect 1098 1418 1110 1421
rect 1114 1418 1366 1421
rect 1518 1421 1521 1428
rect 1518 1418 2046 1421
rect 2090 1418 2102 1421
rect 2170 1418 2190 1421
rect 2258 1418 2350 1421
rect 2354 1418 2414 1421
rect 2702 1421 2705 1428
rect 2426 1418 2705 1421
rect 2898 1418 2910 1421
rect 3122 1418 3126 1421
rect 3154 1418 3158 1421
rect 3258 1418 3406 1421
rect 3410 1418 4142 1421
rect 4146 1418 4150 1421
rect 4338 1418 4446 1421
rect 4450 1418 4665 1421
rect 3070 1412 3073 1418
rect 170 1408 337 1411
rect 658 1408 662 1411
rect 682 1408 742 1411
rect 1162 1408 1270 1411
rect 1402 1408 1422 1411
rect 1642 1408 1758 1411
rect 1858 1408 2038 1411
rect 2058 1408 2062 1411
rect 2090 1408 2286 1411
rect 2362 1408 2486 1411
rect 2682 1408 2742 1411
rect 3114 1408 3182 1411
rect 3266 1408 3422 1411
rect 3858 1408 3950 1411
rect 4018 1408 4022 1411
rect 4042 1408 4246 1411
rect 4258 1408 4510 1411
rect 4514 1408 4534 1411
rect 4662 1411 4665 1418
rect 4782 1412 4785 1418
rect 4662 1408 4694 1411
rect 4698 1408 4766 1411
rect 4802 1408 4854 1411
rect 334 1402 337 1408
rect 536 1403 538 1407
rect 542 1403 545 1407
rect 550 1403 552 1407
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1574 1403 1576 1407
rect 2584 1403 2586 1407
rect 2590 1403 2593 1407
rect 2598 1403 2600 1407
rect 3608 1403 3610 1407
rect 3614 1403 3617 1407
rect 3622 1403 3624 1407
rect 4632 1403 4634 1407
rect 4638 1403 4641 1407
rect 4646 1403 4648 1407
rect 202 1398 230 1401
rect 234 1398 302 1401
rect 338 1398 398 1401
rect 402 1398 454 1401
rect 458 1398 526 1401
rect 570 1398 686 1401
rect 810 1398 854 1401
rect 970 1398 1238 1401
rect 1370 1398 1430 1401
rect 1442 1398 1510 1401
rect 1642 1398 1726 1401
rect 1746 1398 2118 1401
rect 2250 1398 2398 1401
rect 2402 1398 2574 1401
rect 2914 1398 3094 1401
rect 3458 1398 3494 1401
rect 3498 1398 3534 1401
rect 3826 1398 3926 1401
rect 3970 1398 4446 1401
rect 4658 1398 4758 1401
rect 126 1392 129 1398
rect 282 1388 310 1391
rect 314 1388 382 1391
rect 418 1388 422 1391
rect 482 1388 518 1391
rect 634 1388 654 1391
rect 658 1388 734 1391
rect 738 1388 758 1391
rect 762 1388 998 1391
rect 1002 1388 1214 1391
rect 1218 1388 1230 1391
rect 1234 1388 1454 1391
rect 1458 1388 2150 1391
rect 2306 1388 2470 1391
rect 2474 1388 2558 1391
rect 2562 1388 2838 1391
rect 2938 1388 3022 1391
rect 3194 1388 3286 1391
rect 3458 1388 3638 1391
rect 3650 1388 3822 1391
rect 3826 1388 3902 1391
rect 3906 1388 3934 1391
rect 4130 1388 4134 1391
rect 4234 1388 4254 1391
rect 4346 1388 4478 1391
rect 106 1378 134 1381
rect 138 1378 502 1381
rect 530 1378 1086 1381
rect 1250 1378 1638 1381
rect 1674 1378 1710 1381
rect 1906 1378 2478 1381
rect 2578 1378 2606 1381
rect 2610 1378 2918 1381
rect 2926 1381 2929 1388
rect 2926 1378 2958 1381
rect 3066 1378 3334 1381
rect 3338 1378 3390 1381
rect 3394 1378 4390 1381
rect 4394 1378 4422 1381
rect 4522 1378 4862 1381
rect 4930 1378 5030 1381
rect 226 1368 294 1371
rect 666 1368 678 1371
rect 1094 1371 1097 1378
rect 1082 1368 1097 1371
rect 1110 1368 1198 1371
rect 1202 1368 1390 1371
rect 1698 1368 1710 1371
rect 1986 1368 2070 1371
rect 2090 1368 2126 1371
rect 2202 1368 2214 1371
rect 2226 1368 2478 1371
rect 2554 1368 2558 1371
rect 2634 1368 2678 1371
rect 2690 1368 2734 1371
rect 2826 1368 2886 1371
rect 2890 1368 3190 1371
rect 3218 1368 3382 1371
rect 3434 1368 3630 1371
rect 3722 1368 3798 1371
rect 3818 1368 3838 1371
rect 4234 1368 4358 1371
rect 4850 1368 4942 1371
rect 102 1361 105 1368
rect 102 1358 134 1361
rect 154 1358 326 1361
rect 430 1361 433 1368
rect 354 1358 409 1361
rect 430 1358 462 1361
rect 598 1361 601 1368
rect 638 1361 641 1368
rect 846 1362 849 1368
rect 1110 1362 1113 1368
rect 598 1358 641 1361
rect 650 1358 806 1361
rect 834 1358 838 1361
rect 874 1358 902 1361
rect 946 1358 950 1361
rect 1034 1358 1094 1361
rect 1218 1358 1262 1361
rect 1346 1358 1350 1361
rect 1370 1358 1374 1361
rect 1410 1358 1422 1361
rect 1426 1358 1502 1361
rect 1586 1358 1606 1361
rect 1610 1358 1646 1361
rect 1666 1358 1710 1361
rect 1838 1361 1841 1368
rect 3654 1362 3657 1368
rect 1834 1358 1841 1361
rect 1978 1358 1990 1361
rect 2178 1358 2302 1361
rect 2314 1358 2318 1361
rect 2330 1358 2334 1361
rect 2418 1358 2606 1361
rect 2610 1358 2630 1361
rect 2642 1358 2646 1361
rect 2658 1358 2670 1361
rect 2722 1358 2782 1361
rect 2874 1358 2886 1361
rect 3066 1358 3078 1361
rect 3098 1358 3286 1361
rect 3290 1358 3294 1361
rect 3378 1358 3414 1361
rect 3418 1358 3438 1361
rect 3530 1358 3534 1361
rect 3666 1358 3766 1361
rect 3894 1361 3897 1368
rect 3894 1358 3966 1361
rect 4050 1358 4054 1361
rect 4190 1361 4193 1368
rect 4122 1358 4193 1361
rect 4670 1361 4673 1368
rect 4670 1358 4734 1361
rect 4986 1358 4990 1361
rect 5058 1358 5062 1361
rect 406 1352 409 1358
rect 974 1352 977 1358
rect 1102 1352 1105 1358
rect 2006 1352 2009 1358
rect 58 1348 105 1351
rect 102 1342 105 1348
rect 118 1348 294 1351
rect 298 1348 350 1351
rect 410 1348 414 1351
rect 426 1348 470 1351
rect 118 1342 121 1348
rect 570 1348 574 1351
rect 602 1348 606 1351
rect 626 1348 726 1351
rect 778 1348 854 1351
rect 874 1348 886 1351
rect 914 1348 918 1351
rect 938 1348 942 1351
rect 1018 1348 1038 1351
rect 1226 1348 1230 1351
rect 1234 1348 1390 1351
rect 1434 1348 1473 1351
rect 1546 1348 1598 1351
rect 1770 1348 1774 1351
rect 1794 1348 1830 1351
rect 1834 1348 1902 1351
rect 2014 1351 2017 1358
rect 2062 1352 2065 1358
rect 2110 1352 2113 1358
rect 3006 1352 3009 1358
rect 3830 1352 3833 1358
rect 2014 1348 2062 1351
rect 2158 1348 2222 1351
rect 2250 1348 2326 1351
rect 2330 1348 2382 1351
rect 2394 1348 2422 1351
rect 2442 1348 2486 1351
rect 2490 1348 2694 1351
rect 2698 1348 2726 1351
rect 2730 1348 2758 1351
rect 2826 1348 2838 1351
rect 2858 1348 2942 1351
rect 3170 1348 3318 1351
rect 3382 1348 3574 1351
rect 3674 1348 3678 1351
rect 3690 1348 3750 1351
rect 3906 1348 3926 1351
rect 4018 1348 4046 1351
rect 4050 1348 4054 1351
rect 4082 1348 4182 1351
rect 4186 1348 4190 1351
rect 4202 1348 4529 1351
rect 4826 1348 4886 1351
rect 4950 1351 4953 1358
rect 4906 1348 4982 1351
rect 5006 1351 5009 1358
rect 4986 1348 5009 1351
rect 5042 1348 5134 1351
rect 1470 1342 1473 1348
rect 258 1338 342 1341
rect 346 1338 350 1341
rect 418 1338 558 1341
rect 610 1338 678 1341
rect 698 1338 750 1341
rect 882 1338 886 1341
rect 890 1338 1046 1341
rect 1082 1338 1142 1341
rect 1202 1338 1222 1341
rect 1338 1338 1366 1341
rect 1390 1338 1406 1341
rect 1410 1338 1422 1341
rect 1498 1338 1550 1341
rect 1562 1338 1566 1341
rect 1630 1341 1633 1348
rect 2158 1342 2161 1348
rect 3318 1342 3321 1348
rect 3382 1342 3385 1348
rect 3502 1342 3505 1348
rect 3662 1342 3665 1348
rect 1618 1338 1798 1341
rect 1810 1338 2094 1341
rect 2330 1338 2350 1341
rect 2474 1338 2478 1341
rect 2482 1338 2494 1341
rect 2514 1338 2534 1341
rect 2554 1338 2574 1341
rect 2618 1338 2646 1341
rect 2738 1338 2742 1341
rect 2850 1338 2870 1341
rect 2874 1338 3134 1341
rect 3138 1338 3198 1341
rect 3218 1338 3222 1341
rect 3770 1338 3838 1341
rect 3898 1338 3902 1341
rect 3974 1338 4030 1341
rect 4042 1338 4057 1341
rect 4090 1338 4206 1341
rect 4282 1338 4286 1341
rect 4394 1338 4518 1341
rect 4526 1341 4529 1348
rect 4526 1338 4662 1341
rect 4666 1338 4702 1341
rect 4810 1338 4830 1341
rect 4954 1338 4998 1341
rect 5026 1338 5054 1341
rect 354 1328 422 1331
rect 530 1328 574 1331
rect 782 1331 785 1338
rect 778 1328 785 1331
rect 802 1328 806 1331
rect 866 1328 878 1331
rect 914 1328 998 1331
rect 1270 1331 1273 1338
rect 1390 1332 1393 1338
rect 2270 1332 2273 1338
rect 2534 1332 2537 1338
rect 3974 1332 3977 1338
rect 4054 1332 4057 1338
rect 1270 1328 1334 1331
rect 1550 1328 1646 1331
rect 1738 1328 1830 1331
rect 1898 1328 1942 1331
rect 2090 1328 2142 1331
rect 2162 1328 2270 1331
rect 2394 1328 2454 1331
rect 2458 1328 2510 1331
rect 2554 1328 2566 1331
rect 2874 1328 2910 1331
rect 2930 1328 2934 1331
rect 3138 1328 3142 1331
rect 3194 1328 3225 1331
rect 3250 1328 3414 1331
rect 3442 1328 3614 1331
rect 3650 1328 3734 1331
rect 3882 1328 3950 1331
rect 4170 1328 4470 1331
rect 4490 1328 4510 1331
rect 4514 1328 4886 1331
rect 4890 1328 5014 1331
rect 5042 1328 5062 1331
rect 462 1322 465 1328
rect 66 1318 190 1321
rect 194 1318 254 1321
rect 282 1318 366 1321
rect 594 1318 598 1321
rect 834 1318 950 1321
rect 954 1318 1166 1321
rect 1254 1321 1257 1328
rect 1550 1322 1553 1328
rect 1170 1318 1257 1321
rect 1322 1318 1542 1321
rect 1594 1318 1702 1321
rect 1850 1318 2198 1321
rect 2218 1318 2246 1321
rect 2326 1321 2329 1328
rect 2326 1318 2862 1321
rect 2874 1318 2878 1321
rect 3110 1321 3113 1328
rect 3026 1318 3113 1321
rect 3222 1322 3225 1328
rect 4070 1322 4073 1328
rect 3250 1318 3254 1321
rect 3290 1318 3294 1321
rect 3714 1318 3862 1321
rect 4002 1318 4014 1321
rect 4274 1318 4302 1321
rect 4338 1318 4462 1321
rect 4586 1318 4606 1321
rect 4706 1318 4790 1321
rect 282 1308 358 1311
rect 466 1308 934 1311
rect 1122 1308 1174 1311
rect 1194 1308 1222 1311
rect 1242 1308 1286 1311
rect 1290 1308 1334 1311
rect 1346 1308 1742 1311
rect 2098 1308 2214 1311
rect 2402 1308 2702 1311
rect 2842 1308 2950 1311
rect 3202 1308 3222 1311
rect 3234 1308 3238 1311
rect 3882 1308 4022 1311
rect 4258 1308 4422 1311
rect 4602 1308 4734 1311
rect 4874 1308 4894 1311
rect 4898 1308 4982 1311
rect 1048 1303 1050 1307
rect 1054 1303 1057 1307
rect 1062 1303 1064 1307
rect 2072 1303 2074 1307
rect 2078 1303 2081 1307
rect 2086 1303 2088 1307
rect 3096 1303 3098 1307
rect 3102 1303 3105 1307
rect 3110 1303 3112 1307
rect 4112 1303 4114 1307
rect 4118 1303 4121 1307
rect 4126 1303 4128 1307
rect 338 1298 374 1301
rect 514 1298 662 1301
rect 730 1298 782 1301
rect 930 1298 1038 1301
rect 1210 1298 1294 1301
rect 1298 1298 1334 1301
rect 1434 1298 1550 1301
rect 1618 1298 1950 1301
rect 2130 1298 2150 1301
rect 2186 1298 2422 1301
rect 2522 1298 2646 1301
rect 2754 1298 2854 1301
rect 2874 1298 2998 1301
rect 3154 1298 3214 1301
rect 3394 1298 3422 1301
rect 3522 1298 3550 1301
rect 3618 1298 3686 1301
rect 3706 1298 3918 1301
rect 3946 1298 4046 1301
rect 4266 1298 4278 1301
rect 4282 1298 4302 1301
rect 4314 1298 4438 1301
rect 4682 1298 4710 1301
rect 4786 1298 5014 1301
rect 3246 1292 3249 1298
rect 3446 1292 3449 1298
rect 106 1288 134 1291
rect 138 1288 166 1291
rect 190 1288 198 1291
rect 202 1288 334 1291
rect 370 1288 486 1291
rect 578 1288 678 1291
rect 706 1288 750 1291
rect 1058 1288 1126 1291
rect 1226 1288 1310 1291
rect 1326 1288 1342 1291
rect 1490 1288 1574 1291
rect 1602 1288 1630 1291
rect 1714 1288 1726 1291
rect 1858 1288 1910 1291
rect 1946 1288 2022 1291
rect 2026 1288 2046 1291
rect 2058 1288 2094 1291
rect 2210 1288 2230 1291
rect 2290 1288 2462 1291
rect 2594 1288 2686 1291
rect 2706 1288 2929 1291
rect 2986 1288 3126 1291
rect 3154 1288 3230 1291
rect 3362 1288 3382 1291
rect 3434 1288 3438 1291
rect 3458 1288 3798 1291
rect 3810 1288 3838 1291
rect 4010 1288 4086 1291
rect 4170 1288 4206 1291
rect 4226 1288 4246 1291
rect 4298 1288 4361 1291
rect 4378 1288 4390 1291
rect 4486 1291 4489 1298
rect 4474 1288 4489 1291
rect 5090 1288 5174 1291
rect 358 1282 361 1288
rect 186 1278 302 1281
rect 450 1278 550 1281
rect 642 1278 710 1281
rect 794 1278 854 1281
rect 894 1281 897 1288
rect 1326 1282 1329 1288
rect 2926 1282 2929 1288
rect 894 1278 966 1281
rect 970 1278 1142 1281
rect 1458 1278 1465 1281
rect 1474 1278 1582 1281
rect 1690 1278 1726 1281
rect 1730 1278 1750 1281
rect 1754 1278 1926 1281
rect 1946 1278 1998 1281
rect 2002 1278 2534 1281
rect 2746 1278 2902 1281
rect 2930 1278 3166 1281
rect 3186 1278 3262 1281
rect 3402 1278 3414 1281
rect 3418 1278 3470 1281
rect 3614 1278 3822 1281
rect 3826 1278 3830 1281
rect 3850 1278 3878 1281
rect 3898 1278 3902 1281
rect 3974 1281 3977 1288
rect 4358 1282 4361 1288
rect 4702 1282 4705 1288
rect 3906 1278 3977 1281
rect 4074 1278 4142 1281
rect 4146 1278 4238 1281
rect 4242 1278 4326 1281
rect 4602 1278 4702 1281
rect 4754 1278 4766 1281
rect 4770 1278 4774 1281
rect 4978 1278 5102 1281
rect 5170 1278 5182 1281
rect 590 1272 593 1278
rect 226 1268 230 1271
rect 450 1268 454 1271
rect 650 1268 670 1271
rect 854 1271 857 1278
rect 1198 1272 1201 1278
rect 1382 1272 1385 1278
rect 826 1268 857 1271
rect 994 1268 1006 1271
rect 1082 1268 1086 1271
rect 1090 1268 1094 1271
rect 1130 1268 1166 1271
rect 1330 1268 1342 1271
rect 1546 1268 1606 1271
rect 1930 1268 1950 1271
rect 1954 1268 1974 1271
rect 2026 1268 2030 1271
rect 2082 1268 2249 1271
rect 2282 1268 2294 1271
rect 2298 1268 2310 1271
rect 2630 1271 2633 1278
rect 2578 1268 2633 1271
rect 2794 1268 2846 1271
rect 2850 1268 2878 1271
rect 2954 1268 2958 1271
rect 2986 1268 3094 1271
rect 3154 1268 3158 1271
rect 3218 1268 3222 1271
rect 3226 1268 3254 1271
rect 3338 1268 3358 1271
rect 3614 1271 3617 1278
rect 4582 1272 4585 1278
rect 3410 1268 3617 1271
rect 3622 1268 3678 1271
rect 3682 1268 3694 1271
rect 3738 1268 3742 1271
rect 3818 1268 3822 1271
rect 3906 1268 4406 1271
rect 4666 1268 4718 1271
rect 4878 1271 4881 1278
rect 4878 1268 4934 1271
rect 5058 1268 5062 1271
rect 102 1262 105 1268
rect 470 1262 473 1268
rect 1110 1262 1113 1268
rect 1214 1262 1217 1268
rect 354 1258 358 1261
rect 386 1258 390 1261
rect 490 1258 646 1261
rect 658 1258 702 1261
rect 706 1258 710 1261
rect 842 1258 846 1261
rect 874 1258 982 1261
rect 986 1258 1006 1261
rect 1130 1258 1142 1261
rect 1186 1258 1201 1261
rect 1222 1261 1225 1268
rect 1262 1261 1265 1268
rect 1222 1258 1265 1261
rect 1358 1262 1361 1268
rect 1398 1262 1401 1268
rect 1662 1262 1665 1268
rect 1410 1258 1470 1261
rect 1602 1258 1606 1261
rect 1634 1258 1638 1261
rect 1706 1258 1782 1261
rect 1854 1261 1857 1268
rect 1818 1258 1857 1261
rect 1982 1262 1985 1268
rect 2246 1262 2249 1268
rect 3622 1262 3625 1268
rect 5030 1262 5033 1268
rect 2090 1258 2094 1261
rect 2162 1258 2166 1261
rect 2274 1258 2358 1261
rect 2426 1258 2430 1261
rect 2650 1258 2806 1261
rect 2882 1258 2894 1261
rect 2898 1258 2926 1261
rect 2974 1258 2982 1261
rect 2986 1258 3025 1261
rect 3042 1258 3254 1261
rect 3418 1258 3446 1261
rect 3562 1258 3598 1261
rect 3642 1258 4046 1261
rect 4242 1258 4265 1261
rect 4354 1258 4358 1261
rect 4362 1258 4366 1261
rect 4378 1258 4382 1261
rect 4506 1258 4534 1261
rect 4570 1258 4574 1261
rect 4682 1258 4686 1261
rect 4778 1258 4814 1261
rect 4818 1258 4990 1261
rect 4994 1258 5006 1261
rect 5042 1258 5078 1261
rect 1198 1252 1201 1258
rect 2414 1252 2417 1258
rect 3022 1252 3025 1258
rect 4262 1252 4265 1258
rect 5014 1252 5017 1258
rect 42 1248 113 1251
rect 234 1248 238 1251
rect 338 1248 446 1251
rect 538 1248 686 1251
rect 690 1248 758 1251
rect 794 1248 833 1251
rect 110 1242 113 1248
rect 830 1242 833 1248
rect 1110 1248 1137 1251
rect 1218 1248 1278 1251
rect 1386 1248 1414 1251
rect 1426 1248 1678 1251
rect 2066 1248 2094 1251
rect 2274 1248 2302 1251
rect 2578 1248 2582 1251
rect 2618 1248 2750 1251
rect 2962 1248 2990 1251
rect 3154 1248 3158 1251
rect 3186 1248 3190 1251
rect 3234 1248 3238 1251
rect 3298 1248 3454 1251
rect 3482 1248 3593 1251
rect 1110 1242 1113 1248
rect 1134 1242 1137 1248
rect 2142 1242 2145 1248
rect 2206 1242 2209 1248
rect 218 1238 238 1241
rect 394 1238 409 1241
rect 1242 1238 1262 1241
rect 1402 1238 1406 1241
rect 1426 1238 1438 1241
rect 1498 1238 1766 1241
rect 2050 1238 2078 1241
rect 2450 1238 2654 1241
rect 2714 1238 2838 1241
rect 3162 1238 3166 1241
rect 3206 1241 3209 1248
rect 3590 1242 3593 1248
rect 3606 1248 3646 1251
rect 3722 1248 3726 1251
rect 3794 1248 3798 1251
rect 3826 1248 3830 1251
rect 3842 1248 3846 1251
rect 3850 1248 4254 1251
rect 4418 1248 4446 1251
rect 4450 1248 4590 1251
rect 4594 1248 4622 1251
rect 4706 1248 4718 1251
rect 5062 1248 5118 1251
rect 3606 1242 3609 1248
rect 3206 1238 3302 1241
rect 3378 1238 3526 1241
rect 3562 1238 3582 1241
rect 3634 1238 3646 1241
rect 3686 1241 3689 1248
rect 4350 1242 4353 1248
rect 4750 1242 4753 1248
rect 3658 1238 3689 1241
rect 3726 1238 3750 1241
rect 3778 1238 3790 1241
rect 3874 1238 3878 1241
rect 3890 1238 4105 1241
rect 4114 1238 4262 1241
rect 4442 1238 4662 1241
rect 4790 1241 4793 1248
rect 5062 1242 5065 1248
rect 4790 1238 4806 1241
rect 406 1232 409 1238
rect 3726 1232 3729 1238
rect 506 1228 830 1231
rect 1770 1228 2110 1231
rect 2218 1228 2606 1231
rect 2610 1228 3054 1231
rect 3058 1228 3158 1231
rect 3362 1228 3574 1231
rect 3690 1228 3702 1231
rect 3754 1228 4094 1231
rect 4102 1231 4105 1238
rect 5054 1232 5057 1238
rect 4102 1228 4126 1231
rect 4322 1228 4342 1231
rect 4346 1228 4710 1231
rect 4730 1228 4790 1231
rect 4794 1228 4838 1231
rect 166 1222 169 1228
rect 458 1218 838 1221
rect 1098 1218 1206 1221
rect 1210 1218 1310 1221
rect 1738 1218 1758 1221
rect 1978 1218 2006 1221
rect 2106 1218 2198 1221
rect 2202 1218 2254 1221
rect 2258 1218 2390 1221
rect 2570 1218 2662 1221
rect 2714 1218 3350 1221
rect 3370 1218 3398 1221
rect 3402 1218 3526 1221
rect 3674 1218 3990 1221
rect 4090 1218 4246 1221
rect 4426 1218 4854 1221
rect 4858 1218 4950 1221
rect 398 1212 401 1218
rect 170 1208 374 1211
rect 562 1208 630 1211
rect 690 1208 878 1211
rect 1010 1208 1294 1211
rect 1378 1208 1454 1211
rect 1642 1208 1926 1211
rect 1930 1208 2038 1211
rect 2058 1208 2102 1211
rect 2130 1208 2262 1211
rect 2266 1208 2294 1211
rect 2298 1208 2414 1211
rect 2546 1208 2550 1211
rect 2626 1208 2766 1211
rect 2914 1208 3150 1211
rect 3182 1208 3302 1211
rect 3330 1208 3462 1211
rect 3714 1208 3966 1211
rect 4002 1208 4038 1211
rect 4042 1208 4462 1211
rect 536 1203 538 1207
rect 542 1203 545 1207
rect 550 1203 552 1207
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1574 1203 1576 1207
rect 2584 1203 2586 1207
rect 2590 1203 2593 1207
rect 2598 1203 2600 1207
rect 882 1198 902 1201
rect 978 1198 1182 1201
rect 1346 1198 1494 1201
rect 1842 1198 1894 1201
rect 2122 1198 2238 1201
rect 2642 1198 2798 1201
rect 3182 1201 3185 1208
rect 3608 1203 3610 1207
rect 3614 1203 3617 1207
rect 3622 1203 3624 1207
rect 4632 1203 4634 1207
rect 4638 1203 4641 1207
rect 4646 1203 4648 1207
rect 3106 1198 3185 1201
rect 3290 1198 3358 1201
rect 3442 1198 3454 1201
rect 3498 1198 3558 1201
rect 3722 1198 3734 1201
rect 3922 1198 3942 1201
rect 3954 1198 4382 1201
rect 378 1188 390 1191
rect 434 1188 438 1191
rect 1194 1188 1390 1191
rect 1522 1188 1598 1191
rect 1602 1188 1902 1191
rect 1906 1188 2030 1191
rect 2194 1188 2614 1191
rect 2626 1188 3150 1191
rect 3154 1188 3214 1191
rect 3282 1188 3294 1191
rect 3314 1188 4086 1191
rect 4098 1188 4230 1191
rect 4258 1188 4366 1191
rect 4466 1188 4518 1191
rect 4554 1188 4742 1191
rect 202 1178 382 1181
rect 386 1178 718 1181
rect 722 1178 1470 1181
rect 1474 1178 1510 1181
rect 1514 1178 1838 1181
rect 2018 1178 2182 1181
rect 2458 1178 3022 1181
rect 3290 1178 3326 1181
rect 3466 1178 3702 1181
rect 4002 1178 4070 1181
rect 4146 1178 4198 1181
rect 4314 1178 4646 1181
rect 682 1168 750 1171
rect 762 1168 790 1171
rect 874 1168 926 1171
rect 1078 1168 1526 1171
rect 1534 1168 1582 1171
rect 1754 1168 1814 1171
rect 1834 1168 1878 1171
rect 1882 1168 1926 1171
rect 2298 1168 2374 1171
rect 2634 1168 2638 1171
rect 2658 1168 2726 1171
rect 2898 1168 2998 1171
rect 3290 1168 3310 1171
rect 3762 1168 3854 1171
rect 3906 1168 3910 1171
rect 4146 1168 4158 1171
rect 4346 1168 4470 1171
rect 4602 1168 4806 1171
rect 190 1161 193 1168
rect 206 1161 209 1168
rect 190 1158 209 1161
rect 218 1158 222 1161
rect 590 1161 593 1168
rect 1078 1162 1081 1168
rect 1534 1162 1537 1168
rect 586 1158 593 1161
rect 730 1158 766 1161
rect 770 1158 790 1161
rect 938 1158 1078 1161
rect 1154 1158 1174 1161
rect 1178 1158 1414 1161
rect 1426 1158 1446 1161
rect 1458 1158 1486 1161
rect 1522 1158 1534 1161
rect 1558 1158 1566 1161
rect 1570 1158 1646 1161
rect 1810 1158 2014 1161
rect 2050 1158 2054 1161
rect 2118 1161 2121 1168
rect 2114 1158 2121 1161
rect 2178 1158 2318 1161
rect 2406 1161 2409 1168
rect 2422 1161 2425 1168
rect 2406 1158 2425 1161
rect 2462 1161 2465 1168
rect 2450 1158 2465 1161
rect 2474 1158 2678 1161
rect 2698 1158 2766 1161
rect 2786 1158 2846 1161
rect 2906 1158 2998 1161
rect 3178 1158 3230 1161
rect 3502 1161 3505 1168
rect 3870 1162 3873 1168
rect 4174 1162 4177 1168
rect 3466 1158 3505 1161
rect 3746 1158 3766 1161
rect 3922 1158 3982 1161
rect 4026 1158 4046 1161
rect 4050 1158 4054 1161
rect 4106 1158 4150 1161
rect 4214 1161 4217 1168
rect 4342 1162 4345 1168
rect 4214 1158 4302 1161
rect 4354 1158 4358 1161
rect 4482 1158 4486 1161
rect 4506 1158 4510 1161
rect 4522 1158 4526 1161
rect 4530 1158 4566 1161
rect 4634 1158 4670 1161
rect 4674 1158 4710 1161
rect 110 1151 113 1158
rect 470 1152 473 1158
rect 110 1148 134 1151
rect 154 1148 182 1151
rect 186 1148 246 1151
rect 562 1148 566 1151
rect 586 1148 598 1151
rect 618 1148 670 1151
rect 746 1148 782 1151
rect 834 1148 838 1151
rect 898 1148 902 1151
rect 946 1148 958 1151
rect 1018 1148 1022 1151
rect 1050 1148 1054 1151
rect 1130 1148 1158 1151
rect 1242 1148 1246 1151
rect 1346 1148 1382 1151
rect 1386 1148 1430 1151
rect 1442 1148 1454 1151
rect 1498 1148 1502 1151
rect 1562 1148 1566 1151
rect 1706 1148 1710 1151
rect 1794 1148 1854 1151
rect 1938 1148 2254 1151
rect 2258 1148 2262 1151
rect 2342 1151 2345 1158
rect 2342 1148 2430 1151
rect 2694 1151 2697 1158
rect 2530 1148 2697 1151
rect 2706 1148 2710 1151
rect 2778 1148 2841 1151
rect 2866 1148 2926 1151
rect 2946 1148 3022 1151
rect 734 1142 737 1148
rect 2838 1142 2841 1148
rect 3114 1148 3270 1151
rect 3302 1148 3318 1151
rect 3338 1148 3342 1151
rect 3378 1148 3382 1151
rect 3514 1148 3518 1151
rect 3542 1151 3545 1158
rect 3638 1152 3641 1158
rect 3530 1148 3545 1151
rect 3578 1148 3598 1151
rect 3682 1148 3742 1151
rect 3798 1151 3801 1158
rect 3786 1148 3801 1151
rect 3822 1151 3825 1158
rect 3810 1148 3825 1151
rect 3830 1152 3833 1158
rect 3862 1151 3865 1158
rect 4102 1152 4105 1158
rect 3862 1148 3894 1151
rect 3906 1148 3934 1151
rect 4106 1148 4206 1151
rect 4210 1148 4390 1151
rect 4394 1148 4414 1151
rect 4426 1148 4438 1151
rect 4466 1148 4470 1151
rect 4474 1148 4478 1151
rect 4506 1148 4526 1151
rect 4546 1148 4582 1151
rect 4634 1148 4638 1151
rect 4698 1148 4702 1151
rect 4858 1148 4878 1151
rect 4890 1148 4918 1151
rect 4938 1148 4966 1151
rect 5002 1148 5078 1151
rect 3302 1142 3305 1148
rect 4662 1142 4665 1148
rect 18 1138 294 1141
rect 298 1138 502 1141
rect 562 1138 662 1141
rect 666 1138 734 1141
rect 810 1138 822 1141
rect 994 1138 998 1141
rect 1170 1138 1174 1141
rect 1298 1138 1478 1141
rect 1506 1138 1558 1141
rect 1562 1138 1614 1141
rect 1682 1138 1689 1141
rect 1722 1138 1726 1141
rect 1786 1138 1982 1141
rect 2002 1138 2014 1141
rect 2066 1138 2070 1141
rect 2106 1138 2190 1141
rect 2202 1138 2278 1141
rect 2282 1138 2406 1141
rect 2642 1138 2678 1141
rect 2770 1138 2782 1141
rect 2922 1138 2958 1141
rect 2962 1138 2966 1141
rect 3130 1138 3214 1141
rect 3218 1138 3294 1141
rect 3314 1138 4054 1141
rect 4074 1138 4166 1141
rect 4378 1138 4382 1141
rect 4482 1138 4486 1141
rect 4490 1138 4598 1141
rect 4698 1138 4798 1141
rect 4866 1138 4886 1141
rect 4906 1138 4926 1141
rect 4986 1138 5006 1141
rect 66 1128 86 1131
rect 274 1128 366 1131
rect 370 1128 462 1131
rect 510 1131 513 1138
rect 510 1128 614 1131
rect 634 1128 654 1131
rect 746 1128 750 1131
rect 770 1128 886 1131
rect 942 1131 945 1138
rect 1078 1132 1081 1138
rect 1686 1132 1689 1138
rect 942 1128 1054 1131
rect 1154 1128 1182 1131
rect 1258 1128 1294 1131
rect 1354 1128 1406 1131
rect 1410 1128 1446 1131
rect 1466 1128 1518 1131
rect 1862 1128 1870 1131
rect 1874 1128 1990 1131
rect 2038 1131 2041 1138
rect 2046 1131 2049 1138
rect 2702 1132 2705 1138
rect 2942 1132 2945 1138
rect 2038 1128 2049 1131
rect 2194 1128 2342 1131
rect 2406 1128 2526 1131
rect 2982 1131 2985 1138
rect 3046 1131 3049 1138
rect 2982 1128 3049 1131
rect 3210 1128 3230 1131
rect 3326 1128 3494 1131
rect 3518 1128 3782 1131
rect 3866 1128 3878 1131
rect 3890 1128 3902 1131
rect 3938 1128 3942 1131
rect 4098 1128 4110 1131
rect 4290 1128 4414 1131
rect 4422 1131 4425 1138
rect 4422 1128 4550 1131
rect 4778 1128 4950 1131
rect 4954 1128 5014 1131
rect 246 1122 249 1128
rect 362 1118 502 1121
rect 586 1118 902 1121
rect 910 1121 913 1128
rect 2406 1122 2409 1128
rect 2606 1122 2609 1128
rect 906 1118 913 1121
rect 1382 1118 1390 1121
rect 1394 1118 1414 1121
rect 1706 1118 1798 1121
rect 1802 1118 1838 1121
rect 1842 1118 2302 1121
rect 2690 1118 2750 1121
rect 2806 1121 2809 1128
rect 3326 1122 3329 1128
rect 3518 1122 3521 1128
rect 2754 1118 2809 1121
rect 2986 1118 3174 1121
rect 3226 1118 3254 1121
rect 3562 1118 3670 1121
rect 3682 1118 3710 1121
rect 3746 1118 3750 1121
rect 3818 1118 3886 1121
rect 4050 1118 4054 1121
rect 4410 1118 4526 1121
rect 4874 1118 4894 1121
rect 4922 1118 4926 1121
rect 402 1108 790 1111
rect 794 1108 798 1111
rect 810 1108 846 1111
rect 874 1108 958 1111
rect 1154 1108 1758 1111
rect 1810 1108 1910 1111
rect 1978 1108 1990 1111
rect 2250 1108 2270 1111
rect 2290 1108 2470 1111
rect 2626 1108 2654 1111
rect 2666 1108 2878 1111
rect 3130 1108 3358 1111
rect 3402 1108 3422 1111
rect 3426 1108 3686 1111
rect 3714 1108 3838 1111
rect 4522 1108 4726 1111
rect 1048 1103 1050 1107
rect 1054 1103 1057 1107
rect 1062 1103 1064 1107
rect 2072 1103 2074 1107
rect 2078 1103 2081 1107
rect 2086 1103 2088 1107
rect 3096 1103 3098 1107
rect 3102 1103 3105 1107
rect 3110 1103 3112 1107
rect 3694 1102 3697 1108
rect 4112 1103 4114 1107
rect 4118 1103 4121 1107
rect 4126 1103 4128 1107
rect 578 1098 614 1101
rect 842 1098 990 1101
rect 1098 1098 1174 1101
rect 1378 1098 1406 1101
rect 1658 1098 1662 1101
rect 1674 1098 1718 1101
rect 1738 1098 2049 1101
rect 2114 1098 2118 1101
rect 2122 1098 2182 1101
rect 2242 1098 2246 1101
rect 2306 1098 2406 1101
rect 2578 1098 2734 1101
rect 2738 1098 2934 1101
rect 3178 1098 3238 1101
rect 3266 1098 3462 1101
rect 3594 1098 3598 1101
rect 4402 1098 4830 1101
rect 742 1092 745 1098
rect 2046 1092 2049 1098
rect 410 1088 478 1091
rect 482 1088 486 1091
rect 1010 1088 1102 1091
rect 1402 1088 1478 1091
rect 1482 1088 1566 1091
rect 1658 1088 1734 1091
rect 1874 1088 1878 1091
rect 1898 1088 2006 1091
rect 2050 1088 2206 1091
rect 2274 1088 2390 1091
rect 2658 1088 2702 1091
rect 2738 1088 2862 1091
rect 2990 1088 2998 1091
rect 3002 1088 3206 1091
rect 3370 1088 3478 1091
rect 3482 1088 3502 1091
rect 3530 1088 3614 1091
rect 3666 1088 3670 1091
rect 3726 1088 3734 1091
rect 3738 1088 3774 1091
rect 3874 1088 4390 1091
rect 4866 1088 4878 1091
rect 4946 1088 5054 1091
rect 214 1081 217 1088
rect 42 1078 217 1081
rect 330 1078 342 1081
rect 346 1078 590 1081
rect 594 1078 686 1081
rect 806 1081 809 1088
rect 714 1078 809 1081
rect 858 1078 862 1081
rect 1074 1078 1078 1081
rect 1082 1078 1134 1081
rect 1498 1078 1638 1081
rect 1830 1081 1833 1088
rect 1770 1078 1833 1081
rect 1842 1078 1902 1081
rect 1962 1078 1966 1081
rect 1970 1078 2022 1081
rect 2026 1078 2102 1081
rect 2234 1078 2382 1081
rect 2554 1078 2774 1081
rect 2938 1078 3006 1081
rect 3074 1078 3134 1081
rect 3186 1078 3262 1081
rect 3298 1078 3382 1081
rect 3458 1078 3550 1081
rect 3554 1078 3614 1081
rect 3658 1078 3662 1081
rect 3666 1078 3742 1081
rect 3770 1078 4014 1081
rect 4018 1078 4030 1081
rect 4178 1078 4310 1081
rect 4594 1078 4630 1081
rect 4634 1078 4662 1081
rect 4810 1078 4862 1081
rect 114 1068 134 1071
rect 174 1068 182 1071
rect 186 1068 222 1071
rect 234 1068 342 1071
rect 354 1068 414 1071
rect 426 1068 462 1071
rect 714 1068 790 1071
rect 794 1068 806 1071
rect 866 1068 870 1071
rect 890 1068 894 1071
rect 1034 1068 1070 1071
rect 1090 1068 1094 1071
rect 1106 1068 1190 1071
rect 1450 1068 1454 1071
rect 1538 1068 1614 1071
rect 1646 1071 1649 1078
rect 1626 1068 1649 1071
rect 1690 1068 1710 1071
rect 1778 1068 1814 1071
rect 1818 1068 1846 1071
rect 1882 1068 1886 1071
rect 1898 1068 1902 1071
rect 1922 1068 2078 1071
rect 2082 1068 2150 1071
rect 2234 1068 2238 1071
rect 2258 1068 2438 1071
rect 2546 1068 2590 1071
rect 2674 1068 2678 1071
rect 2722 1068 2726 1071
rect 2830 1071 2833 1078
rect 2762 1068 2862 1071
rect 2930 1068 3006 1071
rect 3010 1068 3038 1071
rect 3082 1068 3182 1071
rect 3186 1068 3334 1071
rect 3338 1068 3342 1071
rect 3354 1068 3414 1071
rect 3434 1068 3462 1071
rect 3482 1068 3486 1071
rect 3506 1068 3838 1071
rect 3930 1068 3934 1071
rect 4042 1068 4062 1071
rect 4098 1068 4206 1071
rect 4326 1071 4329 1078
rect 4230 1068 4358 1071
rect 4454 1071 4457 1078
rect 4454 1068 4526 1071
rect 4566 1071 4569 1078
rect 4554 1068 4569 1071
rect 4906 1068 4942 1071
rect 4966 1071 4969 1078
rect 4966 1068 5046 1071
rect 102 1061 105 1068
rect 1910 1062 1913 1068
rect 50 1058 105 1061
rect 130 1058 238 1061
rect 338 1058 398 1061
rect 402 1058 422 1061
rect 738 1058 918 1061
rect 930 1058 934 1061
rect 954 1058 958 1061
rect 1050 1058 1054 1061
rect 1066 1058 1190 1061
rect 1250 1058 1278 1061
rect 1314 1058 1614 1061
rect 1658 1058 1662 1061
rect 2018 1058 2022 1061
rect 2098 1058 2118 1061
rect 2210 1058 2246 1061
rect 2266 1058 2270 1061
rect 2290 1058 2337 1061
rect 2506 1058 2510 1061
rect 2622 1061 2625 1068
rect 2594 1058 2625 1061
rect 2662 1061 2665 1068
rect 2662 1058 2686 1061
rect 2730 1058 2782 1061
rect 2858 1058 2934 1061
rect 3042 1058 3118 1061
rect 3122 1058 3142 1061
rect 3266 1058 3310 1061
rect 3314 1058 3590 1061
rect 3618 1058 3646 1061
rect 3706 1058 3734 1061
rect 3738 1058 3742 1061
rect 3762 1058 3854 1061
rect 3874 1058 3958 1061
rect 4050 1058 4134 1061
rect 4230 1061 4233 1068
rect 4422 1061 4425 1068
rect 4758 1062 4761 1068
rect 4814 1062 4817 1068
rect 4218 1058 4233 1061
rect 4342 1058 4425 1061
rect 4434 1058 4510 1061
rect 4530 1058 4574 1061
rect 4602 1058 4630 1061
rect 4634 1058 4710 1061
rect 4714 1058 4753 1061
rect 4858 1058 4990 1061
rect 5010 1058 5030 1061
rect 98 1048 166 1051
rect 170 1048 182 1051
rect 202 1048 374 1051
rect 430 1051 433 1058
rect 2334 1052 2337 1058
rect 2630 1052 2633 1058
rect 2694 1052 2697 1058
rect 3078 1052 3081 1058
rect 4342 1052 4345 1058
rect 430 1048 534 1051
rect 554 1048 998 1051
rect 1162 1048 1286 1051
rect 1290 1048 1302 1051
rect 1354 1048 1422 1051
rect 1442 1048 1558 1051
rect 1598 1048 1617 1051
rect 198 1038 214 1041
rect 282 1038 353 1041
rect 382 1041 385 1048
rect 1134 1042 1137 1048
rect 370 1038 385 1041
rect 418 1038 558 1041
rect 810 1038 830 1041
rect 898 1038 902 1041
rect 1142 1041 1145 1048
rect 1598 1042 1601 1048
rect 1614 1042 1617 1048
rect 1814 1048 1822 1051
rect 1906 1048 1926 1051
rect 2030 1048 2086 1051
rect 2110 1048 2150 1051
rect 2162 1048 2214 1051
rect 2254 1048 2281 1051
rect 2386 1048 2406 1051
rect 2430 1048 2449 1051
rect 2466 1048 2502 1051
rect 2570 1048 2614 1051
rect 2842 1048 2926 1051
rect 2946 1048 2966 1051
rect 3186 1048 3278 1051
rect 3442 1048 3446 1051
rect 3466 1048 3606 1051
rect 3610 1048 3766 1051
rect 3786 1048 3990 1051
rect 4058 1048 4062 1051
rect 4614 1048 4718 1051
rect 4750 1051 4753 1058
rect 4750 1048 4878 1051
rect 4882 1048 4926 1051
rect 1142 1038 1166 1041
rect 1182 1038 1222 1041
rect 1290 1038 1294 1041
rect 1490 1038 1502 1041
rect 1798 1041 1801 1048
rect 1714 1038 1801 1041
rect 1814 1042 1817 1048
rect 2030 1042 2033 1048
rect 2110 1042 2113 1048
rect 2254 1042 2257 1048
rect 2278 1042 2281 1048
rect 2430 1042 2433 1048
rect 2446 1042 2449 1048
rect 4190 1042 4193 1048
rect 4614 1042 4617 1048
rect 2570 1038 3190 1041
rect 3194 1038 3366 1041
rect 3378 1038 3382 1041
rect 3402 1038 3558 1041
rect 3594 1038 3662 1041
rect 3666 1038 3694 1041
rect 3746 1038 3750 1041
rect 3786 1038 3918 1041
rect 4658 1038 4694 1041
rect 4714 1038 4750 1041
rect 198 1032 201 1038
rect 350 1032 353 1038
rect 1182 1032 1185 1038
rect 2222 1032 2225 1038
rect 714 1028 910 1031
rect 1122 1028 1166 1031
rect 1602 1028 1606 1031
rect 1634 1028 1854 1031
rect 1986 1028 2134 1031
rect 2146 1028 2150 1031
rect 2418 1028 2430 1031
rect 2522 1028 2678 1031
rect 2754 1028 2766 1031
rect 3114 1028 3782 1031
rect 3794 1028 4678 1031
rect 4778 1028 5126 1031
rect 5130 1028 5174 1031
rect 138 1018 446 1021
rect 874 1018 1102 1021
rect 1178 1018 1246 1021
rect 1250 1018 1406 1021
rect 1762 1018 2014 1021
rect 2562 1018 2830 1021
rect 3034 1018 3726 1021
rect 3818 1018 3822 1021
rect 4258 1018 4574 1021
rect 4578 1018 4742 1021
rect 4774 1021 4777 1028
rect 4746 1018 4777 1021
rect 218 1008 414 1011
rect 442 1008 494 1011
rect 982 1008 1326 1011
rect 1778 1008 1974 1011
rect 2010 1008 2286 1011
rect 2618 1008 3022 1011
rect 3082 1008 3390 1011
rect 3506 1008 3510 1011
rect 3514 1008 3598 1011
rect 3674 1008 3758 1011
rect 3770 1008 3950 1011
rect 3954 1008 4086 1011
rect 4202 1008 4622 1011
rect 4682 1008 4790 1011
rect 536 1003 538 1007
rect 542 1003 545 1007
rect 550 1003 552 1007
rect 266 998 390 1001
rect 394 998 518 1001
rect 634 998 646 1001
rect 982 1001 985 1008
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1574 1003 1576 1007
rect 2584 1003 2586 1007
rect 2590 1003 2593 1007
rect 2598 1003 2600 1007
rect 3608 1003 3610 1007
rect 3614 1003 3617 1007
rect 3622 1003 3624 1007
rect 4632 1003 4634 1007
rect 4638 1003 4641 1007
rect 4646 1003 4648 1007
rect 786 998 985 1001
rect 1114 998 1150 1001
rect 1658 998 2022 1001
rect 2026 998 2118 1001
rect 2210 998 2294 1001
rect 2410 998 2542 1001
rect 2546 998 2574 1001
rect 2682 998 2798 1001
rect 2802 998 2830 1001
rect 2906 998 3094 1001
rect 3098 998 3238 1001
rect 3738 998 3902 1001
rect 3994 998 4142 1001
rect 4698 998 4702 1001
rect 106 988 134 991
rect 202 988 230 991
rect 234 988 238 991
rect 322 988 374 991
rect 410 988 454 991
rect 458 988 462 991
rect 506 988 534 991
rect 538 988 678 991
rect 842 988 958 991
rect 962 988 1022 991
rect 1146 988 1422 991
rect 1426 988 1630 991
rect 1810 988 1830 991
rect 1946 988 1966 991
rect 2122 988 2486 991
rect 2490 988 2678 991
rect 3058 988 3062 991
rect 3482 988 3614 991
rect 3618 988 3654 991
rect 3922 988 3942 991
rect 4394 988 4486 991
rect 4578 988 4638 991
rect 4738 988 4798 991
rect 3990 982 3993 988
rect 162 978 414 981
rect 418 978 662 981
rect 666 978 1134 981
rect 1226 978 1318 981
rect 1402 978 1606 981
rect 1986 978 2046 981
rect 2058 978 2550 981
rect 2818 978 2966 981
rect 3122 978 3166 981
rect 3274 978 3422 981
rect 3802 978 3926 981
rect 4402 978 4425 981
rect 4458 978 4998 981
rect 5002 978 5062 981
rect 106 968 198 971
rect 274 968 406 971
rect 410 968 718 971
rect 826 968 830 971
rect 922 968 1030 971
rect 1066 968 1134 971
rect 1186 968 1214 971
rect 1218 968 1398 971
rect 1466 968 1566 971
rect 1570 968 1614 971
rect 1666 968 1806 971
rect 1810 968 1830 971
rect 1906 968 2014 971
rect 2018 968 2094 971
rect 2098 968 2454 971
rect 2458 968 2542 971
rect 2546 968 2870 971
rect 2874 968 3126 971
rect 3354 968 3470 971
rect 3946 968 3998 971
rect 4026 968 4214 971
rect 4422 971 4425 978
rect 4422 968 4542 971
rect 4786 968 4870 971
rect 206 961 209 968
rect 138 958 209 961
rect 346 958 358 961
rect 362 958 1118 961
rect 1122 958 1238 961
rect 1258 958 1366 961
rect 1450 958 1462 961
rect 1466 958 1470 961
rect 1530 958 1550 961
rect 1590 958 1598 961
rect 1602 958 1678 961
rect 1838 961 1841 968
rect 4390 962 4393 968
rect 4414 962 4417 968
rect 1834 958 1841 961
rect 2002 958 2110 961
rect 2166 958 2174 961
rect 2562 958 2566 961
rect 2578 958 2758 961
rect 2826 958 2926 961
rect 3026 958 3126 961
rect 3146 958 3174 961
rect 3258 958 3302 961
rect 3306 958 3326 961
rect 3362 958 3398 961
rect 3418 958 3422 961
rect 3498 958 3550 961
rect 3770 958 3830 961
rect 3922 958 3974 961
rect 4038 958 4094 961
rect 4330 958 4342 961
rect 4418 958 4718 961
rect 4758 961 4761 968
rect 4758 958 4814 961
rect 4890 958 4894 961
rect 4914 958 5030 961
rect 1774 952 1777 958
rect 370 948 374 951
rect 474 948 494 951
rect 614 948 646 951
rect 658 948 670 951
rect 706 948 798 951
rect 802 948 814 951
rect 818 948 830 951
rect 854 948 905 951
rect 1138 948 1142 951
rect 1258 948 1302 951
rect 110 941 113 948
rect 614 942 617 948
rect 854 942 857 948
rect 902 942 905 948
rect 1174 942 1177 948
rect 1394 948 1438 951
rect 1442 948 1478 951
rect 1498 948 1502 951
rect 1506 948 1582 951
rect 1586 948 1662 951
rect 1834 948 1910 951
rect 2090 948 2190 951
rect 2226 948 2230 951
rect 2382 951 2385 958
rect 2486 952 2489 958
rect 2346 948 2385 951
rect 2466 948 2486 951
rect 2610 948 2625 951
rect 66 938 174 941
rect 346 938 446 941
rect 474 938 606 941
rect 698 938 702 941
rect 730 938 734 941
rect 818 938 822 941
rect 994 938 998 941
rect 1178 938 1198 941
rect 1354 938 1518 941
rect 1522 938 1526 941
rect 1610 938 1638 941
rect 1702 941 1705 948
rect 1702 938 1734 941
rect 1738 938 1918 941
rect 2066 938 2094 941
rect 2186 938 2198 941
rect 2326 941 2329 948
rect 2622 942 2625 948
rect 2658 948 2662 951
rect 2666 948 2782 951
rect 2874 948 2918 951
rect 2958 951 2961 958
rect 2958 948 2974 951
rect 3082 948 3118 951
rect 3210 948 3270 951
rect 3274 948 3281 951
rect 3322 948 3462 951
rect 3466 948 3526 951
rect 3530 948 3638 951
rect 3662 948 3750 951
rect 3886 951 3889 958
rect 3810 948 3889 951
rect 3974 951 3977 958
rect 3990 951 3993 958
rect 3974 948 3993 951
rect 4006 952 4009 958
rect 4038 952 4041 958
rect 4018 948 4038 951
rect 4070 948 4078 951
rect 4082 948 4158 951
rect 2646 942 2649 948
rect 3030 942 3033 948
rect 2326 938 2350 941
rect 2354 938 2454 941
rect 2530 938 2574 941
rect 2858 938 2894 941
rect 2898 938 3014 941
rect 3174 941 3177 948
rect 3662 942 3665 948
rect 3098 938 3177 941
rect 3274 938 3278 941
rect 3410 938 3414 941
rect 3554 938 3641 941
rect 3794 938 3798 941
rect 3826 938 3830 941
rect 3926 941 3929 948
rect 4282 948 4342 951
rect 4354 948 4446 951
rect 4466 948 4510 951
rect 4674 948 4678 951
rect 4714 948 4726 951
rect 4770 948 4774 951
rect 4778 948 4798 951
rect 4898 948 4902 951
rect 4930 948 4942 951
rect 5102 951 5105 958
rect 5102 948 5150 951
rect 4694 942 4697 948
rect 3922 938 3929 941
rect 3938 938 4054 941
rect 4058 938 4070 941
rect 4074 938 4198 941
rect 4218 938 4321 941
rect 262 932 265 938
rect 2214 932 2217 938
rect 3470 932 3473 938
rect 3638 932 3641 938
rect 4318 932 4321 938
rect 4386 938 4510 941
rect 4722 938 4774 941
rect 4786 938 4886 941
rect 4990 941 4993 948
rect 4990 938 5006 941
rect 5042 938 5134 941
rect 5162 938 5166 941
rect 4358 932 4361 938
rect 250 928 254 931
rect 530 928 646 931
rect 650 928 774 931
rect 842 928 1086 931
rect 1194 928 1246 931
rect 1250 928 1358 931
rect 1482 928 1486 931
rect 1530 928 1678 931
rect 1794 928 1806 931
rect 1834 928 2174 931
rect 2386 928 2390 931
rect 2442 928 2654 931
rect 2802 928 2881 931
rect 2970 928 2974 931
rect 2986 928 3110 931
rect 3138 928 3158 931
rect 3162 928 3214 931
rect 3258 928 3286 931
rect 3730 928 3774 931
rect 3810 928 3814 931
rect 3986 928 4022 931
rect 4034 928 4038 931
rect 4154 928 4278 931
rect 4438 928 4446 931
rect 4450 928 4478 931
rect 5018 928 5062 931
rect 5066 928 5126 931
rect 5146 928 5166 931
rect 5170 928 5182 931
rect 2350 922 2353 928
rect 2878 922 2881 928
rect 250 918 406 921
rect 410 918 486 921
rect 490 918 526 921
rect 570 918 614 921
rect 618 918 702 921
rect 810 918 862 921
rect 866 918 918 921
rect 994 918 1158 921
rect 1170 918 1182 921
rect 1186 918 1382 921
rect 1386 918 1398 921
rect 1402 918 1534 921
rect 1778 918 2150 921
rect 2258 918 2262 921
rect 2370 918 2438 921
rect 2442 918 2510 921
rect 2538 918 2838 921
rect 3018 918 3278 921
rect 3362 918 3934 921
rect 4194 918 4214 921
rect 4218 918 4302 921
rect 4306 918 4374 921
rect 4378 918 4526 921
rect 4826 918 5126 921
rect 1726 912 1729 918
rect 346 908 441 911
rect 602 908 670 911
rect 794 908 886 911
rect 1194 908 1198 911
rect 1218 908 1278 911
rect 1282 908 1342 911
rect 1362 908 1430 911
rect 1434 908 1598 911
rect 1778 908 1798 911
rect 1802 908 1846 911
rect 1914 908 1966 911
rect 2010 908 2022 911
rect 2130 908 2166 911
rect 2482 908 2630 911
rect 2634 908 3078 911
rect 3210 908 3782 911
rect 3954 908 4086 911
rect 4090 908 4102 911
rect 4202 908 4414 911
rect 4418 908 4438 911
rect 4474 908 4502 911
rect 4506 908 4614 911
rect 4722 908 4870 911
rect 438 902 441 908
rect 894 902 897 908
rect 1048 903 1050 907
rect 1054 903 1057 907
rect 1062 903 1064 907
rect 2072 903 2074 907
rect 2078 903 2081 907
rect 2086 903 2088 907
rect 2206 902 2209 908
rect 3096 903 3098 907
rect 3102 903 3105 907
rect 3110 903 3112 907
rect 4112 903 4114 907
rect 4118 903 4121 907
rect 4126 903 4128 907
rect 442 898 510 901
rect 562 898 878 901
rect 1210 898 1230 901
rect 1322 898 1374 901
rect 1394 898 1462 901
rect 1466 898 1526 901
rect 1538 898 1550 901
rect 1554 898 1678 901
rect 1770 898 1790 901
rect 1874 898 2022 901
rect 2314 898 2582 901
rect 2586 898 2630 901
rect 2858 898 2870 901
rect 2954 898 3030 901
rect 3122 898 3206 901
rect 3322 898 3710 901
rect 3786 898 3806 901
rect 3874 898 3950 901
rect 4306 898 4982 901
rect 422 892 425 898
rect 3246 892 3249 898
rect 106 888 134 891
rect 138 888 358 891
rect 566 888 574 891
rect 578 888 598 891
rect 606 888 838 891
rect 986 888 1206 891
rect 1234 888 1262 891
rect 1266 888 1382 891
rect 1426 888 1502 891
rect 1546 888 1566 891
rect 1570 888 1606 891
rect 1842 888 1910 891
rect 1962 888 2078 891
rect 2082 888 2086 891
rect 2106 888 2110 891
rect 2138 888 2222 891
rect 2226 888 2278 891
rect 2322 888 2406 891
rect 2466 888 2502 891
rect 2506 888 2526 891
rect 2614 888 2622 891
rect 2626 888 2638 891
rect 2650 888 2694 891
rect 2898 888 2929 891
rect 3106 888 3150 891
rect 3314 888 3470 891
rect 3506 888 3510 891
rect 3762 888 3822 891
rect 3930 888 3966 891
rect 4082 888 4126 891
rect 4250 888 4350 891
rect 4474 888 4478 891
rect 4490 888 4526 891
rect 4570 888 4726 891
rect 4730 888 4758 891
rect 210 878 214 881
rect 290 878 326 881
rect 606 881 609 888
rect 2926 882 2929 888
rect 330 878 609 881
rect 634 878 758 881
rect 762 878 798 881
rect 978 878 990 881
rect 1010 878 1102 881
rect 1130 878 1166 881
rect 1258 878 1350 881
rect 1354 878 1430 881
rect 1618 878 1638 881
rect 1642 878 1870 881
rect 1962 878 2038 881
rect 2154 878 2254 881
rect 2258 878 2366 881
rect 2442 878 2686 881
rect 2690 878 2814 881
rect 2834 878 2910 881
rect 2930 878 2966 881
rect 3178 878 3238 881
rect 3406 878 3414 881
rect 3418 878 3446 881
rect 3466 878 3486 881
rect 3690 878 3838 881
rect 3930 878 4054 881
rect 4210 878 4230 881
rect 4234 878 4246 881
rect 4314 878 4446 881
rect 4498 878 4582 881
rect 4698 878 4702 881
rect 4730 878 4862 881
rect 114 868 126 871
rect 314 868 326 871
rect 330 868 430 871
rect 722 868 814 871
rect 822 871 825 878
rect 822 868 926 871
rect 1074 868 1153 871
rect 1258 868 1302 871
rect 1454 871 1457 878
rect 1334 868 1457 871
rect 1506 868 1622 871
rect 1626 868 1638 871
rect 1706 868 1710 871
rect 1722 868 1742 871
rect 1746 868 1750 871
rect 1802 868 1806 871
rect 1818 868 1822 871
rect 1970 868 2070 871
rect 2074 868 2126 871
rect 2138 868 2142 871
rect 2602 868 2646 871
rect 2890 868 2894 871
rect 2954 868 2958 871
rect 3010 868 3190 871
rect 3194 868 3254 871
rect 3306 868 3342 871
rect 3346 868 3350 871
rect 3378 868 3382 871
rect 3450 868 3502 871
rect 3582 871 3585 878
rect 4454 872 4457 878
rect 3582 868 3670 871
rect 3738 868 3750 871
rect 3754 868 3918 871
rect 3954 868 3958 871
rect 3986 868 4022 871
rect 4562 868 4654 871
rect 4658 868 4814 871
rect 4994 868 5014 871
rect 150 861 153 868
rect 590 862 593 868
rect 606 862 609 868
rect 870 862 873 868
rect 50 858 121 861
rect 150 858 246 861
rect 250 858 286 861
rect 322 858 390 861
rect 410 858 478 861
rect 522 858 574 861
rect 642 858 697 861
rect 786 858 790 861
rect 962 858 966 861
rect 1006 861 1009 868
rect 1150 862 1153 868
rect 1334 862 1337 868
rect 1006 858 1086 861
rect 1130 858 1142 861
rect 1170 858 1198 861
rect 1242 858 1246 861
rect 1426 858 1430 861
rect 1478 861 1481 868
rect 1478 858 1574 861
rect 1706 858 1718 861
rect 1722 858 1838 861
rect 1954 858 2270 861
rect 2274 858 2302 861
rect 2306 858 2342 861
rect 2346 858 2534 861
rect 2538 858 2622 861
rect 2694 861 2697 868
rect 2634 858 2894 861
rect 3130 858 3166 861
rect 3174 858 3246 861
rect 3266 858 3270 861
rect 3290 858 3294 861
rect 3378 858 3414 861
rect 3442 858 3486 861
rect 3570 858 3614 861
rect 3682 858 3702 861
rect 3762 858 3926 861
rect 3938 858 3950 861
rect 3978 858 4030 861
rect 4130 858 4182 861
rect 4258 858 4310 861
rect 4406 861 4409 868
rect 4370 858 4409 861
rect 4554 858 4558 861
rect 4610 858 4638 861
rect 4738 858 4814 861
rect 4858 858 5134 861
rect 118 852 121 858
rect 694 852 697 858
rect 886 852 889 858
rect 178 848 198 851
rect 298 848 654 851
rect 746 848 782 851
rect 802 848 806 851
rect 914 848 1310 851
rect 1394 848 1406 851
rect 1410 848 1542 851
rect 1610 848 1614 851
rect 1642 848 1646 851
rect 1698 848 1766 851
rect 1770 848 1894 851
rect 2018 848 2022 851
rect 2138 848 2214 851
rect 2338 848 2454 851
rect 2522 848 2566 851
rect 2570 848 2606 851
rect 2618 848 2646 851
rect 2666 848 2686 851
rect 2690 848 2918 851
rect 3042 848 3134 851
rect 3174 851 3177 858
rect 3926 852 3929 858
rect 5182 852 5185 858
rect 3162 848 3177 851
rect 3242 848 3710 851
rect 3762 848 3774 851
rect 3822 848 3870 851
rect 4066 848 4190 851
rect 4378 848 4422 851
rect 4594 848 4694 851
rect 4990 848 5078 851
rect 1550 842 1553 848
rect 1598 842 1601 848
rect 354 838 374 841
rect 410 838 454 841
rect 458 838 662 841
rect 666 838 934 841
rect 962 838 1550 841
rect 1634 838 1638 841
rect 1754 838 1838 841
rect 2014 841 2017 848
rect 2054 841 2057 848
rect 3822 842 3825 848
rect 4470 842 4473 848
rect 4990 842 4993 848
rect 2014 838 2057 841
rect 2066 838 2558 841
rect 2670 838 2758 841
rect 2770 838 2982 841
rect 3122 838 3182 841
rect 3282 838 3342 841
rect 3346 838 3406 841
rect 3422 838 3558 841
rect 3682 838 3694 841
rect 3834 838 3870 841
rect 4250 838 4254 841
rect 4594 838 4662 841
rect 4666 838 4686 841
rect 4690 838 4710 841
rect 4714 838 4750 841
rect 2670 832 2673 838
rect 3422 832 3425 838
rect 138 828 454 831
rect 914 828 918 831
rect 930 828 966 831
rect 1418 828 1518 831
rect 1522 828 1662 831
rect 1666 828 1726 831
rect 1818 828 1822 831
rect 1850 828 2262 831
rect 2698 828 2702 831
rect 2786 828 2822 831
rect 2850 828 2958 831
rect 2962 828 3014 831
rect 3266 828 3326 831
rect 3442 828 3446 831
rect 3458 828 3462 831
rect 3546 828 3982 831
rect 4018 828 4486 831
rect 4626 828 4758 831
rect 4762 828 4790 831
rect 4794 828 4806 831
rect 186 818 190 821
rect 370 818 614 821
rect 806 821 809 828
rect 618 818 809 821
rect 874 818 934 821
rect 938 818 942 821
rect 1434 818 1438 821
rect 1554 818 2270 821
rect 2506 818 3110 821
rect 3130 818 3166 821
rect 3170 818 3230 821
rect 3234 818 3294 821
rect 3578 818 3734 821
rect 3802 818 3822 821
rect 3998 821 4001 828
rect 3998 818 4022 821
rect 4274 818 4294 821
rect 4294 812 4297 818
rect 226 808 438 811
rect 594 808 782 811
rect 834 808 1134 811
rect 1138 808 1334 811
rect 1394 808 1542 811
rect 1858 808 2078 811
rect 2130 808 2254 811
rect 2258 808 2326 811
rect 2346 808 2350 811
rect 2354 808 2486 811
rect 2610 808 2862 811
rect 2866 808 3542 811
rect 3634 808 3782 811
rect 3850 808 3854 811
rect 4306 808 4502 811
rect 536 803 538 807
rect 542 803 545 807
rect 550 803 552 807
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1574 803 1576 807
rect 2584 803 2586 807
rect 2590 803 2593 807
rect 2598 803 2600 807
rect 3608 803 3610 807
rect 3614 803 3617 807
rect 3622 803 3624 807
rect 4632 803 4634 807
rect 4638 803 4641 807
rect 4646 803 4648 807
rect 58 798 110 801
rect 114 798 126 801
rect 130 798 366 801
rect 570 798 694 801
rect 698 798 894 801
rect 954 798 1182 801
rect 1714 798 1862 801
rect 2130 798 2318 801
rect 2482 798 2502 801
rect 2642 798 2894 801
rect 2954 798 3286 801
rect 3290 798 3310 801
rect 3698 798 3774 801
rect 3786 798 3894 801
rect 3898 798 4518 801
rect 5122 798 5174 801
rect 242 788 598 791
rect 602 788 822 791
rect 826 788 862 791
rect 866 788 918 791
rect 930 788 1238 791
rect 1482 788 1558 791
rect 1738 788 1814 791
rect 1898 788 2070 791
rect 2098 788 2374 791
rect 2378 788 2550 791
rect 2554 788 2662 791
rect 2666 788 2678 791
rect 2970 788 3182 791
rect 3298 788 3422 791
rect 3482 788 3982 791
rect 3990 788 4302 791
rect 4378 788 4654 791
rect 4810 788 4910 791
rect 5026 788 5046 791
rect 5162 788 5174 791
rect 202 778 214 781
rect 218 778 910 781
rect 1242 778 1286 781
rect 1290 778 1294 781
rect 1578 778 1654 781
rect 1658 778 1662 781
rect 1706 778 2286 781
rect 2338 778 2710 781
rect 2946 778 3054 781
rect 3074 778 3174 781
rect 3258 778 3374 781
rect 3522 778 3766 781
rect 3990 781 3993 788
rect 3802 778 3993 781
rect 4010 778 4350 781
rect 4442 778 4926 781
rect 4930 778 4950 781
rect 4954 778 4998 781
rect 210 768 241 771
rect 466 768 510 771
rect 522 768 614 771
rect 658 768 886 771
rect 890 768 902 771
rect 970 768 1022 771
rect 1034 768 1150 771
rect 1186 768 1254 771
rect 1346 768 1358 771
rect 1434 768 1462 771
rect 1658 768 1718 771
rect 2366 768 2542 771
rect 2930 768 3038 771
rect 3362 768 3406 771
rect 3434 768 3438 771
rect 3442 768 3686 771
rect 3690 768 3910 771
rect 3946 768 4062 771
rect 4434 768 4510 771
rect 4754 768 5054 771
rect 5058 768 5062 771
rect 5066 768 5166 771
rect 238 762 241 768
rect 494 762 497 768
rect 266 758 278 761
rect 402 758 478 761
rect 586 758 630 761
rect 690 758 718 761
rect 798 758 806 761
rect 810 758 822 761
rect 842 758 878 761
rect 906 758 974 761
rect 994 758 998 761
rect 1066 758 1070 761
rect 1130 758 1246 761
rect 1274 758 1286 761
rect 1406 761 1409 768
rect 1306 758 1409 761
rect 1422 762 1425 768
rect 1462 761 1465 768
rect 2366 762 2369 768
rect 1462 758 1638 761
rect 1698 758 1758 761
rect 2130 758 2238 761
rect 2418 758 2438 761
rect 2654 761 2657 768
rect 3134 762 3137 768
rect 3174 762 3177 768
rect 2654 758 2726 761
rect 2802 758 2806 761
rect 2978 758 3022 761
rect 3050 758 3102 761
rect 3154 758 3158 761
rect 3250 758 3302 761
rect 3410 758 3470 761
rect 3834 758 3878 761
rect 4218 758 4294 761
rect 4330 758 4334 761
rect 4394 758 4398 761
rect 4522 758 4870 761
rect 114 748 134 751
rect 186 748 222 751
rect 226 748 230 751
rect 258 748 270 751
rect 482 748 702 751
rect 722 748 750 751
rect 770 748 774 751
rect 778 748 1062 751
rect 1090 748 1094 751
rect 1242 748 1254 751
rect 1378 748 1446 751
rect 1674 748 1678 751
rect 1686 751 1689 758
rect 2614 752 2617 758
rect 3822 752 3825 758
rect 3830 752 3833 758
rect 4014 752 4017 758
rect 1686 748 1694 751
rect 1706 748 1726 751
rect 1930 748 1945 751
rect 2034 748 2118 751
rect 2130 748 2169 751
rect 2194 748 2270 751
rect 2298 748 2302 751
rect 2322 748 2446 751
rect 2450 748 2518 751
rect 2626 748 2670 751
rect 2794 748 2809 751
rect 2906 748 2950 751
rect 2954 748 3006 751
rect 3210 748 3214 751
rect 3266 748 3270 751
rect 3298 748 3326 751
rect 3390 748 3518 751
rect 3686 748 3710 751
rect 3722 748 3726 751
rect 3778 748 3782 751
rect 3930 748 3934 751
rect 3962 748 4006 751
rect 4134 751 4137 758
rect 4074 748 4137 751
rect 4242 748 4254 751
rect 4306 748 4310 751
rect 4362 748 4366 751
rect 4438 751 4441 758
rect 4394 748 4441 751
rect 4522 748 4590 751
rect 4606 748 4737 751
rect 4770 748 4798 751
rect 4958 751 4961 758
rect 4810 748 4961 751
rect 5022 751 5025 758
rect 5022 748 5094 751
rect 238 742 241 748
rect 462 742 465 748
rect 590 742 593 748
rect 1358 742 1361 748
rect 98 738 150 741
rect 154 738 190 741
rect 306 738 310 741
rect 634 738 662 741
rect 666 738 990 741
rect 1050 738 1054 741
rect 1098 738 1110 741
rect 1122 738 1126 741
rect 1178 738 1262 741
rect 1330 738 1353 741
rect 1458 738 1502 741
rect 1534 741 1537 748
rect 1942 742 1945 748
rect 2166 742 2169 748
rect 2806 742 2809 748
rect 3070 742 3073 748
rect 3390 742 3393 748
rect 3686 742 3689 748
rect 3838 742 3841 748
rect 4606 742 4609 748
rect 4734 742 4737 748
rect 1506 738 1590 741
rect 1626 738 1798 741
rect 1818 738 1822 741
rect 1978 738 2153 741
rect 2242 738 2246 741
rect 2362 738 2366 741
rect 2418 738 2430 741
rect 2618 738 2622 741
rect 3186 738 3334 741
rect 3362 738 3366 741
rect 3722 738 3726 741
rect 3938 738 4574 741
rect 4578 738 4598 741
rect 4602 738 4606 741
rect 4666 738 4678 741
rect 4738 738 4766 741
rect 4790 738 4862 741
rect 4894 738 4974 741
rect 5066 738 5070 741
rect 998 732 1001 738
rect 1350 732 1353 738
rect 1406 732 1409 738
rect 2150 732 2153 738
rect 4790 732 4793 738
rect 4894 732 4897 738
rect 42 728 121 731
rect 170 728 206 731
rect 234 728 270 731
rect 594 728 598 731
rect 682 728 702 731
rect 786 728 830 731
rect 834 728 950 731
rect 1130 728 1134 731
rect 1154 728 1302 731
rect 1394 728 1398 731
rect 1450 728 1646 731
rect 1658 728 1670 731
rect 1970 728 2094 731
rect 2274 728 2302 731
rect 2394 728 2470 731
rect 2594 728 2710 731
rect 3010 728 3022 731
rect 3026 728 3118 731
rect 3154 728 3174 731
rect 3178 728 3198 731
rect 3202 728 3350 731
rect 3354 728 3430 731
rect 3938 728 3958 731
rect 3962 728 3998 731
rect 4106 728 4206 731
rect 4274 728 4278 731
rect 4354 728 4374 731
rect 4402 728 4558 731
rect 5042 728 5094 731
rect 118 722 121 728
rect 178 718 262 721
rect 266 718 702 721
rect 706 718 878 721
rect 970 718 1342 721
rect 1394 718 1494 721
rect 1498 718 1542 721
rect 1546 718 1998 721
rect 2002 718 2318 721
rect 2362 718 2398 721
rect 2410 718 2422 721
rect 2650 718 2686 721
rect 2790 721 2793 728
rect 3974 722 3977 728
rect 2690 718 2793 721
rect 2874 718 3078 721
rect 3106 718 3222 721
rect 4074 718 4190 721
rect 4378 718 4414 721
rect 4522 718 4774 721
rect 4778 718 4806 721
rect 5186 718 5190 721
rect 74 708 102 711
rect 106 708 294 711
rect 450 708 734 711
rect 770 708 862 711
rect 946 708 966 711
rect 978 708 1022 711
rect 1090 708 1166 711
rect 1170 708 1278 711
rect 1282 708 1390 711
rect 1410 708 1438 711
rect 1626 708 1638 711
rect 1642 708 1854 711
rect 1962 708 2006 711
rect 2018 708 2054 711
rect 2266 708 2302 711
rect 2378 708 2902 711
rect 3154 708 3414 711
rect 3474 708 3742 711
rect 3746 708 3814 711
rect 3890 708 3966 711
rect 4290 708 4294 711
rect 4330 708 4422 711
rect 4482 708 4502 711
rect 4698 708 4766 711
rect 5106 708 5126 711
rect 106 698 126 701
rect 130 698 174 701
rect 266 698 294 701
rect 298 698 486 701
rect 578 698 686 701
rect 698 698 758 701
rect 762 698 822 701
rect 862 701 865 708
rect 1048 703 1050 707
rect 1054 703 1057 707
rect 1062 703 1064 707
rect 2072 703 2074 707
rect 2078 703 2081 707
rect 2086 703 2088 707
rect 3096 703 3098 707
rect 3102 703 3105 707
rect 3110 703 3112 707
rect 4112 703 4114 707
rect 4118 703 4121 707
rect 4126 703 4128 707
rect 4886 702 4889 708
rect 4918 702 4921 708
rect 862 698 1022 701
rect 1346 698 1430 701
rect 1450 698 1454 701
rect 1594 698 1622 701
rect 1634 698 1638 701
rect 1762 698 1894 701
rect 1898 698 2062 701
rect 2114 698 2174 701
rect 2178 698 2318 701
rect 2338 698 2598 701
rect 2634 698 2846 701
rect 2914 698 2942 701
rect 2946 698 3086 701
rect 3482 698 3494 701
rect 3902 698 4046 701
rect 4250 698 4318 701
rect 4490 698 4558 701
rect 4594 698 4710 701
rect 4754 698 4758 701
rect 4762 698 4862 701
rect 3902 692 3905 698
rect 226 688 1078 691
rect 1082 688 1566 691
rect 1570 688 1766 691
rect 1770 688 1774 691
rect 2034 688 2126 691
rect 2178 688 2374 691
rect 2482 688 2566 691
rect 2570 688 2686 691
rect 2922 688 3062 691
rect 3146 688 3238 691
rect 3242 688 3262 691
rect 3314 688 3382 691
rect 3450 688 3502 691
rect 3506 688 3526 691
rect 3818 688 3902 691
rect 3946 688 4014 691
rect 4034 688 4054 691
rect 4066 688 4206 691
rect 4210 688 4310 691
rect 4442 688 4462 691
rect 4546 688 4782 691
rect 4906 688 4910 691
rect 210 678 214 681
rect 386 678 398 681
rect 402 678 446 681
rect 450 678 518 681
rect 634 678 766 681
rect 1042 678 1222 681
rect 1274 678 1350 681
rect 1418 678 1422 681
rect 1610 678 1974 681
rect 1990 681 1993 688
rect 1990 678 1998 681
rect 2018 678 2038 681
rect 2042 678 2086 681
rect 2130 678 2206 681
rect 2290 678 2358 681
rect 2466 678 2646 681
rect 2762 678 2822 681
rect 2826 678 2854 681
rect 3170 678 3182 681
rect 3194 678 3310 681
rect 3530 678 3798 681
rect 3858 678 4078 681
rect 4226 678 4246 681
rect 4354 678 4366 681
rect 4426 678 4454 681
rect 4570 678 4585 681
rect 4618 678 4654 681
rect 4738 678 5049 681
rect 86 671 89 678
rect 18 668 89 671
rect 254 671 257 678
rect 582 672 585 678
rect 830 672 833 678
rect 910 672 913 678
rect 982 672 985 678
rect 254 668 294 671
rect 338 668 358 671
rect 362 668 398 671
rect 498 668 529 671
rect 642 668 726 671
rect 794 668 830 671
rect 1034 668 1110 671
rect 1146 668 1174 671
rect 1462 671 1465 678
rect 2654 672 2657 678
rect 2934 672 2937 678
rect 4582 672 4585 678
rect 5046 672 5049 678
rect 1230 668 1465 671
rect 1498 668 1590 671
rect 1666 668 1670 671
rect 1690 668 1694 671
rect 1770 668 1902 671
rect 1946 668 2006 671
rect 2042 668 2134 671
rect 2186 668 2294 671
rect 2354 668 2374 671
rect 2450 668 2510 671
rect 2906 668 2910 671
rect 3010 668 3017 671
rect 3066 668 3110 671
rect 3154 668 3158 671
rect 3218 668 3286 671
rect 3290 668 3846 671
rect 3922 668 3934 671
rect 4050 668 4390 671
rect 4410 668 4430 671
rect 4626 668 4630 671
rect 4770 668 4862 671
rect 5050 668 5086 671
rect 190 661 193 668
rect 122 658 193 661
rect 214 662 217 668
rect 330 658 414 661
rect 418 658 470 661
rect 482 658 518 661
rect 526 661 529 668
rect 526 658 654 661
rect 714 658 718 661
rect 846 661 849 668
rect 1230 662 1233 668
rect 1246 662 1249 668
rect 778 658 849 661
rect 906 658 918 661
rect 970 658 1022 661
rect 1114 658 1142 661
rect 1418 658 1422 661
rect 1458 658 1502 661
rect 1546 658 1622 661
rect 1674 658 1678 661
rect 1730 658 1742 661
rect 1754 658 1758 661
rect 1762 658 1862 661
rect 1866 658 1902 661
rect 1906 658 2038 661
rect 2042 658 2366 661
rect 2386 658 2454 661
rect 2614 661 2617 668
rect 3014 662 3017 668
rect 3166 662 3169 668
rect 2614 658 2630 661
rect 2650 658 2798 661
rect 2930 658 2934 661
rect 3058 658 3078 661
rect 3082 658 3118 661
rect 3206 661 3209 668
rect 3950 662 3953 668
rect 4446 662 4449 668
rect 3202 658 3209 661
rect 3322 658 3425 661
rect 3498 658 3582 661
rect 3730 658 3750 661
rect 3754 658 3774 661
rect 4050 658 4214 661
rect 4410 658 4414 661
rect 4534 658 4590 661
rect 4738 658 4750 661
rect 4762 658 4926 661
rect 4930 658 4982 661
rect 4990 661 4993 668
rect 4986 658 4993 661
rect 5002 658 5014 661
rect 5062 658 5142 661
rect 178 648 206 651
rect 286 648 305 651
rect 330 648 446 651
rect 482 648 518 651
rect 522 648 550 651
rect 826 648 870 651
rect 874 648 894 651
rect 970 648 982 651
rect 1138 648 1222 651
rect 1226 648 1278 651
rect 1282 648 1294 651
rect 1298 648 1382 651
rect 1386 648 1606 651
rect 1610 648 1630 651
rect 1634 648 1718 651
rect 1758 648 1766 651
rect 1770 648 1822 651
rect 1922 648 1950 651
rect 2002 648 2070 651
rect 2146 648 2150 651
rect 2170 648 2222 651
rect 2266 648 2334 651
rect 2354 648 2366 651
rect 2458 648 2470 651
rect 2610 648 2622 651
rect 2682 648 2790 651
rect 2890 648 2902 651
rect 2926 648 2934 651
rect 2938 648 2950 651
rect 3026 648 3254 651
rect 3422 651 3425 658
rect 4534 652 4537 658
rect 4598 652 4601 658
rect 5062 652 5065 658
rect 3422 648 3494 651
rect 3522 648 3526 651
rect 3682 648 3753 651
rect 3938 648 3982 651
rect 4202 648 4206 651
rect 4474 648 4486 651
rect 4722 648 4726 651
rect 4754 648 4798 651
rect 286 642 289 648
rect 302 642 305 648
rect 354 638 366 641
rect 370 638 377 641
rect 426 638 478 641
rect 498 638 606 641
rect 730 638 846 641
rect 874 638 878 641
rect 890 638 1318 641
rect 1326 638 1374 641
rect 1482 638 1518 641
rect 1594 638 1609 641
rect 1634 638 1646 641
rect 1734 641 1737 648
rect 3750 642 3753 648
rect 4070 642 4073 648
rect 1734 638 1766 641
rect 1970 638 2054 641
rect 2090 638 3054 641
rect 3186 638 3190 641
rect 3258 638 3470 641
rect 3506 638 3534 641
rect 4162 638 4182 641
rect 4386 638 4462 641
rect 4706 638 4750 641
rect 1326 632 1329 638
rect 1606 632 1609 638
rect 3862 632 3865 638
rect 274 628 566 631
rect 826 628 1006 631
rect 1450 628 1494 631
rect 1986 628 1990 631
rect 2426 628 2462 631
rect 2570 628 2598 631
rect 2618 628 2622 631
rect 2670 628 2718 631
rect 2754 628 3006 631
rect 3010 628 3014 631
rect 3178 628 3486 631
rect 3890 628 4086 631
rect 4098 628 4190 631
rect 4282 628 4822 631
rect 2670 622 2673 628
rect 298 618 422 621
rect 426 618 494 621
rect 1002 618 1070 621
rect 1274 618 1366 621
rect 1482 618 1814 621
rect 2578 618 2630 621
rect 2850 618 3166 621
rect 3170 618 3478 621
rect 3514 618 3670 621
rect 3674 618 3742 621
rect 3746 618 3950 621
rect 4026 618 4606 621
rect 4610 618 4622 621
rect 4650 618 4654 621
rect 1002 608 1006 611
rect 1234 608 1510 611
rect 2890 608 2958 611
rect 3002 608 3214 611
rect 3226 608 3502 611
rect 3506 608 3566 611
rect 3730 608 3742 611
rect 3794 608 3806 611
rect 3810 608 3926 611
rect 3930 608 4238 611
rect 4242 608 4454 611
rect 536 603 538 607
rect 542 603 545 607
rect 550 603 552 607
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1574 603 1576 607
rect 2584 603 2586 607
rect 2590 603 2593 607
rect 2598 603 2600 607
rect 3608 603 3610 607
rect 3614 603 3617 607
rect 3622 603 3624 607
rect 4632 603 4634 607
rect 4638 603 4641 607
rect 4646 603 4648 607
rect 594 598 750 601
rect 1338 598 1526 601
rect 1682 598 1702 601
rect 2338 598 2414 601
rect 2418 598 2446 601
rect 3314 598 3382 601
rect 3386 598 3398 601
rect 3458 598 3518 601
rect 3866 598 3958 601
rect 4098 598 4374 601
rect 3566 592 3569 598
rect 362 588 534 591
rect 538 588 950 591
rect 1018 588 1502 591
rect 1658 588 1702 591
rect 1706 588 1974 591
rect 2034 588 2246 591
rect 2322 588 2838 591
rect 2874 588 2990 591
rect 3018 588 3046 591
rect 3050 588 3118 591
rect 3346 588 3406 591
rect 3434 588 3526 591
rect 3530 588 3542 591
rect 3818 588 3838 591
rect 3850 588 3854 591
rect 3954 588 4270 591
rect 4374 588 4926 591
rect 4930 588 5030 591
rect 234 578 238 581
rect 242 578 254 581
rect 570 578 622 581
rect 1282 578 1473 581
rect 1890 578 2022 581
rect 2026 578 2046 581
rect 2066 578 2398 581
rect 2402 578 2726 581
rect 2970 578 2974 581
rect 3026 578 3094 581
rect 3098 578 3438 581
rect 3522 578 3590 581
rect 3594 578 3782 581
rect 3786 578 3822 581
rect 3850 578 3902 581
rect 4374 581 4377 588
rect 4194 578 4377 581
rect 4602 578 4758 581
rect 4762 578 4766 581
rect 106 568 137 571
rect 154 568 254 571
rect 258 568 382 571
rect 386 568 454 571
rect 458 568 574 571
rect 610 568 646 571
rect 650 568 846 571
rect 850 568 886 571
rect 926 571 929 578
rect 1470 572 1473 578
rect 926 568 1078 571
rect 1194 568 1262 571
rect 1318 568 1350 571
rect 1818 568 1862 571
rect 2006 568 2022 571
rect 2098 568 2190 571
rect 2194 568 2214 571
rect 2930 568 2990 571
rect 3394 568 3438 571
rect 3554 568 3582 571
rect 3626 568 3646 571
rect 3738 568 3758 571
rect 3770 568 3790 571
rect 3810 568 3814 571
rect 3830 571 3833 578
rect 3830 568 3878 571
rect 4070 571 4073 578
rect 4070 568 4166 571
rect 4890 568 5062 571
rect 5066 568 5078 571
rect 134 562 137 568
rect 1318 562 1321 568
rect 2006 562 2009 568
rect 42 558 118 561
rect 138 558 182 561
rect 346 558 478 561
rect 614 558 622 561
rect 626 558 686 561
rect 786 558 790 561
rect 906 558 910 561
rect 930 558 934 561
rect 946 558 950 561
rect 1682 558 1694 561
rect 1770 558 1862 561
rect 2018 558 2022 561
rect 2026 558 2054 561
rect 2122 558 2158 561
rect 2210 558 2310 561
rect 2314 558 2366 561
rect 2370 558 2382 561
rect 2478 561 2481 568
rect 2478 558 2638 561
rect 2842 558 2966 561
rect 2974 558 3086 561
rect 3090 558 3198 561
rect 3214 561 3217 568
rect 3366 561 3369 568
rect 3470 562 3473 568
rect 3214 558 3369 561
rect 3378 558 3398 561
rect 3402 558 3454 561
rect 3570 558 3574 561
rect 3578 558 4094 561
rect 4390 561 4393 568
rect 4390 558 4454 561
rect 4654 561 4657 568
rect 4634 558 4657 561
rect 4914 558 4974 561
rect 206 552 209 558
rect 262 552 265 558
rect 886 552 889 558
rect 1014 552 1017 558
rect 1030 552 1033 558
rect 98 548 158 551
rect 194 548 201 551
rect 274 548 390 551
rect 618 548 622 551
rect 634 548 758 551
rect 874 548 878 551
rect 922 548 990 551
rect 1066 548 1070 551
rect 1146 548 1182 551
rect 1246 551 1249 558
rect 1486 552 1489 558
rect 1246 548 1270 551
rect 1334 548 1406 551
rect 1546 548 1550 551
rect 1626 548 1678 551
rect 1730 548 1734 551
rect 1810 548 1902 551
rect 1926 551 1929 558
rect 1926 548 2030 551
rect 2110 548 2174 551
rect 2250 548 2262 551
rect 2306 548 2326 551
rect 2694 551 2697 558
rect 2474 548 2518 551
rect 862 542 865 548
rect 1334 542 1337 548
rect 1702 542 1705 548
rect 2110 542 2113 548
rect 98 538 126 541
rect 218 538 310 541
rect 570 538 574 541
rect 618 538 630 541
rect 650 538 686 541
rect 722 538 766 541
rect 794 538 814 541
rect 850 538 854 541
rect 930 538 934 541
rect 1034 538 1038 541
rect 1074 538 1158 541
rect 1162 538 1286 541
rect 1602 538 1670 541
rect 1722 538 1830 541
rect 1834 538 1958 541
rect 1994 538 2057 541
rect 2122 538 2126 541
rect 2278 541 2281 548
rect 2694 548 2750 551
rect 2802 548 2806 551
rect 2858 548 2958 551
rect 2974 551 2977 558
rect 4102 552 4105 558
rect 2962 548 2977 551
rect 3014 548 3142 551
rect 3146 548 3174 551
rect 3266 548 3318 551
rect 3338 548 3358 551
rect 3426 548 3430 551
rect 3450 548 3478 551
rect 3522 548 3526 551
rect 3562 548 3582 551
rect 3666 548 4006 551
rect 4034 548 4046 551
rect 4058 548 4062 551
rect 4186 548 4230 551
rect 4234 548 4262 551
rect 4482 548 4518 551
rect 4522 548 4598 551
rect 4602 548 4646 551
rect 4850 548 4862 551
rect 4882 548 4934 551
rect 5050 548 5134 551
rect 2146 538 2281 541
rect 2298 538 2302 541
rect 2386 538 2497 541
rect 2746 538 2774 541
rect 2778 538 2918 541
rect 2922 538 2950 541
rect 3014 541 3017 548
rect 3182 542 3185 548
rect 2954 538 3017 541
rect 3074 538 3134 541
rect 3186 538 3254 541
rect 3314 538 3326 541
rect 3406 541 3409 548
rect 3406 538 3438 541
rect 3450 538 3454 541
rect 3630 541 3633 548
rect 4414 542 4417 548
rect 4422 542 4425 548
rect 4742 542 4745 548
rect 3514 538 3633 541
rect 3682 538 3790 541
rect 3810 538 3862 541
rect 3906 538 3926 541
rect 4002 538 4086 541
rect 4210 538 4214 541
rect 4218 538 4294 541
rect 4298 538 4390 541
rect 4450 538 4606 541
rect 4626 538 4638 541
rect 4786 538 4798 541
rect 4818 538 4862 541
rect 4866 538 4870 541
rect 5050 538 5054 541
rect 5058 538 5078 541
rect 90 528 94 531
rect 166 531 169 538
rect 1014 532 1017 538
rect 2054 532 2057 538
rect 2494 532 2497 538
rect 3342 532 3345 538
rect 4654 532 4657 538
rect 162 528 169 531
rect 442 528 886 531
rect 1034 528 1182 531
rect 1194 528 1198 531
rect 1306 528 1398 531
rect 1418 528 1566 531
rect 1570 528 1646 531
rect 1650 528 1742 531
rect 1762 528 1878 531
rect 1882 528 1966 531
rect 2302 528 2310 531
rect 2314 528 2398 531
rect 2682 528 2729 531
rect 2762 528 2958 531
rect 3154 528 3334 531
rect 3370 528 3414 531
rect 3586 528 4430 531
rect 4562 528 4582 531
rect 4810 528 4894 531
rect 4898 528 4918 531
rect 4922 528 5054 531
rect 2726 522 2729 528
rect 4478 522 4481 528
rect 4494 522 4497 528
rect 4750 522 4753 528
rect 66 518 198 521
rect 506 518 670 521
rect 690 518 766 521
rect 842 518 846 521
rect 1074 518 1102 521
rect 1402 518 1478 521
rect 1514 518 1710 521
rect 1714 518 1758 521
rect 1762 518 1934 521
rect 1938 518 2014 521
rect 2314 518 2318 521
rect 2330 518 2430 521
rect 2818 518 2830 521
rect 2938 518 2950 521
rect 2994 518 3334 521
rect 3338 518 3374 521
rect 3378 518 3526 521
rect 3578 518 3654 521
rect 3818 518 3854 521
rect 3930 518 4054 521
rect 4138 518 4398 521
rect 4554 518 4593 521
rect 886 512 889 518
rect 4590 512 4593 518
rect 106 508 246 511
rect 306 508 638 511
rect 650 508 782 511
rect 1234 508 1238 511
rect 1242 508 1534 511
rect 1802 508 1806 511
rect 2314 508 2342 511
rect 2506 508 2566 511
rect 3418 508 3422 511
rect 3458 508 3470 511
rect 3482 508 3582 511
rect 3626 508 3686 511
rect 3786 508 3798 511
rect 3802 508 3822 511
rect 3826 508 3886 511
rect 4034 508 4094 511
rect 4162 508 4254 511
rect 4602 508 4622 511
rect 1048 503 1050 507
rect 1054 503 1057 507
rect 1062 503 1064 507
rect 2072 503 2074 507
rect 2078 503 2081 507
rect 2086 503 2088 507
rect 3096 503 3098 507
rect 3102 503 3105 507
rect 3110 503 3112 507
rect 3174 502 3177 508
rect 4112 503 4114 507
rect 4118 503 4121 507
rect 4126 503 4128 507
rect 482 498 590 501
rect 602 498 630 501
rect 778 498 950 501
rect 1690 498 1758 501
rect 2042 498 2062 501
rect 2106 498 2462 501
rect 2466 498 2878 501
rect 2922 498 3038 501
rect 3258 498 3278 501
rect 3466 498 3486 501
rect 3882 498 3894 501
rect 3898 498 3926 501
rect 4194 498 4230 501
rect 4258 498 4318 501
rect 4362 498 4718 501
rect 4826 498 4846 501
rect 562 488 758 491
rect 906 488 1190 491
rect 1354 488 1438 491
rect 1618 488 1734 491
rect 1826 488 1990 491
rect 2042 488 2174 491
rect 2178 488 2270 491
rect 2354 488 2662 491
rect 2866 488 2902 491
rect 3002 488 3390 491
rect 3394 488 3574 491
rect 3594 488 3745 491
rect 3874 488 3934 491
rect 3938 488 3982 491
rect 4242 488 4278 491
rect 4378 488 4470 491
rect 4490 488 4758 491
rect 4762 488 4766 491
rect 4954 488 5038 491
rect 14 481 17 488
rect 1494 482 1497 488
rect 14 478 86 481
rect 90 478 150 481
rect 154 478 158 481
rect 754 478 790 481
rect 794 478 822 481
rect 834 478 926 481
rect 942 478 1086 481
rect 1282 478 1366 481
rect 1466 478 1470 481
rect 1742 481 1745 488
rect 3742 482 3745 488
rect 1682 478 1745 481
rect 1778 478 1782 481
rect 1826 478 1846 481
rect 1850 478 1886 481
rect 2010 478 2046 481
rect 2074 478 2126 481
rect 2258 478 2334 481
rect 2346 478 2510 481
rect 2514 478 2646 481
rect 2722 478 2782 481
rect 2818 478 2862 481
rect 3042 478 3174 481
rect 3178 478 3270 481
rect 3450 478 3462 481
rect 3466 478 3510 481
rect 3642 478 3678 481
rect 3746 478 3846 481
rect 3954 478 3974 481
rect 3978 478 4046 481
rect 4266 478 4510 481
rect 4514 478 4534 481
rect 4686 478 4710 481
rect 34 468 102 471
rect 274 468 321 471
rect 354 468 358 471
rect 410 468 414 471
rect 422 468 430 471
rect 490 468 494 471
rect 654 471 657 478
rect 942 472 945 478
rect 654 468 694 471
rect 770 468 782 471
rect 810 468 838 471
rect 930 468 934 471
rect 1042 468 1046 471
rect 1082 468 1134 471
rect 1206 471 1209 478
rect 1278 472 1281 478
rect 1766 472 1769 478
rect 2654 472 2657 478
rect 2670 472 2673 478
rect 2966 472 2969 478
rect 3406 472 3409 478
rect 4086 472 4089 478
rect 4182 472 4185 478
rect 4686 472 4689 478
rect 4734 472 4737 478
rect 1206 468 1214 471
rect 1342 468 1350 471
rect 1354 468 1382 471
rect 1418 468 1502 471
rect 1514 468 1518 471
rect 1562 468 1606 471
rect 1610 468 1737 471
rect 1858 468 1934 471
rect 2266 468 2382 471
rect 2402 468 2406 471
rect 2426 468 2430 471
rect 2498 468 2542 471
rect 2826 468 2830 471
rect 2834 468 2878 471
rect 3138 468 3190 471
rect 3218 468 3294 471
rect 3434 468 3438 471
rect 3458 468 3494 471
rect 3738 468 3782 471
rect 3970 468 4038 471
rect 4202 468 4222 471
rect 4226 468 4254 471
rect 4314 468 4318 471
rect 4330 468 4374 471
rect 4394 468 4438 471
rect 4458 468 4662 471
rect 4666 468 4686 471
rect 4830 468 4878 471
rect 5058 468 5070 471
rect 42 458 78 461
rect 150 461 153 468
rect 318 462 321 468
rect 454 462 457 468
rect 150 458 182 461
rect 194 458 286 461
rect 338 458 398 461
rect 402 458 406 461
rect 618 458 622 461
rect 778 458 806 461
rect 818 458 870 461
rect 962 458 966 461
rect 1002 458 1006 461
rect 1010 458 1166 461
rect 1170 458 1694 461
rect 1722 458 1726 461
rect 1734 461 1737 468
rect 2022 462 2025 468
rect 1734 458 2006 461
rect 2054 461 2057 468
rect 2118 461 2121 468
rect 2054 458 2121 461
rect 2150 461 2153 468
rect 2150 458 2262 461
rect 2282 458 2430 461
rect 2490 458 2614 461
rect 2634 458 2678 461
rect 2798 461 2801 468
rect 2730 458 2801 461
rect 2810 458 2830 461
rect 2850 458 2982 461
rect 2986 458 3038 461
rect 3110 461 3113 468
rect 3042 458 3113 461
rect 3130 458 3254 461
rect 3314 458 3494 461
rect 3654 461 3657 468
rect 3634 458 3657 461
rect 3670 461 3673 468
rect 3670 458 3774 461
rect 3826 459 3870 461
rect 4830 462 4833 468
rect 3826 458 3873 459
rect 4018 458 4430 461
rect 4434 458 4446 461
rect 4594 458 4782 461
rect 4794 458 4806 461
rect 4858 458 4894 461
rect 5006 461 5009 468
rect 5006 458 5062 461
rect 114 448 142 451
rect 146 448 238 451
rect 242 448 342 451
rect 546 448 617 451
rect 634 448 638 451
rect 698 448 769 451
rect 162 438 177 441
rect 186 438 222 441
rect 438 441 441 448
rect 410 438 441 441
rect 614 442 617 448
rect 766 442 769 448
rect 782 448 809 451
rect 826 448 902 451
rect 938 448 1030 451
rect 1082 448 1118 451
rect 1486 448 1505 451
rect 782 442 785 448
rect 806 442 809 448
rect 1486 442 1489 448
rect 1502 442 1505 448
rect 1726 448 1734 451
rect 2314 448 2350 451
rect 2414 448 2446 451
rect 2554 448 2694 451
rect 2778 448 2814 451
rect 2818 448 2830 451
rect 3058 448 3718 451
rect 3722 448 3878 451
rect 4170 448 4406 451
rect 4426 448 4502 451
rect 4506 448 4526 451
rect 4538 448 4814 451
rect 1518 442 1521 448
rect 666 438 678 441
rect 842 438 950 441
rect 1018 438 1342 441
rect 1346 438 1470 441
rect 1710 441 1713 448
rect 1626 438 1713 441
rect 1726 442 1729 448
rect 2382 442 2385 448
rect 2414 442 2417 448
rect 2494 442 2497 448
rect 4414 442 4417 448
rect 2274 438 2374 441
rect 2666 438 2790 441
rect 2938 438 2990 441
rect 3106 438 3438 441
rect 3554 438 3982 441
rect 3986 438 4230 441
rect 4362 438 4366 441
rect 4942 441 4945 448
rect 4498 438 4945 441
rect 174 432 177 438
rect 290 428 470 431
rect 634 428 774 431
rect 782 428 926 431
rect 1018 428 1102 431
rect 1346 428 1422 431
rect 1458 428 1878 431
rect 1882 428 2086 431
rect 2442 428 3014 431
rect 3018 428 3134 431
rect 3178 428 3398 431
rect 3478 431 3481 438
rect 3478 428 3566 431
rect 3834 428 3862 431
rect 4266 428 4806 431
rect 162 418 206 421
rect 782 421 785 428
rect 602 418 785 421
rect 794 418 822 421
rect 858 418 870 421
rect 1066 418 1270 421
rect 1698 418 1782 421
rect 1914 418 2054 421
rect 2098 418 2110 421
rect 2346 418 2406 421
rect 2866 418 2886 421
rect 2890 418 2990 421
rect 2994 418 3102 421
rect 3530 418 3790 421
rect 3794 418 3798 421
rect 4242 418 4382 421
rect 4386 418 4406 421
rect 4410 418 4558 421
rect 4746 418 5182 421
rect 762 408 766 411
rect 802 408 846 411
rect 858 408 1030 411
rect 1434 408 1542 411
rect 1722 408 1910 411
rect 2058 408 2334 411
rect 2354 408 2470 411
rect 2658 408 2702 411
rect 2706 408 2742 411
rect 2778 408 2846 411
rect 2962 408 2974 411
rect 3002 408 3374 411
rect 3754 408 3814 411
rect 4074 408 4150 411
rect 4154 408 4182 411
rect 4186 408 4334 411
rect 4338 408 4430 411
rect 536 403 538 407
rect 542 403 545 407
rect 550 403 552 407
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1574 403 1576 407
rect 2584 403 2586 407
rect 2590 403 2593 407
rect 2598 403 2600 407
rect 3608 403 3610 407
rect 3614 403 3617 407
rect 3622 403 3624 407
rect 4632 403 4634 407
rect 4638 403 4641 407
rect 4646 403 4648 407
rect 618 398 1014 401
rect 1106 398 1174 401
rect 1226 398 1230 401
rect 1258 398 1502 401
rect 2010 398 2110 401
rect 2114 398 2190 401
rect 2322 398 2438 401
rect 2658 398 2774 401
rect 2794 398 2846 401
rect 2850 398 3038 401
rect 3042 398 3150 401
rect 3450 398 3470 401
rect 3642 398 3646 401
rect 3658 398 3678 401
rect 3682 398 3694 401
rect 3850 398 4030 401
rect 4274 398 4382 401
rect 4386 398 4622 401
rect 74 388 86 391
rect 90 388 158 391
rect 170 388 174 391
rect 178 388 366 391
rect 370 388 814 391
rect 818 388 1086 391
rect 1130 388 1182 391
rect 1422 388 1430 391
rect 1434 388 1438 391
rect 1466 388 1526 391
rect 1970 388 2174 391
rect 2178 388 2302 391
rect 2306 388 2350 391
rect 2358 388 2366 391
rect 2370 388 2454 391
rect 2626 388 2718 391
rect 2738 388 2814 391
rect 2838 388 2846 391
rect 2850 388 3006 391
rect 3018 388 3118 391
rect 3122 388 3150 391
rect 3298 388 3790 391
rect 3794 388 3806 391
rect 3810 388 3886 391
rect 4426 388 4854 391
rect 282 378 350 381
rect 506 378 590 381
rect 682 378 1270 381
rect 1402 378 1446 381
rect 1514 378 1550 381
rect 2034 378 2054 381
rect 2130 378 2774 381
rect 2882 378 3046 381
rect 3578 378 3982 381
rect 4690 378 4862 381
rect 1758 372 1761 378
rect 326 368 393 371
rect 326 362 329 368
rect 390 362 393 368
rect 810 368 814 371
rect 914 368 974 371
rect 1074 368 1078 371
rect 1098 368 1118 371
rect 1170 368 1214 371
rect 1226 368 1230 371
rect 1242 368 1246 371
rect 1290 368 1294 371
rect 1330 368 1334 371
rect 1394 368 1414 371
rect 1426 368 1462 371
rect 1530 368 1545 371
rect 1578 368 1654 371
rect 1658 368 1662 371
rect 2094 371 2097 378
rect 3454 372 3457 378
rect 1978 368 2097 371
rect 2150 368 2158 371
rect 2162 368 2262 371
rect 2266 368 2278 371
rect 2290 368 2329 371
rect 414 362 417 368
rect 1542 362 1545 368
rect 1734 362 1737 368
rect 358 358 382 361
rect 394 358 406 361
rect 450 358 478 361
rect 626 358 654 361
rect 658 358 1534 361
rect 1570 358 1670 361
rect 1698 358 1702 361
rect 1750 361 1753 368
rect 1766 361 1769 368
rect 2326 362 2329 368
rect 2418 368 2510 371
rect 2514 368 2606 371
rect 2866 368 2998 371
rect 3026 368 3206 371
rect 3282 368 3310 371
rect 3314 368 3334 371
rect 3466 368 3486 371
rect 3502 371 3505 378
rect 3502 368 3518 371
rect 3682 368 3686 371
rect 3818 368 3838 371
rect 3850 368 3854 371
rect 3922 368 4078 371
rect 4082 368 4166 371
rect 4394 368 4406 371
rect 4410 368 4513 371
rect 1750 358 1769 361
rect 2066 358 2318 361
rect 2374 361 2377 368
rect 2390 361 2393 368
rect 2374 358 2393 361
rect 2694 361 2697 368
rect 2562 358 2697 361
rect 2714 358 2718 361
rect 2806 361 2809 368
rect 2802 358 2809 361
rect 2954 358 2974 361
rect 2986 358 2998 361
rect 3058 358 3646 361
rect 3650 358 3822 361
rect 3826 358 3902 361
rect 4198 361 4201 368
rect 4510 362 4513 368
rect 4570 368 4798 371
rect 4858 368 4918 371
rect 4922 368 5062 371
rect 5066 368 5086 371
rect 4198 358 4206 361
rect 4346 358 4358 361
rect 4526 361 4529 368
rect 4526 358 4534 361
rect 4586 358 4678 361
rect 4778 358 4966 361
rect 358 352 361 358
rect 122 348 150 351
rect 154 348 174 351
rect 210 348 214 351
rect 346 348 350 351
rect 450 348 542 351
rect 102 342 105 348
rect 550 348 606 351
rect 610 348 782 351
rect 786 348 1430 351
rect 1442 348 1462 351
rect 1466 348 1502 351
rect 1506 348 1870 351
rect 1910 351 1913 358
rect 3966 352 3969 358
rect 4030 352 4033 358
rect 4070 352 4073 358
rect 4134 352 4137 358
rect 4478 352 4481 358
rect 4518 352 4521 358
rect 1910 348 1934 351
rect 2018 348 2654 351
rect 2682 348 2686 351
rect 2690 348 2710 351
rect 2714 348 2782 351
rect 2818 348 2854 351
rect 2874 348 2966 351
rect 3030 348 3097 351
rect 82 338 102 341
rect 130 338 222 341
rect 410 338 438 341
rect 550 341 553 348
rect 2982 342 2985 348
rect 3030 342 3033 348
rect 3094 342 3097 348
rect 3226 348 3278 351
rect 3298 348 3310 351
rect 3410 348 3457 351
rect 3466 348 3478 351
rect 3482 348 3526 351
rect 3546 348 3673 351
rect 3682 348 3726 351
rect 3834 348 3854 351
rect 4170 348 4190 351
rect 4210 348 4214 351
rect 4354 348 4406 351
rect 4538 348 4542 351
rect 4742 351 4745 358
rect 4562 348 4782 351
rect 5006 351 5009 358
rect 4794 348 5009 351
rect 5018 348 5054 351
rect 458 338 553 341
rect 578 338 614 341
rect 666 338 670 341
rect 738 338 822 341
rect 866 338 870 341
rect 914 338 953 341
rect 1114 338 1118 341
rect 1178 338 1305 341
rect 1426 338 1494 341
rect 1498 338 1542 341
rect 1714 338 1734 341
rect 1754 338 1838 341
rect 1850 338 1945 341
rect 1994 338 2022 341
rect 2042 338 2134 341
rect 2146 338 2174 341
rect 2178 338 2286 341
rect 2290 338 2358 341
rect 2722 338 2774 341
rect 2778 338 2974 341
rect 3190 341 3193 348
rect 3454 342 3457 348
rect 3670 342 3673 348
rect 3798 342 3801 348
rect 3878 342 3881 348
rect 3130 338 3193 341
rect 3258 338 3270 341
rect 3274 338 3366 341
rect 3490 338 3550 341
rect 3682 338 3734 341
rect 3818 338 3870 341
rect 4066 338 4198 341
rect 4474 338 4526 341
rect 4562 338 4758 341
rect 4794 338 5046 341
rect 5050 338 5062 341
rect 5066 338 5094 341
rect 950 332 953 338
rect 1302 332 1305 338
rect 1942 332 1945 338
rect 178 328 182 331
rect 186 328 190 331
rect 338 328 798 331
rect 1058 328 1070 331
rect 1090 328 1110 331
rect 1114 328 1206 331
rect 1306 328 1414 331
rect 1466 328 1502 331
rect 1526 328 1606 331
rect 2018 328 2126 331
rect 2130 328 2318 331
rect 2690 328 2734 331
rect 2738 328 2894 331
rect 3162 328 3326 331
rect 3338 328 3558 331
rect 3918 331 3921 338
rect 3842 328 3921 331
rect 4018 328 4422 331
rect 4426 328 4566 331
rect 4762 328 4870 331
rect 4874 328 4910 331
rect 166 322 169 328
rect 1526 322 1529 328
rect 234 318 422 321
rect 466 318 574 321
rect 586 318 598 321
rect 1226 318 1446 321
rect 1474 318 1478 321
rect 1546 318 1726 321
rect 1730 318 1766 321
rect 1770 318 1830 321
rect 2158 318 2166 321
rect 2170 318 2214 321
rect 2242 318 2334 321
rect 2338 318 2342 321
rect 2378 318 2398 321
rect 2686 318 2798 321
rect 2802 318 2902 321
rect 2906 318 3006 321
rect 3010 318 3150 321
rect 3242 318 3366 321
rect 3442 318 3590 321
rect 3858 318 4062 321
rect 4106 318 4230 321
rect 4234 318 4238 321
rect 4522 318 4734 321
rect 4750 321 4753 328
rect 4750 318 4766 321
rect 4802 318 4814 321
rect 4834 318 4886 321
rect 2686 312 2689 318
rect 202 308 286 311
rect 402 308 422 311
rect 442 308 726 311
rect 978 308 1006 311
rect 1266 308 1270 311
rect 1434 308 1534 311
rect 1538 308 1606 311
rect 1962 308 2014 311
rect 2138 308 2278 311
rect 2282 308 2326 311
rect 2330 308 2374 311
rect 2386 308 2686 311
rect 2762 308 2870 311
rect 2882 308 3022 311
rect 3130 308 3446 311
rect 3450 308 3662 311
rect 3842 308 3950 311
rect 3962 308 3998 311
rect 4242 308 4286 311
rect 4306 308 4358 311
rect 4410 308 4590 311
rect 4594 308 4614 311
rect 4626 308 4670 311
rect 1048 303 1050 307
rect 1054 303 1057 307
rect 1062 303 1064 307
rect 2072 303 2074 307
rect 2078 303 2081 307
rect 2086 303 2088 307
rect 3096 303 3098 307
rect 3102 303 3105 307
rect 3110 303 3112 307
rect 4112 303 4114 307
rect 4118 303 4121 307
rect 4126 303 4128 307
rect 162 298 174 301
rect 186 298 310 301
rect 314 298 374 301
rect 378 298 430 301
rect 434 298 470 301
rect 474 298 566 301
rect 578 298 598 301
rect 1210 298 1302 301
rect 1546 298 1950 301
rect 2098 298 2206 301
rect 2290 298 2318 301
rect 2442 298 2734 301
rect 2738 298 2870 301
rect 3130 298 3166 301
rect 3258 298 3326 301
rect 3338 298 3422 301
rect 3674 298 3710 301
rect 3714 298 3750 301
rect 4410 298 4518 301
rect 4526 298 4574 301
rect 4594 298 4686 301
rect 4698 298 4806 301
rect 5066 298 5126 301
rect 50 288 222 291
rect 322 288 366 291
rect 410 288 606 291
rect 722 288 750 291
rect 890 288 966 291
rect 970 288 982 291
rect 1066 288 1102 291
rect 1106 288 1270 291
rect 1610 288 1718 291
rect 1810 288 1958 291
rect 2186 288 2214 291
rect 2218 288 2230 291
rect 2274 288 2286 291
rect 2394 288 2406 291
rect 2418 288 2446 291
rect 2642 288 2646 291
rect 2834 288 2862 291
rect 3002 288 3014 291
rect 3066 288 3198 291
rect 3202 288 3294 291
rect 3314 288 3358 291
rect 3362 288 3430 291
rect 3634 288 3726 291
rect 3754 288 3758 291
rect 3762 288 3782 291
rect 4050 288 4350 291
rect 4358 291 4361 298
rect 4358 288 4374 291
rect 4526 291 4529 298
rect 4474 288 4529 291
rect 4658 288 4702 291
rect 4706 288 4726 291
rect 4898 288 4918 291
rect 4922 288 5038 291
rect 5106 288 5110 291
rect 5186 288 5190 291
rect 1534 282 1537 288
rect 66 278 102 281
rect 106 278 638 281
rect 642 278 734 281
rect 738 278 750 281
rect 754 278 918 281
rect 922 278 982 281
rect 986 278 1270 281
rect 1274 278 1310 281
rect 1330 278 1358 281
rect 1362 278 1470 281
rect 1586 278 1726 281
rect 1858 278 1870 281
rect 2194 278 2302 281
rect 2450 278 2462 281
rect 2794 278 2806 281
rect 2978 278 3022 281
rect 3034 278 3126 281
rect 3250 278 3318 281
rect 3322 278 3342 281
rect 3346 278 3478 281
rect 3554 278 3598 281
rect 3602 278 3630 281
rect 3746 278 3838 281
rect 3898 278 3934 281
rect 4186 278 4366 281
rect 4458 278 4854 281
rect 1502 272 1505 278
rect 1526 272 1529 278
rect 1926 272 1929 278
rect 2774 272 2777 278
rect 442 268 446 271
rect 458 268 462 271
rect 506 268 614 271
rect 666 268 670 271
rect 690 268 694 271
rect 802 268 918 271
rect 1082 268 1086 271
rect 1154 268 1238 271
rect 1282 268 1302 271
rect 1354 268 1358 271
rect 1402 268 1406 271
rect 1450 268 1486 271
rect 1554 268 1590 271
rect 1602 268 1662 271
rect 1746 268 1798 271
rect 1826 268 1926 271
rect 1946 268 2014 271
rect 2186 268 2382 271
rect 2386 268 2702 271
rect 2730 268 2774 271
rect 2986 268 3310 271
rect 3362 268 3366 271
rect 3550 271 3553 278
rect 3514 268 3553 271
rect 3666 268 3694 271
rect 3718 271 3721 278
rect 4454 272 4457 278
rect 3718 268 3806 271
rect 3810 268 3902 271
rect 3906 268 4014 271
rect 4034 268 4046 271
rect 4058 268 4126 271
rect 4178 268 4190 271
rect 4474 268 4718 271
rect 4770 268 4774 271
rect 4894 268 4942 271
rect 5110 271 5113 278
rect 5110 268 5118 271
rect 1270 262 1273 268
rect 2958 262 2961 268
rect 98 258 134 261
rect 146 258 542 261
rect 546 258 710 261
rect 786 258 817 261
rect 842 258 998 261
rect 1002 258 1070 261
rect 1074 258 1222 261
rect 1338 258 1358 261
rect 1506 258 1622 261
rect 1738 258 1790 261
rect 1794 258 1878 261
rect 1986 258 2070 261
rect 2170 258 2174 261
rect 2218 258 2233 261
rect 2242 258 2254 261
rect 2442 258 2566 261
rect 2610 258 2702 261
rect 2746 258 2958 261
rect 3010 259 3070 261
rect 3310 262 3313 268
rect 3010 258 3073 259
rect 3314 258 3758 261
rect 3778 258 3846 261
rect 3954 258 4110 261
rect 4114 258 4278 261
rect 4382 261 4385 268
rect 4378 258 4385 261
rect 4446 262 4449 268
rect 4894 262 4897 268
rect 4526 258 4606 261
rect 4666 258 4710 261
rect 4714 258 4782 261
rect 4866 258 4870 261
rect 4974 261 4977 268
rect 4974 258 5014 261
rect 5050 258 5078 261
rect 5130 258 5134 261
rect 42 248 113 251
rect 210 248 222 251
rect 426 248 550 251
rect 562 248 606 251
rect 610 248 638 251
rect 710 251 713 258
rect 814 252 817 258
rect 710 248 718 251
rect 722 248 798 251
rect 898 248 910 251
rect 1034 248 1102 251
rect 1238 251 1241 258
rect 1302 252 1305 258
rect 1238 248 1286 251
rect 1478 251 1481 258
rect 2230 252 2233 258
rect 3174 252 3177 258
rect 1378 248 1481 251
rect 1598 248 1617 251
rect 110 242 113 248
rect 1598 242 1601 248
rect 1614 242 1617 248
rect 1746 248 1774 251
rect 1798 248 1806 251
rect 1810 248 1870 251
rect 1962 248 1990 251
rect 2438 248 2510 251
rect 2678 248 2697 251
rect 3114 248 3174 251
rect 3346 248 3390 251
rect 3594 248 3697 251
rect 602 238 614 241
rect 634 238 798 241
rect 802 238 806 241
rect 1058 238 1062 241
rect 1298 238 1486 241
rect 1630 241 1633 248
rect 1630 238 1718 241
rect 1774 241 1777 248
rect 1910 242 1913 248
rect 1774 238 1806 241
rect 1990 241 1993 248
rect 2022 241 2025 248
rect 1990 238 2025 241
rect 2262 241 2265 248
rect 2234 238 2265 241
rect 2438 242 2441 248
rect 2678 242 2681 248
rect 2694 242 2697 248
rect 3694 242 3697 248
rect 3754 248 3758 251
rect 3910 251 3913 258
rect 4526 252 4529 258
rect 3910 248 3974 251
rect 4002 248 4174 251
rect 4214 248 4241 251
rect 4594 248 4710 251
rect 4762 248 4774 251
rect 4858 248 4870 251
rect 2818 238 3022 241
rect 3074 238 3462 241
rect 3538 238 3630 241
rect 3734 241 3737 248
rect 3774 241 3777 248
rect 4214 242 4217 248
rect 4238 242 4241 248
rect 3734 238 3777 241
rect 3786 238 3886 241
rect 4498 238 4542 241
rect 4554 238 4878 241
rect 362 228 478 231
rect 486 228 670 231
rect 922 228 1214 231
rect 1218 228 1254 231
rect 1314 228 1582 231
rect 1690 228 1846 231
rect 1850 228 1950 231
rect 1994 228 2254 231
rect 2258 228 2382 231
rect 2498 228 2790 231
rect 2858 228 2974 231
rect 3042 228 3414 231
rect 3418 228 3502 231
rect 3506 228 3558 231
rect 3562 228 3590 231
rect 3594 228 3638 231
rect 4210 228 4230 231
rect 4234 228 4390 231
rect 4394 228 4622 231
rect 486 221 489 228
rect 330 218 489 221
rect 498 218 646 221
rect 698 218 758 221
rect 762 218 830 221
rect 1114 218 1326 221
rect 1386 218 1582 221
rect 1610 218 1750 221
rect 1754 218 1758 221
rect 1762 218 2014 221
rect 2018 218 2174 221
rect 2178 218 2238 221
rect 2242 218 2286 221
rect 2530 218 2862 221
rect 3034 218 3222 221
rect 3290 218 3382 221
rect 3530 218 3726 221
rect 3730 218 3830 221
rect 4218 218 4238 221
rect 4466 218 4830 221
rect 5026 218 5070 221
rect 762 208 878 211
rect 1258 208 1502 211
rect 1962 208 2054 211
rect 2186 208 2446 211
rect 2698 208 3161 211
rect 3170 208 3470 211
rect 3658 208 4262 211
rect 4530 208 4606 211
rect 4762 208 5110 211
rect 536 203 538 207
rect 542 203 545 207
rect 550 203 552 207
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1574 203 1576 207
rect 2584 203 2586 207
rect 2590 203 2593 207
rect 2598 203 2600 207
rect 570 198 670 201
rect 794 198 926 201
rect 1050 198 1078 201
rect 1114 198 1206 201
rect 1210 198 1310 201
rect 1666 198 1790 201
rect 1850 198 1942 201
rect 2690 198 2721 201
rect 2730 198 2750 201
rect 2754 198 2766 201
rect 3158 201 3161 208
rect 3608 203 3610 207
rect 3614 203 3617 207
rect 3622 203 3624 207
rect 4632 203 4634 207
rect 4638 203 4641 207
rect 4646 203 4648 207
rect 3158 198 3374 201
rect 4058 198 4094 201
rect 4098 198 4102 201
rect 4410 198 4414 201
rect 4418 198 4422 201
rect 4674 198 4734 201
rect 4778 198 4966 201
rect 222 192 225 198
rect 2718 192 2721 198
rect 106 188 166 191
rect 434 188 462 191
rect 466 188 846 191
rect 1074 188 1337 191
rect 1434 188 1550 191
rect 1586 188 1750 191
rect 1754 188 1878 191
rect 1922 188 2030 191
rect 2034 188 2246 191
rect 2722 188 2782 191
rect 2786 188 2894 191
rect 3330 188 3438 191
rect 3442 188 3526 191
rect 3666 188 3710 191
rect 4018 188 4062 191
rect 4146 188 4494 191
rect 4498 188 4502 191
rect 4754 188 4902 191
rect 5106 188 5110 191
rect 1334 182 1337 188
rect 202 178 294 181
rect 514 178 686 181
rect 1202 178 1222 181
rect 1226 178 1246 181
rect 1338 178 1734 181
rect 1890 178 1894 181
rect 1898 178 1910 181
rect 2210 178 2294 181
rect 2702 181 2705 188
rect 2658 178 2705 181
rect 2730 178 3158 181
rect 3402 178 3470 181
rect 3538 178 3710 181
rect 3714 178 3854 181
rect 4074 178 4182 181
rect 4186 178 4254 181
rect 4730 178 4790 181
rect 4794 178 4846 181
rect 4874 178 4998 181
rect 138 168 278 171
rect 290 168 310 171
rect 410 168 494 171
rect 642 168 734 171
rect 854 168 942 171
rect 946 168 966 171
rect 1218 168 1358 171
rect 1714 168 1769 171
rect 1778 168 2158 171
rect 2162 168 2225 171
rect 2326 171 2329 178
rect 2314 168 2329 171
rect 2342 168 2430 171
rect 2434 168 2494 171
rect 2642 168 2686 171
rect 2690 168 2718 171
rect 2738 168 2742 171
rect 2754 168 2758 171
rect 2762 168 2798 171
rect 2814 168 2822 171
rect 2826 168 2830 171
rect 2850 168 2854 171
rect 3178 168 3198 171
rect 3494 171 3497 178
rect 3862 172 3865 178
rect 3218 168 3497 171
rect 3522 168 3638 171
rect 3642 168 3670 171
rect 4010 168 4142 171
rect 4170 168 4198 171
rect 4202 168 4238 171
rect 4258 168 4374 171
rect 4378 168 4446 171
rect 4650 168 4769 171
rect 4818 168 4822 171
rect 854 162 857 168
rect 1454 162 1457 168
rect 1766 162 1769 168
rect 2222 162 2225 168
rect 2342 162 2345 168
rect 4766 162 4769 168
rect 42 158 121 161
rect 186 158 190 161
rect 234 158 430 161
rect 538 158 582 161
rect 586 158 630 161
rect 650 158 702 161
rect 778 158 838 161
rect 1066 158 1254 161
rect 1274 158 1454 161
rect 1466 158 1478 161
rect 1650 158 1726 161
rect 1746 158 1758 161
rect 1770 158 1806 161
rect 1882 158 1974 161
rect 2106 158 2158 161
rect 2282 158 2326 161
rect 2682 158 2854 161
rect 2866 158 2870 161
rect 3354 158 3414 161
rect 3494 158 4174 161
rect 4202 158 4254 161
rect 4330 158 4366 161
rect 4706 158 4750 161
rect 4894 161 4897 168
rect 4894 158 5054 161
rect 118 151 121 158
rect 214 152 217 158
rect 1862 152 1865 158
rect 2510 152 2513 158
rect 118 148 206 151
rect 242 148 254 151
rect 314 148 342 151
rect 378 148 454 151
rect 490 148 510 151
rect 602 148 710 151
rect 754 148 774 151
rect 786 148 790 151
rect 826 148 846 151
rect 1002 148 1086 151
rect 1146 148 1230 151
rect 1314 148 1350 151
rect 1354 148 1406 151
rect 1498 148 1502 151
rect 110 141 113 148
rect 66 138 113 141
rect 238 141 241 148
rect 234 138 241 141
rect 498 138 526 141
rect 530 138 694 141
rect 746 138 798 141
rect 818 138 894 141
rect 1262 141 1265 148
rect 1374 142 1377 148
rect 1446 142 1449 148
rect 1462 142 1465 148
rect 1562 148 1710 151
rect 1714 148 1742 151
rect 1754 148 1758 151
rect 1874 148 1910 151
rect 1914 148 2022 151
rect 2058 148 2126 151
rect 2146 148 2214 151
rect 2322 148 2377 151
rect 2610 148 2662 151
rect 2786 148 2806 151
rect 2826 148 2886 151
rect 2938 148 3086 151
rect 3142 151 3145 158
rect 3090 148 3145 151
rect 3206 152 3209 158
rect 3494 152 3497 158
rect 3314 148 3454 151
rect 3490 148 3494 151
rect 3506 148 3790 151
rect 3818 148 3838 151
rect 4050 148 4118 151
rect 4122 148 4230 151
rect 4246 148 4358 151
rect 4442 148 4510 151
rect 4522 148 4606 151
rect 4754 148 4758 151
rect 4838 151 4841 158
rect 4834 148 4841 151
rect 5166 151 5169 158
rect 5166 148 5174 151
rect 2286 142 2289 148
rect 2374 142 2377 148
rect 2702 142 2705 148
rect 3790 142 3793 148
rect 1258 138 1334 141
rect 1418 138 1430 141
rect 1594 138 1702 141
rect 1706 138 1758 141
rect 1810 138 1854 141
rect 1882 138 1902 141
rect 1938 138 2118 141
rect 2122 138 2182 141
rect 2202 138 2222 141
rect 2250 138 2270 141
rect 2706 138 2782 141
rect 2858 138 2862 141
rect 3242 138 3390 141
rect 3410 138 3414 141
rect 3458 138 3598 141
rect 3650 138 3726 141
rect 3814 138 3910 141
rect 3974 141 3977 148
rect 4246 142 4249 148
rect 4382 142 4385 148
rect 4438 142 4441 148
rect 3954 138 3977 141
rect 3982 138 4110 141
rect 4114 138 4158 141
rect 4210 138 4214 141
rect 4610 138 4742 141
rect 4750 138 4798 141
rect 4902 141 4905 148
rect 4858 138 4905 141
rect 4970 138 5054 141
rect 318 131 321 138
rect 298 128 321 131
rect 426 128 438 131
rect 442 128 550 131
rect 554 128 758 131
rect 802 128 1062 131
rect 1362 128 1510 131
rect 1722 128 1742 131
rect 1802 128 1806 131
rect 2190 131 2193 138
rect 3814 132 3817 138
rect 1814 128 2193 131
rect 2282 128 2318 131
rect 2434 128 2582 131
rect 2682 128 2734 131
rect 2746 128 2918 131
rect 3026 128 3566 131
rect 3570 128 3590 131
rect 3982 131 3985 138
rect 4222 132 4225 138
rect 3826 128 3985 131
rect 4002 128 4078 131
rect 4234 128 4358 131
rect 4362 128 4470 131
rect 4570 128 4574 131
rect 4750 131 4753 138
rect 4626 128 4753 131
rect 4762 128 4894 131
rect 314 118 414 121
rect 418 118 574 121
rect 690 118 790 121
rect 802 118 830 121
rect 834 118 1198 121
rect 1202 118 1318 121
rect 1322 118 1406 121
rect 1814 121 1817 128
rect 1770 118 1817 121
rect 1826 118 1918 121
rect 2254 121 2257 128
rect 2030 118 2257 121
rect 2338 118 2366 121
rect 2690 118 2846 121
rect 3370 118 3670 121
rect 4194 118 4798 121
rect 4810 118 5078 121
rect 2030 112 2033 118
rect 546 108 766 111
rect 770 108 798 111
rect 1074 108 1294 111
rect 1306 108 1358 111
rect 1474 108 1582 111
rect 1586 108 1998 111
rect 2106 108 2174 111
rect 2178 108 2814 111
rect 2826 108 2862 111
rect 3366 111 3369 118
rect 3202 108 3369 111
rect 3498 108 3662 111
rect 3674 108 3982 111
rect 4202 108 4342 111
rect 4602 108 4606 111
rect 4706 108 4894 111
rect 4898 108 5174 111
rect 1048 103 1050 107
rect 1054 103 1057 107
rect 1062 103 1064 107
rect 2072 103 2074 107
rect 2078 103 2081 107
rect 2086 103 2088 107
rect 3096 103 3098 107
rect 3102 103 3105 107
rect 3110 103 3112 107
rect 4022 102 4025 108
rect 4112 103 4114 107
rect 4118 103 4121 107
rect 4126 103 4128 107
rect 538 98 654 101
rect 746 98 750 101
rect 762 98 918 101
rect 1154 98 1342 101
rect 1474 98 1774 101
rect 1786 98 1798 101
rect 2618 98 2838 101
rect 3234 98 3398 101
rect 3442 98 3510 101
rect 3514 98 3774 101
rect 3826 98 4014 101
rect 4034 98 4070 101
rect 4202 98 4230 101
rect 4242 98 4366 101
rect 4386 98 4510 101
rect 4522 98 4782 101
rect 4786 98 4854 101
rect 1990 92 1993 98
rect 4958 92 4961 98
rect 282 88 302 91
rect 306 88 638 91
rect 698 88 806 91
rect 914 88 966 91
rect 1250 88 1329 91
rect 1602 88 1678 91
rect 1682 88 1686 91
rect 1714 88 1774 91
rect 2014 88 2038 91
rect 2074 88 2446 91
rect 2546 88 2742 91
rect 2794 88 2894 91
rect 2898 88 2998 91
rect 3114 88 3230 91
rect 3266 88 3350 91
rect 3642 88 3686 91
rect 3690 88 3950 91
rect 4010 88 4062 91
rect 4066 88 4238 91
rect 4346 88 4462 91
rect 4514 88 4830 91
rect 5010 88 5014 91
rect 1326 82 1329 88
rect 2014 82 2017 88
rect 330 78 454 81
rect 482 78 566 81
rect 914 78 918 81
rect 1010 78 1270 81
rect 1498 78 1614 81
rect 1818 78 1870 81
rect 2050 78 2206 81
rect 2242 78 2350 81
rect 2354 78 2478 81
rect 2570 78 2678 81
rect 2690 78 2750 81
rect 2758 78 2902 81
rect 2986 78 3022 81
rect 3026 78 3310 81
rect 3446 81 3449 88
rect 3478 81 3481 88
rect 3322 78 3449 81
rect 3454 78 3481 81
rect 3986 78 4198 81
rect 4294 78 4302 81
rect 4306 78 4390 81
rect 4402 78 4406 81
rect 4578 78 4838 81
rect 4842 78 4942 81
rect 4954 78 4958 81
rect 5002 78 5038 81
rect 150 71 153 78
rect 82 68 153 71
rect 230 71 233 78
rect 326 71 329 78
rect 758 72 761 78
rect 982 72 985 78
rect 162 68 329 71
rect 506 68 569 71
rect 810 68 934 71
rect 986 68 1225 71
rect 1330 68 1342 71
rect 1346 68 1542 71
rect 1546 68 1582 71
rect 1910 71 1913 78
rect 1782 68 1913 71
rect 1938 68 2022 71
rect 2166 68 2449 71
rect 2758 71 2761 78
rect 2706 68 2761 71
rect 2770 68 2822 71
rect 2850 68 2934 71
rect 2946 68 3054 71
rect 3090 68 3198 71
rect 3218 68 3246 71
rect 3454 71 3457 78
rect 3654 72 3657 78
rect 3662 72 3665 78
rect 3386 68 3457 71
rect 3482 68 3654 71
rect 3854 68 3942 71
rect 3962 68 3990 71
rect 4018 68 4046 71
rect 4098 68 4190 71
rect 4210 68 4214 71
rect 4226 68 4318 71
rect 4370 68 4518 71
rect 4906 68 5126 71
rect 5130 68 5158 71
rect 210 58 350 61
rect 430 61 433 68
rect 566 62 569 68
rect 370 58 433 61
rect 766 61 769 68
rect 1126 62 1129 68
rect 1222 62 1225 68
rect 714 59 769 61
rect 710 58 769 59
rect 794 58 798 61
rect 858 58 926 61
rect 946 58 958 61
rect 962 58 1030 61
rect 1034 58 1070 61
rect 1306 58 1310 61
rect 1426 58 1446 61
rect 1466 58 1542 61
rect 1546 58 1558 61
rect 1578 59 1638 61
rect 1782 62 1785 68
rect 1830 62 1833 68
rect 2166 62 2169 68
rect 2254 62 2257 68
rect 2446 62 2449 68
rect 1578 58 1641 59
rect 1898 58 2102 61
rect 2282 58 2286 61
rect 2378 58 2382 61
rect 2482 58 2630 61
rect 2674 58 2742 61
rect 2762 58 2830 61
rect 3002 58 3030 61
rect 3166 58 3222 61
rect 3474 58 3494 61
rect 3670 61 3673 68
rect 3854 62 3857 68
rect 3870 62 3873 68
rect 4542 62 4545 68
rect 4582 62 4585 68
rect 4686 62 4689 68
rect 3586 58 3673 61
rect 3714 58 3822 61
rect 3914 58 3969 61
rect 3986 58 4017 61
rect 4026 58 4414 61
rect 4754 58 4758 61
rect 4826 58 4846 61
rect 4854 58 4990 61
rect 4994 58 5134 61
rect 438 51 441 58
rect 3166 52 3169 58
rect 3406 52 3409 58
rect 3966 52 3969 58
rect 4014 52 4017 58
rect 4854 52 4857 58
rect 438 48 494 51
rect 658 48 782 51
rect 946 48 953 51
rect 962 48 1390 51
rect 1530 48 1798 51
rect 1802 48 1910 51
rect 2650 48 2654 51
rect 2738 48 2878 51
rect 2882 48 3014 51
rect 3038 48 3046 51
rect 3426 48 3438 51
rect 3490 48 3502 51
rect 3514 48 3598 51
rect 3602 48 3718 51
rect 3722 48 3886 51
rect 3994 48 3998 51
rect 4034 48 4038 51
rect 4058 48 4065 51
rect 4090 48 4110 51
rect 4122 48 4126 51
rect 4234 48 4241 51
rect 950 42 953 48
rect 2686 41 2689 48
rect 2602 38 2689 41
rect 3038 42 3041 48
rect 3990 41 3993 48
rect 3962 38 3993 41
rect 4062 42 4065 48
rect 4238 42 4241 48
rect 4366 48 4393 51
rect 4366 42 4369 48
rect 4390 42 4393 48
rect 4406 48 4446 51
rect 4554 48 4558 51
rect 4818 48 4822 51
rect 4406 42 4409 48
rect 2754 28 2774 31
rect 2778 28 3214 31
rect 3794 28 4606 31
rect 3226 8 3254 11
rect 536 3 538 7
rect 542 3 545 7
rect 550 3 552 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1574 3 1576 7
rect 2584 3 2586 7
rect 2590 3 2593 7
rect 2598 3 2600 7
rect 3608 3 3610 7
rect 3614 3 3617 7
rect 3622 3 3624 7
rect 4632 3 4634 7
rect 4638 3 4641 7
rect 4646 3 4648 7
<< m4contact >>
rect 1050 4903 1054 4907
rect 1058 4903 1061 4907
rect 1061 4903 1062 4907
rect 2074 4903 2078 4907
rect 2082 4903 2085 4907
rect 2085 4903 2086 4907
rect 3098 4903 3102 4907
rect 3106 4903 3109 4907
rect 3109 4903 3110 4907
rect 4114 4903 4118 4907
rect 4122 4903 4125 4907
rect 4125 4903 4126 4907
rect 958 4888 962 4892
rect 582 4868 586 4872
rect 750 4868 754 4872
rect 1814 4868 1818 4872
rect 2350 4868 2354 4872
rect 2438 4868 2442 4872
rect 3678 4868 3682 4872
rect 4806 4868 4810 4872
rect 4878 4868 4882 4872
rect 5062 4868 5066 4872
rect 574 4858 578 4862
rect 1238 4858 1242 4862
rect 1550 4858 1554 4862
rect 1814 4858 1818 4862
rect 2366 4858 2370 4862
rect 2686 4858 2690 4862
rect 3198 4858 3202 4862
rect 3222 4858 3226 4862
rect 4254 4858 4258 4862
rect 4614 4858 4618 4862
rect 4822 4858 4826 4862
rect 4870 4858 4874 4862
rect 4934 4858 4938 4862
rect 5046 4858 5050 4862
rect 5070 4858 5074 4862
rect 5102 4858 5106 4862
rect 4894 4848 4898 4852
rect 4134 4838 4138 4842
rect 4782 4838 4786 4842
rect 5102 4838 5106 4842
rect 750 4828 754 4832
rect 1302 4828 1306 4832
rect 4950 4828 4954 4832
rect 710 4818 714 4822
rect 1422 4818 1426 4822
rect 1886 4818 1890 4822
rect 2438 4818 2442 4822
rect 4046 4818 4050 4822
rect 4934 4818 4938 4822
rect 4982 4818 4986 4822
rect 1670 4808 1674 4812
rect 1750 4808 1754 4812
rect 1766 4808 1770 4812
rect 4366 4808 4370 4812
rect 5014 4808 5018 4812
rect 5094 4808 5098 4812
rect 538 4803 542 4807
rect 546 4803 549 4807
rect 549 4803 550 4807
rect 1562 4803 1566 4807
rect 1570 4803 1573 4807
rect 1573 4803 1574 4807
rect 2586 4803 2590 4807
rect 2594 4803 2597 4807
rect 2597 4803 2598 4807
rect 3610 4803 3614 4807
rect 3618 4803 3621 4807
rect 3621 4803 3622 4807
rect 4634 4803 4638 4807
rect 4642 4803 4645 4807
rect 4645 4803 4646 4807
rect 3246 4798 3250 4802
rect 4446 4798 4450 4802
rect 990 4788 994 4792
rect 2214 4788 2218 4792
rect 4774 4788 4778 4792
rect 5022 4788 5026 4792
rect 4134 4778 4138 4782
rect 2430 4768 2434 4772
rect 4254 4768 4258 4772
rect 174 4758 178 4762
rect 2518 4758 2522 4762
rect 4918 4758 4922 4762
rect 678 4748 682 4752
rect 1182 4748 1186 4752
rect 1358 4748 1362 4752
rect 1510 4748 1514 4752
rect 1622 4748 1626 4752
rect 1638 4748 1642 4752
rect 1686 4748 1690 4752
rect 1702 4748 1706 4752
rect 1814 4748 1818 4752
rect 486 4738 490 4742
rect 646 4738 650 4742
rect 758 4738 762 4742
rect 766 4738 770 4742
rect 1206 4738 1210 4742
rect 4350 4748 4354 4752
rect 4710 4748 4714 4752
rect 2230 4738 2234 4742
rect 2334 4738 2338 4742
rect 2654 4738 2658 4742
rect 3014 4738 3018 4742
rect 4102 4738 4106 4742
rect 4294 4738 4298 4742
rect 1766 4728 1770 4732
rect 2158 4728 2162 4732
rect 2526 4728 2530 4732
rect 294 4718 298 4722
rect 758 4718 762 4722
rect 1326 4718 1330 4722
rect 1902 4718 1906 4722
rect 3870 4718 3874 4722
rect 4510 4718 4514 4722
rect 262 4708 266 4712
rect 574 4708 578 4712
rect 678 4708 682 4712
rect 718 4708 722 4712
rect 1542 4708 1546 4712
rect 4142 4708 4146 4712
rect 1050 4703 1054 4707
rect 1058 4703 1061 4707
rect 1061 4703 1062 4707
rect 2074 4703 2078 4707
rect 2082 4703 2085 4707
rect 2085 4703 2086 4707
rect 3098 4703 3102 4707
rect 3106 4703 3109 4707
rect 3109 4703 3110 4707
rect 4114 4703 4118 4707
rect 4122 4703 4125 4707
rect 4125 4703 4126 4707
rect 1318 4698 1322 4702
rect 3390 4698 3394 4702
rect 3510 4698 3514 4702
rect 4550 4698 4554 4702
rect 4870 4698 4874 4702
rect 134 4688 138 4692
rect 1198 4688 1202 4692
rect 2350 4688 2354 4692
rect 2742 4688 2746 4692
rect 3022 4688 3026 4692
rect 4366 4688 4370 4692
rect 342 4678 346 4682
rect 1230 4678 1234 4682
rect 1894 4678 1898 4682
rect 3246 4678 3250 4682
rect 4214 4678 4218 4682
rect 566 4668 570 4672
rect 878 4668 882 4672
rect 1150 4668 1154 4672
rect 1334 4668 1338 4672
rect 1766 4668 1770 4672
rect 3574 4668 3578 4672
rect 3678 4668 3682 4672
rect 4350 4668 4354 4672
rect 5054 4668 5058 4672
rect 5118 4668 5122 4672
rect 150 4658 154 4662
rect 342 4658 346 4662
rect 430 4658 434 4662
rect 494 4658 498 4662
rect 1214 4658 1218 4662
rect 1310 4658 1314 4662
rect 1390 4658 1394 4662
rect 1622 4658 1626 4662
rect 2030 4658 2034 4662
rect 2230 4658 2234 4662
rect 2262 4658 2266 4662
rect 2694 4658 2698 4662
rect 2990 4658 2994 4662
rect 3030 4658 3034 4662
rect 3558 4658 3562 4662
rect 3646 4658 3650 4662
rect 4054 4658 4058 4662
rect 4166 4658 4170 4662
rect 4446 4658 4450 4662
rect 4598 4658 4602 4662
rect 878 4648 882 4652
rect 1590 4648 1594 4652
rect 1606 4648 1610 4652
rect 654 4638 658 4642
rect 2718 4648 2722 4652
rect 3190 4648 3194 4652
rect 4590 4648 4594 4652
rect 4766 4648 4770 4652
rect 4862 4648 4866 4652
rect 1318 4638 1322 4642
rect 2566 4638 2570 4642
rect 3302 4638 3306 4642
rect 3862 4638 3866 4642
rect 4046 4638 4050 4642
rect 4582 4638 4586 4642
rect 4598 4638 4602 4642
rect 870 4628 874 4632
rect 1310 4628 1314 4632
rect 2262 4628 2266 4632
rect 2534 4628 2538 4632
rect 2758 4628 2762 4632
rect 3086 4628 3090 4632
rect 3222 4628 3226 4632
rect 4134 4628 4138 4632
rect 4422 4628 4426 4632
rect 4550 4628 4554 4632
rect 942 4618 946 4622
rect 1182 4618 1186 4622
rect 1502 4618 1506 4622
rect 2542 4618 2546 4622
rect 2550 4618 2554 4622
rect 3486 4618 3490 4622
rect 3750 4618 3754 4622
rect 4606 4618 4610 4622
rect 558 4608 562 4612
rect 1582 4608 1586 4612
rect 4622 4608 4626 4612
rect 538 4603 542 4607
rect 546 4603 549 4607
rect 549 4603 550 4607
rect 1562 4603 1566 4607
rect 1570 4603 1573 4607
rect 1573 4603 1574 4607
rect 2586 4603 2590 4607
rect 2594 4603 2597 4607
rect 2597 4603 2598 4607
rect 3610 4603 3614 4607
rect 3618 4603 3621 4607
rect 3621 4603 3622 4607
rect 4634 4603 4638 4607
rect 4642 4603 4645 4607
rect 4645 4603 4646 4607
rect 638 4598 642 4602
rect 1382 4598 1386 4602
rect 1230 4588 1234 4592
rect 1526 4588 1530 4592
rect 2038 4588 2042 4592
rect 2798 4588 2802 4592
rect 3878 4588 3882 4592
rect 4246 4588 4250 4592
rect 286 4578 290 4582
rect 558 4578 562 4582
rect 2526 4578 2530 4582
rect 2702 4578 2706 4582
rect 4102 4578 4106 4582
rect 4550 4578 4554 4582
rect 710 4568 714 4572
rect 766 4568 770 4572
rect 822 4568 826 4572
rect 950 4568 954 4572
rect 990 4568 994 4572
rect 2286 4568 2290 4572
rect 3814 4568 3818 4572
rect 1814 4558 1818 4562
rect 2318 4558 2322 4562
rect 2974 4558 2978 4562
rect 3014 4558 3018 4562
rect 4102 4558 4106 4562
rect 4886 4558 4890 4562
rect 5166 4558 5170 4562
rect 486 4548 490 4552
rect 1246 4548 1250 4552
rect 1278 4548 1282 4552
rect 1446 4548 1450 4552
rect 1494 4548 1498 4552
rect 1534 4548 1538 4552
rect 1726 4548 1730 4552
rect 2526 4548 2530 4552
rect 318 4538 322 4542
rect 2910 4548 2914 4552
rect 2990 4548 2994 4552
rect 2998 4548 3002 4552
rect 3054 4548 3058 4552
rect 3486 4548 3490 4552
rect 4006 4548 4010 4552
rect 4430 4548 4434 4552
rect 4486 4548 4490 4552
rect 4494 4548 4498 4552
rect 734 4538 738 4542
rect 758 4538 762 4542
rect 982 4538 986 4542
rect 1382 4538 1386 4542
rect 1614 4538 1618 4542
rect 1638 4538 1642 4542
rect 1974 4538 1978 4542
rect 2182 4538 2186 4542
rect 2254 4538 2258 4542
rect 2502 4538 2506 4542
rect 2534 4538 2538 4542
rect 2678 4538 2682 4542
rect 2966 4538 2970 4542
rect 2990 4538 2994 4542
rect 3078 4538 3082 4542
rect 3526 4538 3530 4542
rect 3590 4538 3594 4542
rect 3678 4538 3682 4542
rect 4062 4538 4066 4542
rect 4278 4538 4282 4542
rect 4398 4538 4402 4542
rect 4510 4538 4514 4542
rect 4526 4538 4530 4542
rect 4750 4538 4754 4542
rect 5158 4538 5162 4542
rect 854 4528 858 4532
rect 1574 4528 1578 4532
rect 1606 4528 1610 4532
rect 1710 4528 1714 4532
rect 1910 4528 1914 4532
rect 1982 4528 1986 4532
rect 2214 4528 2218 4532
rect 2526 4528 2530 4532
rect 2982 4528 2986 4532
rect 3534 4528 3538 4532
rect 3894 4528 3898 4532
rect 4094 4528 4098 4532
rect 4558 4528 4562 4532
rect 4870 4528 4874 4532
rect 4942 4528 4946 4532
rect 582 4518 586 4522
rect 686 4518 690 4522
rect 998 4518 1002 4522
rect 1214 4518 1218 4522
rect 1622 4518 1626 4522
rect 1926 4518 1930 4522
rect 2230 4518 2234 4522
rect 3886 4518 3890 4522
rect 4350 4518 4354 4522
rect 4406 4518 4410 4522
rect 822 4508 826 4512
rect 1630 4508 1634 4512
rect 1774 4508 1778 4512
rect 2270 4508 2274 4512
rect 2566 4508 2570 4512
rect 2694 4508 2698 4512
rect 3014 4508 3018 4512
rect 3086 4508 3090 4512
rect 3382 4508 3386 4512
rect 3526 4508 3530 4512
rect 3550 4508 3554 4512
rect 4158 4508 4162 4512
rect 4710 4508 4714 4512
rect 1050 4503 1054 4507
rect 1058 4503 1061 4507
rect 1061 4503 1062 4507
rect 2074 4503 2078 4507
rect 2082 4503 2085 4507
rect 2085 4503 2086 4507
rect 3098 4503 3102 4507
rect 3106 4503 3109 4507
rect 3109 4503 3110 4507
rect 4114 4503 4118 4507
rect 4122 4503 4125 4507
rect 4125 4503 4126 4507
rect 1758 4498 1762 4502
rect 2246 4498 2250 4502
rect 2398 4498 2402 4502
rect 3966 4498 3970 4502
rect 5182 4498 5186 4502
rect 1070 4488 1074 4492
rect 1766 4488 1770 4492
rect 2478 4488 2482 4492
rect 2726 4488 2730 4492
rect 2750 4488 2754 4492
rect 3518 4488 3522 4492
rect 3542 4488 3546 4492
rect 3950 4488 3954 4492
rect 4142 4488 4146 4492
rect 4454 4488 4458 4492
rect 110 4478 114 4482
rect 1310 4478 1314 4482
rect 1886 4478 1890 4482
rect 2310 4478 2314 4482
rect 2678 4478 2682 4482
rect 3406 4478 3410 4482
rect 5038 4478 5042 4482
rect 1150 4468 1154 4472
rect 1190 4468 1194 4472
rect 1334 4468 1338 4472
rect 1422 4468 1426 4472
rect 1598 4468 1602 4472
rect 1854 4468 1858 4472
rect 1918 4468 1922 4472
rect 2238 4468 2242 4472
rect 2270 4468 2274 4472
rect 2302 4468 2306 4472
rect 2422 4468 2426 4472
rect 2702 4468 2706 4472
rect 2718 4468 2722 4472
rect 2974 4468 2978 4472
rect 3198 4468 3202 4472
rect 3806 4468 3810 4472
rect 4438 4468 4442 4472
rect 4662 4468 4666 4472
rect 4918 4468 4922 4472
rect 246 4458 250 4462
rect 710 4458 714 4462
rect 726 4458 730 4462
rect 1158 4458 1162 4462
rect 1454 4458 1458 4462
rect 1494 4458 1498 4462
rect 1510 4458 1514 4462
rect 1590 4458 1594 4462
rect 1622 4458 1626 4462
rect 1854 4458 1858 4462
rect 2030 4458 2034 4462
rect 2270 4458 2274 4462
rect 2366 4458 2370 4462
rect 2406 4458 2410 4462
rect 2734 4458 2738 4462
rect 3030 4458 3034 4462
rect 3134 4458 3138 4462
rect 3262 4458 3266 4462
rect 3862 4458 3866 4462
rect 3902 4458 3906 4462
rect 4022 4458 4026 4462
rect 4078 4458 4082 4462
rect 4326 4458 4330 4462
rect 4430 4458 4434 4462
rect 4758 4458 4762 4462
rect 4814 4458 4818 4462
rect 5054 4458 5058 4462
rect 1238 4448 1242 4452
rect 1894 4448 1898 4452
rect 2030 4448 2034 4452
rect 2062 4448 2066 4452
rect 2294 4448 2298 4452
rect 2382 4448 2386 4452
rect 2886 4448 2890 4452
rect 2974 4448 2978 4452
rect 4814 4448 4818 4452
rect 934 4438 938 4442
rect 990 4438 994 4442
rect 1558 4438 1562 4442
rect 1958 4438 1962 4442
rect 3566 4438 3570 4442
rect 3886 4438 3890 4442
rect 4134 4438 4138 4442
rect 4326 4438 4330 4442
rect 4502 4438 4506 4442
rect 4582 4438 4586 4442
rect 2494 4428 2498 4432
rect 1558 4418 1562 4422
rect 1838 4418 1842 4422
rect 2526 4418 2530 4422
rect 3238 4418 3242 4422
rect 102 4408 106 4412
rect 590 4408 594 4412
rect 1270 4408 1274 4412
rect 3510 4408 3514 4412
rect 3822 4408 3826 4412
rect 3982 4408 3986 4412
rect 4270 4408 4274 4412
rect 4534 4408 4538 4412
rect 4830 4408 4834 4412
rect 538 4403 542 4407
rect 546 4403 549 4407
rect 549 4403 550 4407
rect 1562 4403 1566 4407
rect 1570 4403 1573 4407
rect 1573 4403 1574 4407
rect 2586 4403 2590 4407
rect 2594 4403 2597 4407
rect 2597 4403 2598 4407
rect 3610 4403 3614 4407
rect 3618 4403 3621 4407
rect 3621 4403 3622 4407
rect 4634 4403 4638 4407
rect 4642 4403 4645 4407
rect 4645 4403 4646 4407
rect 1094 4398 1098 4402
rect 1222 4398 1226 4402
rect 2246 4398 2250 4402
rect 2262 4398 2266 4402
rect 3150 4398 3154 4402
rect 3206 4398 3210 4402
rect 3214 4398 3218 4402
rect 1222 4388 1226 4392
rect 2302 4388 2306 4392
rect 3646 4388 3650 4392
rect 3710 4388 3714 4392
rect 4150 4388 4154 4392
rect 4358 4388 4362 4392
rect 1030 4378 1034 4382
rect 1806 4378 1810 4382
rect 1926 4378 1930 4382
rect 1998 4378 2002 4382
rect 2534 4378 2538 4382
rect 3750 4378 3754 4382
rect 4222 4378 4226 4382
rect 4510 4378 4514 4382
rect 4918 4378 4922 4382
rect 94 4368 98 4372
rect 286 4368 290 4372
rect 1598 4368 1602 4372
rect 1902 4368 1906 4372
rect 2366 4368 2370 4372
rect 2702 4368 2706 4372
rect 2726 4368 2730 4372
rect 3494 4368 3498 4372
rect 3758 4368 3762 4372
rect 4206 4368 4210 4372
rect 4422 4368 4426 4372
rect 4430 4368 4434 4372
rect 294 4358 298 4362
rect 998 4358 1002 4362
rect 1582 4358 1586 4362
rect 2262 4358 2266 4362
rect 2278 4358 2282 4362
rect 2286 4358 2290 4362
rect 2478 4358 2482 4362
rect 2534 4358 2538 4362
rect 3558 4358 3562 4362
rect 3966 4358 3970 4362
rect 4702 4358 4706 4362
rect 4870 4358 4874 4362
rect 246 4348 250 4352
rect 270 4348 274 4352
rect 1446 4348 1450 4352
rect 2406 4348 2410 4352
rect 2750 4348 2754 4352
rect 2774 4348 2778 4352
rect 2798 4348 2802 4352
rect 3150 4348 3154 4352
rect 3174 4348 3178 4352
rect 3670 4348 3674 4352
rect 3782 4348 3786 4352
rect 3958 4348 3962 4352
rect 4078 4348 4082 4352
rect 4310 4348 4314 4352
rect 4334 4348 4338 4352
rect 4446 4348 4450 4352
rect 4590 4348 4594 4352
rect 262 4338 266 4342
rect 350 4338 354 4342
rect 630 4338 634 4342
rect 854 4338 858 4342
rect 1006 4338 1010 4342
rect 1118 4328 1122 4332
rect 1550 4328 1554 4332
rect 2174 4338 2178 4342
rect 2190 4338 2194 4342
rect 2550 4338 2554 4342
rect 2798 4338 2802 4342
rect 2878 4338 2882 4342
rect 2886 4338 2890 4342
rect 3486 4338 3490 4342
rect 3774 4338 3778 4342
rect 3934 4338 3938 4342
rect 4030 4338 4034 4342
rect 4294 4338 4298 4342
rect 4558 4338 4562 4342
rect 4694 4338 4698 4342
rect 2446 4328 2450 4332
rect 2646 4328 2650 4332
rect 2782 4328 2786 4332
rect 2966 4328 2970 4332
rect 3326 4328 3330 4332
rect 3422 4328 3426 4332
rect 3846 4328 3850 4332
rect 3958 4328 3962 4332
rect 142 4318 146 4322
rect 862 4318 866 4322
rect 1694 4318 1698 4322
rect 2342 4318 2346 4322
rect 2502 4318 2506 4322
rect 4014 4318 4018 4322
rect 4150 4318 4154 4322
rect 4230 4318 4234 4322
rect 4350 4318 4354 4322
rect 582 4308 586 4312
rect 1910 4308 1914 4312
rect 3462 4308 3466 4312
rect 3998 4308 4002 4312
rect 4102 4308 4106 4312
rect 4134 4308 4138 4312
rect 4502 4308 4506 4312
rect 4870 4308 4874 4312
rect 1050 4303 1054 4307
rect 1058 4303 1061 4307
rect 1061 4303 1062 4307
rect 2074 4303 2078 4307
rect 2082 4303 2085 4307
rect 2085 4303 2086 4307
rect 3098 4303 3102 4307
rect 3106 4303 3109 4307
rect 3109 4303 3110 4307
rect 4114 4303 4118 4307
rect 4122 4303 4125 4307
rect 4125 4303 4126 4307
rect 926 4298 930 4302
rect 1230 4298 1234 4302
rect 1462 4298 1466 4302
rect 2606 4298 2610 4302
rect 2630 4298 2634 4302
rect 2830 4298 2834 4302
rect 2838 4298 2842 4302
rect 3326 4298 3330 4302
rect 3886 4298 3890 4302
rect 3934 4298 3938 4302
rect 4046 4298 4050 4302
rect 4134 4298 4138 4302
rect 4710 4298 4714 4302
rect 774 4288 778 4292
rect 1622 4288 1626 4292
rect 1750 4288 1754 4292
rect 2206 4288 2210 4292
rect 2222 4288 2226 4292
rect 2710 4288 2714 4292
rect 2846 4288 2850 4292
rect 3126 4288 3130 4292
rect 3470 4288 3474 4292
rect 3526 4288 3530 4292
rect 4246 4288 4250 4292
rect 1166 4278 1170 4282
rect 1326 4278 1330 4282
rect 1782 4278 1786 4282
rect 2142 4278 2146 4282
rect 2430 4278 2434 4282
rect 3222 4278 3226 4282
rect 3558 4278 3562 4282
rect 4246 4278 4250 4282
rect 334 4268 338 4272
rect 430 4268 434 4272
rect 638 4268 642 4272
rect 782 4268 786 4272
rect 878 4268 882 4272
rect 966 4268 970 4272
rect 1006 4268 1010 4272
rect 1070 4268 1074 4272
rect 1166 4268 1170 4272
rect 1542 4268 1546 4272
rect 1726 4268 1730 4272
rect 2150 4268 2154 4272
rect 2350 4268 2354 4272
rect 2438 4268 2442 4272
rect 2742 4268 2746 4272
rect 3150 4268 3154 4272
rect 3782 4268 3786 4272
rect 3870 4268 3874 4272
rect 3878 4268 3882 4272
rect 3918 4268 3922 4272
rect 3942 4268 3946 4272
rect 4038 4268 4042 4272
rect 4046 4268 4050 4272
rect 4238 4268 4242 4272
rect 4262 4268 4266 4272
rect 4902 4268 4906 4272
rect 5062 4268 5066 4272
rect 110 4258 114 4262
rect 550 4258 554 4262
rect 806 4258 810 4262
rect 1014 4258 1018 4262
rect 1206 4258 1210 4262
rect 1734 4258 1738 4262
rect 1822 4258 1826 4262
rect 2038 4258 2042 4262
rect 2286 4258 2290 4262
rect 2342 4258 2346 4262
rect 2374 4258 2378 4262
rect 2670 4258 2674 4262
rect 2750 4258 2754 4262
rect 2918 4258 2922 4262
rect 2958 4258 2962 4262
rect 3142 4258 3146 4262
rect 3182 4258 3186 4262
rect 3430 4258 3434 4262
rect 3534 4258 3538 4262
rect 1006 4248 1010 4252
rect 1166 4248 1170 4252
rect 3806 4258 3810 4262
rect 3870 4258 3874 4262
rect 4022 4258 4026 4262
rect 4038 4258 4042 4262
rect 4310 4258 4314 4262
rect 4430 4258 4434 4262
rect 4606 4258 4610 4262
rect 4670 4258 4674 4262
rect 1814 4248 1818 4252
rect 1838 4248 1842 4252
rect 2182 4248 2186 4252
rect 2302 4248 2306 4252
rect 2310 4248 2314 4252
rect 2382 4248 2386 4252
rect 3150 4248 3154 4252
rect 3598 4248 3602 4252
rect 3638 4248 3642 4252
rect 3742 4248 3746 4252
rect 3870 4248 3874 4252
rect 590 4238 594 4242
rect 1614 4238 1618 4242
rect 2926 4238 2930 4242
rect 3718 4238 3722 4242
rect 3798 4238 3802 4242
rect 3886 4238 3890 4242
rect 4230 4248 4234 4252
rect 4558 4248 4562 4252
rect 4814 4238 4818 4242
rect 446 4228 450 4232
rect 702 4228 706 4232
rect 1078 4228 1082 4232
rect 1686 4228 1690 4232
rect 1990 4228 1994 4232
rect 3078 4228 3082 4232
rect 4006 4228 4010 4232
rect 4430 4228 4434 4232
rect 134 4218 138 4222
rect 670 4218 674 4222
rect 1430 4218 1434 4222
rect 2454 4218 2458 4222
rect 3422 4218 3426 4222
rect 4622 4218 4626 4222
rect 1406 4208 1410 4212
rect 1750 4208 1754 4212
rect 2102 4208 2106 4212
rect 2510 4208 2514 4212
rect 2966 4208 2970 4212
rect 4214 4208 4218 4212
rect 538 4203 542 4207
rect 546 4203 549 4207
rect 549 4203 550 4207
rect 1562 4203 1566 4207
rect 1570 4203 1573 4207
rect 1573 4203 1574 4207
rect 2586 4203 2590 4207
rect 2594 4203 2597 4207
rect 2597 4203 2598 4207
rect 3610 4203 3614 4207
rect 3618 4203 3621 4207
rect 3621 4203 3622 4207
rect 4634 4203 4638 4207
rect 4642 4203 4645 4207
rect 4645 4203 4646 4207
rect 886 4198 890 4202
rect 974 4198 978 4202
rect 1638 4198 1642 4202
rect 1870 4198 1874 4202
rect 2366 4198 2370 4202
rect 2606 4198 2610 4202
rect 2694 4198 2698 4202
rect 3598 4198 3602 4202
rect 3782 4198 3786 4202
rect 3814 4198 3818 4202
rect 4598 4198 4602 4202
rect 262 4188 266 4192
rect 1126 4188 1130 4192
rect 1974 4188 1978 4192
rect 2374 4188 2378 4192
rect 2390 4188 2394 4192
rect 2870 4188 2874 4192
rect 3134 4188 3138 4192
rect 4214 4188 4218 4192
rect 4454 4188 4458 4192
rect 358 4178 362 4182
rect 518 4178 522 4182
rect 718 4178 722 4182
rect 1910 4178 1914 4182
rect 3398 4178 3402 4182
rect 3406 4178 3410 4182
rect 3526 4178 3530 4182
rect 3542 4178 3546 4182
rect 3822 4178 3826 4182
rect 3990 4178 3994 4182
rect 382 4168 386 4172
rect 2198 4168 2202 4172
rect 2318 4168 2322 4172
rect 2326 4168 2330 4172
rect 2910 4168 2914 4172
rect 2926 4168 2930 4172
rect 4374 4168 4378 4172
rect 254 4158 258 4162
rect 926 4158 930 4162
rect 998 4158 1002 4162
rect 1526 4158 1530 4162
rect 1862 4158 1866 4162
rect 2366 4158 2370 4162
rect 2430 4158 2434 4162
rect 3254 4158 3258 4162
rect 3478 4158 3482 4162
rect 3638 4158 3642 4162
rect 4174 4158 4178 4162
rect 4654 4158 4658 4162
rect 4694 4158 4698 4162
rect 302 4148 306 4152
rect 366 4148 370 4152
rect 422 4148 426 4152
rect 798 4148 802 4152
rect 1006 4148 1010 4152
rect 1022 4148 1026 4152
rect 1358 4148 1362 4152
rect 1710 4148 1714 4152
rect 1734 4148 1738 4152
rect 2166 4148 2170 4152
rect 2286 4148 2290 4152
rect 2318 4148 2322 4152
rect 2422 4148 2426 4152
rect 2470 4148 2474 4152
rect 2726 4148 2730 4152
rect 2798 4148 2802 4152
rect 2950 4148 2954 4152
rect 2966 4148 2970 4152
rect 3214 4148 3218 4152
rect 3246 4148 3250 4152
rect 3430 4148 3434 4152
rect 3558 4148 3562 4152
rect 3598 4148 3602 4152
rect 4078 4148 4082 4152
rect 278 4138 282 4142
rect 318 4138 322 4142
rect 342 4138 346 4142
rect 430 4138 434 4142
rect 894 4138 898 4142
rect 998 4138 1002 4142
rect 1038 4138 1042 4142
rect 1182 4138 1186 4142
rect 1230 4138 1234 4142
rect 1310 4138 1314 4142
rect 1494 4138 1498 4142
rect 1638 4138 1642 4142
rect 4526 4148 4530 4152
rect 4630 4148 4634 4152
rect 4942 4148 4946 4152
rect 5054 4148 5058 4152
rect 1718 4138 1722 4142
rect 1966 4138 1970 4142
rect 2334 4138 2338 4142
rect 2446 4138 2450 4142
rect 2814 4138 2818 4142
rect 2822 4138 2826 4142
rect 3238 4138 3242 4142
rect 3270 4138 3274 4142
rect 3598 4138 3602 4142
rect 3750 4138 3754 4142
rect 3974 4138 3978 4142
rect 3998 4138 4002 4142
rect 4094 4138 4098 4142
rect 4246 4138 4250 4142
rect 4286 4138 4290 4142
rect 4478 4138 4482 4142
rect 4542 4138 4546 4142
rect 4550 4138 4554 4142
rect 4710 4138 4714 4142
rect 4734 4138 4738 4142
rect 390 4128 394 4132
rect 598 4128 602 4132
rect 1006 4128 1010 4132
rect 1310 4128 1314 4132
rect 1518 4128 1522 4132
rect 1718 4128 1722 4132
rect 2142 4128 2146 4132
rect 2750 4128 2754 4132
rect 2846 4128 2850 4132
rect 3478 4128 3482 4132
rect 3766 4128 3770 4132
rect 3990 4128 3994 4132
rect 966 4118 970 4122
rect 1286 4118 1290 4122
rect 1366 4118 1370 4122
rect 1750 4118 1754 4122
rect 2894 4118 2898 4122
rect 3502 4118 3506 4122
rect 3902 4118 3906 4122
rect 4446 4118 4450 4122
rect 4566 4118 4570 4122
rect 1214 4108 1218 4112
rect 1294 4108 1298 4112
rect 1702 4108 1706 4112
rect 2806 4108 2810 4112
rect 3214 4108 3218 4112
rect 3398 4108 3402 4112
rect 3582 4108 3586 4112
rect 3934 4108 3938 4112
rect 4086 4108 4090 4112
rect 1050 4103 1054 4107
rect 1058 4103 1061 4107
rect 1061 4103 1062 4107
rect 2074 4103 2078 4107
rect 2082 4103 2085 4107
rect 2085 4103 2086 4107
rect 3098 4103 3102 4107
rect 3106 4103 3109 4107
rect 3109 4103 3110 4107
rect 4114 4103 4118 4107
rect 4122 4103 4125 4107
rect 4125 4103 4126 4107
rect 486 4098 490 4102
rect 1038 4098 1042 4102
rect 1998 4098 2002 4102
rect 2222 4098 2226 4102
rect 2262 4098 2266 4102
rect 2302 4098 2306 4102
rect 2310 4098 2314 4102
rect 2702 4098 2706 4102
rect 2790 4098 2794 4102
rect 2830 4098 2834 4102
rect 3550 4098 3554 4102
rect 3574 4098 3578 4102
rect 4654 4098 4658 4102
rect 5062 4098 5066 4102
rect 1206 4088 1210 4092
rect 1374 4088 1378 4092
rect 1398 4088 1402 4092
rect 1806 4088 1810 4092
rect 2526 4088 2530 4092
rect 2638 4088 2642 4092
rect 3030 4088 3034 4092
rect 3198 4088 3202 4092
rect 3222 4088 3226 4092
rect 3526 4088 3530 4092
rect 3950 4088 3954 4092
rect 4262 4088 4266 4092
rect 4270 4088 4274 4092
rect 502 4078 506 4082
rect 1342 4078 1346 4082
rect 1486 4078 1490 4082
rect 1726 4078 1730 4082
rect 1982 4078 1986 4082
rect 2046 4078 2050 4082
rect 2350 4078 2354 4082
rect 2422 4078 2426 4082
rect 3222 4078 3226 4082
rect 3230 4078 3234 4082
rect 3742 4078 3746 4082
rect 3942 4078 3946 4082
rect 4590 4078 4594 4082
rect 4742 4078 4746 4082
rect 494 4068 498 4072
rect 518 4068 522 4072
rect 574 4068 578 4072
rect 606 4068 610 4072
rect 662 4068 666 4072
rect 790 4068 794 4072
rect 926 4068 930 4072
rect 958 4068 962 4072
rect 1046 4068 1050 4072
rect 1150 4068 1154 4072
rect 1534 4068 1538 4072
rect 1902 4068 1906 4072
rect 1934 4068 1938 4072
rect 2518 4068 2522 4072
rect 2606 4068 2610 4072
rect 2758 4068 2762 4072
rect 2934 4068 2938 4072
rect 102 4058 106 4062
rect 310 4058 314 4062
rect 334 4058 338 4062
rect 382 4058 386 4062
rect 582 4058 586 4062
rect 870 4058 874 4062
rect 918 4058 922 4062
rect 942 4058 946 4062
rect 1222 4058 1226 4062
rect 1238 4058 1242 4062
rect 1414 4058 1418 4062
rect 3446 4068 3450 4072
rect 3510 4068 3514 4072
rect 3558 4068 3562 4072
rect 3758 4068 3762 4072
rect 3782 4068 3786 4072
rect 3990 4068 3994 4072
rect 4006 4068 4010 4072
rect 4038 4068 4042 4072
rect 4230 4068 4234 4072
rect 4270 4068 4274 4072
rect 4310 4068 4314 4072
rect 4342 4068 4346 4072
rect 1526 4058 1530 4062
rect 1614 4058 1618 4062
rect 1694 4058 1698 4062
rect 1766 4058 1770 4062
rect 1830 4058 1834 4062
rect 1894 4058 1898 4062
rect 2350 4058 2354 4062
rect 2358 4058 2362 4062
rect 2390 4058 2394 4062
rect 2438 4058 2442 4062
rect 2470 4058 2474 4062
rect 2822 4058 2826 4062
rect 3198 4058 3202 4062
rect 3414 4058 3418 4062
rect 3486 4058 3490 4062
rect 3550 4058 3554 4062
rect 3630 4058 3634 4062
rect 3726 4058 3730 4062
rect 3758 4058 3762 4062
rect 3790 4058 3794 4062
rect 3806 4058 3810 4062
rect 3950 4058 3954 4062
rect 4054 4058 4058 4062
rect 4246 4058 4250 4062
rect 4262 4058 4266 4062
rect 4358 4058 4362 4062
rect 4422 4058 4426 4062
rect 334 4048 338 4052
rect 902 4048 906 4052
rect 1070 4048 1074 4052
rect 1534 4048 1538 4052
rect 1934 4048 1938 4052
rect 2206 4048 2210 4052
rect 2454 4048 2458 4052
rect 2574 4048 2578 4052
rect 2654 4048 2658 4052
rect 2710 4048 2714 4052
rect 3070 4048 3074 4052
rect 3326 4048 3330 4052
rect 4174 4048 4178 4052
rect 4286 4048 4290 4052
rect 4678 4048 4682 4052
rect 382 4038 386 4042
rect 510 4038 514 4042
rect 734 4038 738 4042
rect 878 4038 882 4042
rect 966 4038 970 4042
rect 1230 4038 1234 4042
rect 1310 4038 1314 4042
rect 1542 4038 1546 4042
rect 2142 4038 2146 4042
rect 3470 4038 3474 4042
rect 3638 4038 3642 4042
rect 4046 4038 4050 4042
rect 4094 4038 4098 4042
rect 4430 4038 4434 4042
rect 4870 4038 4874 4042
rect 630 4028 634 4032
rect 814 4028 818 4032
rect 1222 4028 1226 4032
rect 1654 4028 1658 4032
rect 1886 4028 1890 4032
rect 1910 4028 1914 4032
rect 2662 4028 2666 4032
rect 910 4018 914 4022
rect 1022 4018 1026 4022
rect 1622 4018 1626 4022
rect 2054 4018 2058 4022
rect 2142 4018 2146 4022
rect 2606 4018 2610 4022
rect 3670 4028 3674 4032
rect 3950 4028 3954 4032
rect 4022 4028 4026 4032
rect 4446 4028 4450 4032
rect 2838 4018 2842 4022
rect 2846 4018 2850 4022
rect 3006 4018 3010 4022
rect 3502 4018 3506 4022
rect 3750 4018 3754 4022
rect 142 4008 146 4012
rect 486 4008 490 4012
rect 1270 4008 1274 4012
rect 2206 4008 2210 4012
rect 2550 4008 2554 4012
rect 2958 4008 2962 4012
rect 3398 4008 3402 4012
rect 3486 4008 3490 4012
rect 3686 4008 3690 4012
rect 4518 4008 4522 4012
rect 538 4003 542 4007
rect 546 4003 549 4007
rect 549 4003 550 4007
rect 1562 4003 1566 4007
rect 1570 4003 1573 4007
rect 1573 4003 1574 4007
rect 2586 4003 2590 4007
rect 2594 4003 2597 4007
rect 2597 4003 2598 4007
rect 3610 4003 3614 4007
rect 3618 4003 3621 4007
rect 3621 4003 3622 4007
rect 4634 4003 4638 4007
rect 4642 4003 4645 4007
rect 4645 4003 4646 4007
rect 1142 3998 1146 4002
rect 2654 3998 2658 4002
rect 3974 3998 3978 4002
rect 4286 3998 4290 4002
rect 4654 3998 4658 4002
rect 1726 3988 1730 3992
rect 1926 3988 1930 3992
rect 2366 3988 2370 3992
rect 2806 3988 2810 3992
rect 4006 3988 4010 3992
rect 4294 3988 4298 3992
rect 358 3978 362 3982
rect 590 3978 594 3982
rect 1014 3978 1018 3982
rect 1142 3978 1146 3982
rect 1198 3978 1202 3982
rect 1246 3978 1250 3982
rect 1502 3978 1506 3982
rect 1926 3978 1930 3982
rect 3214 3978 3218 3982
rect 3998 3978 4002 3982
rect 4214 3978 4218 3982
rect 4502 3978 4506 3982
rect 950 3968 954 3972
rect 1014 3968 1018 3972
rect 1038 3968 1042 3972
rect 1150 3968 1154 3972
rect 1174 3968 1178 3972
rect 1206 3968 1210 3972
rect 1518 3968 1522 3972
rect 1550 3968 1554 3972
rect 2158 3968 2162 3972
rect 2606 3968 2610 3972
rect 2758 3968 2762 3972
rect 3518 3968 3522 3972
rect 4102 3968 4106 3972
rect 4302 3968 4306 3972
rect 4918 3968 4922 3972
rect 94 3958 98 3962
rect 406 3958 410 3962
rect 590 3958 594 3962
rect 1278 3958 1282 3962
rect 1342 3958 1346 3962
rect 1742 3958 1746 3962
rect 1774 3958 1778 3962
rect 1806 3958 1810 3962
rect 1862 3958 1866 3962
rect 2166 3958 2170 3962
rect 2398 3958 2402 3962
rect 2838 3958 2842 3962
rect 2886 3958 2890 3962
rect 3766 3958 3770 3962
rect 3846 3958 3850 3962
rect 4142 3958 4146 3962
rect 4230 3958 4234 3962
rect 4390 3958 4394 3962
rect 134 3948 138 3952
rect 174 3948 178 3952
rect 734 3948 738 3952
rect 942 3948 946 3952
rect 1038 3948 1042 3952
rect 1054 3948 1058 3952
rect 1078 3948 1082 3952
rect 1838 3948 1842 3952
rect 2038 3948 2042 3952
rect 2182 3948 2186 3952
rect 2766 3948 2770 3952
rect 2982 3948 2986 3952
rect 3038 3948 3042 3952
rect 3254 3948 3258 3952
rect 4174 3948 4178 3952
rect 4222 3948 4226 3952
rect 4326 3948 4330 3952
rect 4390 3948 4394 3952
rect 4446 3948 4450 3952
rect 4454 3948 4458 3952
rect 4550 3948 4554 3952
rect 4654 3948 4658 3952
rect 166 3938 170 3942
rect 326 3938 330 3942
rect 710 3938 714 3942
rect 862 3938 866 3942
rect 1182 3938 1186 3942
rect 1486 3938 1490 3942
rect 1558 3938 1562 3942
rect 1814 3938 1818 3942
rect 2014 3938 2018 3942
rect 2118 3938 2122 3942
rect 2366 3938 2370 3942
rect 2630 3938 2634 3942
rect 3014 3938 3018 3942
rect 3342 3938 3346 3942
rect 3462 3938 3466 3942
rect 3934 3938 3938 3942
rect 4398 3938 4402 3942
rect 4694 3938 4698 3942
rect 4766 3938 4770 3942
rect 4902 3938 4906 3942
rect 438 3928 442 3932
rect 1078 3928 1082 3932
rect 1214 3928 1218 3932
rect 1374 3928 1378 3932
rect 1462 3928 1466 3932
rect 1662 3928 1666 3932
rect 2190 3928 2194 3932
rect 2822 3928 2826 3932
rect 2878 3928 2882 3932
rect 2902 3928 2906 3932
rect 3390 3928 3394 3932
rect 3414 3928 3418 3932
rect 3838 3928 3842 3932
rect 3854 3928 3858 3932
rect 4254 3928 4258 3932
rect 4582 3928 4586 3932
rect 4678 3928 4682 3932
rect 1766 3918 1770 3922
rect 2022 3918 2026 3922
rect 2334 3918 2338 3922
rect 2678 3918 2682 3922
rect 2854 3918 2858 3922
rect 3894 3918 3898 3922
rect 4070 3918 4074 3922
rect 4182 3918 4186 3922
rect 4206 3918 4210 3922
rect 4270 3918 4274 3922
rect 4358 3918 4362 3922
rect 126 3908 130 3912
rect 1334 3908 1338 3912
rect 1606 3908 1610 3912
rect 1702 3908 1706 3912
rect 1790 3908 1794 3912
rect 2214 3908 2218 3912
rect 2526 3908 2530 3912
rect 2806 3908 2810 3912
rect 3022 3908 3026 3912
rect 3374 3908 3378 3912
rect 1050 3903 1054 3907
rect 1058 3903 1061 3907
rect 1061 3903 1062 3907
rect 2074 3903 2078 3907
rect 2082 3903 2085 3907
rect 2085 3903 2086 3907
rect 3098 3903 3102 3907
rect 3106 3903 3109 3907
rect 3109 3903 3110 3907
rect 4114 3903 4118 3907
rect 4122 3903 4125 3907
rect 4125 3903 4126 3907
rect 958 3898 962 3902
rect 1798 3898 1802 3902
rect 4374 3898 4378 3902
rect 4558 3898 4562 3902
rect 1102 3888 1106 3892
rect 2062 3888 2066 3892
rect 3678 3888 3682 3892
rect 4454 3888 4458 3892
rect 4814 3888 4818 3892
rect 414 3878 418 3882
rect 910 3878 914 3882
rect 1742 3878 1746 3882
rect 1870 3878 1874 3882
rect 2262 3878 2266 3882
rect 2326 3878 2330 3882
rect 2422 3878 2426 3882
rect 3438 3878 3442 3882
rect 4166 3878 4170 3882
rect 4246 3878 4250 3882
rect 4262 3878 4266 3882
rect 4574 3878 4578 3882
rect 4918 3878 4922 3882
rect 430 3868 434 3872
rect 974 3868 978 3872
rect 1022 3868 1026 3872
rect 1094 3868 1098 3872
rect 1150 3868 1154 3872
rect 1158 3868 1162 3872
rect 1414 3868 1418 3872
rect 1446 3868 1450 3872
rect 1574 3868 1578 3872
rect 1878 3868 1882 3872
rect 2342 3868 2346 3872
rect 2782 3868 2786 3872
rect 3046 3868 3050 3872
rect 3070 3868 3074 3872
rect 3262 3868 3266 3872
rect 3382 3868 3386 3872
rect 3542 3868 3546 3872
rect 3606 3868 3610 3872
rect 3750 3868 3754 3872
rect 4054 3868 4058 3872
rect 4230 3868 4234 3872
rect 4270 3868 4274 3872
rect 4318 3868 4322 3872
rect 4374 3868 4378 3872
rect 270 3858 274 3862
rect 766 3858 770 3862
rect 822 3858 826 3862
rect 1070 3858 1074 3862
rect 1478 3858 1482 3862
rect 1526 3858 1530 3862
rect 1550 3858 1554 3862
rect 1590 3858 1594 3862
rect 1782 3858 1786 3862
rect 2126 3858 2130 3862
rect 2158 3858 2162 3862
rect 2198 3858 2202 3862
rect 2430 3858 2434 3862
rect 2558 3858 2562 3862
rect 2598 3858 2602 3862
rect 2622 3858 2626 3862
rect 2726 3858 2730 3862
rect 2774 3858 2778 3862
rect 2942 3858 2946 3862
rect 2958 3858 2962 3862
rect 2998 3858 3002 3862
rect 3078 3858 3082 3862
rect 3294 3858 3298 3862
rect 3334 3858 3338 3862
rect 3366 3858 3370 3862
rect 4134 3858 4138 3862
rect 4286 3858 4290 3862
rect 4398 3858 4402 3862
rect 4438 3858 4442 3862
rect 4470 3858 4474 3862
rect 4526 3858 4530 3862
rect 5078 3858 5082 3862
rect 1078 3848 1082 3852
rect 1334 3848 1338 3852
rect 2398 3848 2402 3852
rect 2422 3848 2426 3852
rect 3214 3848 3218 3852
rect 3238 3848 3242 3852
rect 3342 3848 3346 3852
rect 3654 3848 3658 3852
rect 3678 3848 3682 3852
rect 3774 3848 3778 3852
rect 3942 3848 3946 3852
rect 4918 3848 4922 3852
rect 5054 3848 5058 3852
rect 1118 3838 1122 3842
rect 1814 3838 1818 3842
rect 2038 3838 2042 3842
rect 2870 3838 2874 3842
rect 3494 3838 3498 3842
rect 4262 3838 4266 3842
rect 4414 3838 4418 3842
rect 4542 3838 4546 3842
rect 1430 3828 1434 3832
rect 2302 3828 2306 3832
rect 2542 3828 2546 3832
rect 2718 3828 2722 3832
rect 2918 3828 2922 3832
rect 2942 3828 2946 3832
rect 3398 3828 3402 3832
rect 3494 3828 3498 3832
rect 4398 3828 4402 3832
rect 5054 3828 5058 3832
rect 358 3818 362 3822
rect 806 3818 810 3822
rect 1862 3818 1866 3822
rect 2334 3818 2338 3822
rect 2374 3818 2378 3822
rect 2686 3818 2690 3822
rect 3718 3818 3722 3822
rect 3894 3818 3898 3822
rect 4462 3818 4466 3822
rect 526 3808 530 3812
rect 1206 3808 1210 3812
rect 1534 3808 1538 3812
rect 1582 3808 1586 3812
rect 2110 3808 2114 3812
rect 2310 3808 2314 3812
rect 2374 3808 2378 3812
rect 2414 3808 2418 3812
rect 2542 3808 2546 3812
rect 2950 3808 2954 3812
rect 4422 3808 4426 3812
rect 4486 3808 4490 3812
rect 538 3803 542 3807
rect 546 3803 549 3807
rect 549 3803 550 3807
rect 1562 3803 1566 3807
rect 1570 3803 1573 3807
rect 1573 3803 1574 3807
rect 2586 3803 2590 3807
rect 2594 3803 2597 3807
rect 2597 3803 2598 3807
rect 3610 3803 3614 3807
rect 3618 3803 3621 3807
rect 3621 3803 3622 3807
rect 4634 3803 4638 3807
rect 4642 3803 4645 3807
rect 4645 3803 4646 3807
rect 1166 3798 1170 3802
rect 1862 3798 1866 3802
rect 2798 3798 2802 3802
rect 3710 3798 3714 3802
rect 4198 3798 4202 3802
rect 1486 3788 1490 3792
rect 1894 3788 1898 3792
rect 2278 3788 2282 3792
rect 2390 3788 2394 3792
rect 2806 3788 2810 3792
rect 2966 3788 2970 3792
rect 4734 3788 4738 3792
rect 526 3778 530 3782
rect 838 3778 842 3782
rect 1078 3778 1082 3782
rect 1350 3778 1354 3782
rect 1782 3778 1786 3782
rect 2662 3778 2666 3782
rect 2998 3778 3002 3782
rect 3814 3778 3818 3782
rect 4350 3778 4354 3782
rect 358 3768 362 3772
rect 1286 3768 1290 3772
rect 1758 3768 1762 3772
rect 2758 3768 2762 3772
rect 3286 3768 3290 3772
rect 3366 3768 3370 3772
rect 3886 3768 3890 3772
rect 102 3758 106 3762
rect 958 3758 962 3762
rect 1030 3758 1034 3762
rect 1262 3758 1266 3762
rect 2030 3758 2034 3762
rect 2198 3758 2202 3762
rect 2230 3758 2234 3762
rect 2534 3758 2538 3762
rect 2702 3758 2706 3762
rect 2902 3758 2906 3762
rect 3030 3758 3034 3762
rect 3374 3758 3378 3762
rect 3590 3758 3594 3762
rect 3638 3758 3642 3762
rect 3870 3758 3874 3762
rect 382 3748 386 3752
rect 686 3748 690 3752
rect 886 3748 890 3752
rect 1134 3748 1138 3752
rect 1806 3748 1810 3752
rect 1854 3748 1858 3752
rect 2270 3748 2274 3752
rect 2494 3748 2498 3752
rect 2638 3748 2642 3752
rect 2838 3748 2842 3752
rect 3406 3748 3410 3752
rect 3582 3748 3586 3752
rect 318 3738 322 3742
rect 670 3738 674 3742
rect 902 3738 906 3742
rect 1150 3738 1154 3742
rect 1318 3738 1322 3742
rect 1366 3738 1370 3742
rect 1390 3738 1394 3742
rect 1670 3738 1674 3742
rect 1678 3738 1682 3742
rect 1710 3738 1714 3742
rect 2382 3738 2386 3742
rect 2430 3738 2434 3742
rect 2566 3738 2570 3742
rect 2622 3738 2626 3742
rect 2646 3738 2650 3742
rect 2662 3738 2666 3742
rect 2846 3738 2850 3742
rect 2902 3738 2906 3742
rect 3318 3738 3322 3742
rect 3702 3748 3706 3752
rect 3726 3748 3730 3752
rect 3734 3748 3738 3752
rect 3902 3748 3906 3752
rect 3990 3748 3994 3752
rect 4318 3748 4322 3752
rect 4510 3748 4514 3752
rect 4598 3748 4602 3752
rect 3662 3738 3666 3742
rect 3670 3738 3674 3742
rect 3862 3738 3866 3742
rect 3934 3738 3938 3742
rect 4046 3738 4050 3742
rect 4574 3738 4578 3742
rect 4606 3738 4610 3742
rect 4686 3738 4690 3742
rect 4758 3738 4762 3742
rect 590 3728 594 3732
rect 646 3728 650 3732
rect 1094 3728 1098 3732
rect 1174 3728 1178 3732
rect 2094 3728 2098 3732
rect 2174 3728 2178 3732
rect 2342 3728 2346 3732
rect 3518 3728 3522 3732
rect 3542 3728 3546 3732
rect 3798 3728 3802 3732
rect 4742 3728 4746 3732
rect 358 3718 362 3722
rect 1446 3718 1450 3722
rect 1542 3718 1546 3722
rect 1694 3718 1698 3722
rect 1734 3718 1738 3722
rect 2126 3718 2130 3722
rect 2462 3718 2466 3722
rect 3438 3718 3442 3722
rect 4662 3718 4666 3722
rect 4670 3718 4674 3722
rect 4822 3718 4826 3722
rect 1398 3708 1402 3712
rect 1934 3708 1938 3712
rect 2606 3708 2610 3712
rect 3030 3708 3034 3712
rect 4094 3708 4098 3712
rect 4190 3708 4194 3712
rect 1050 3703 1054 3707
rect 1058 3703 1061 3707
rect 1061 3703 1062 3707
rect 2074 3703 2078 3707
rect 2082 3703 2085 3707
rect 2085 3703 2086 3707
rect 3098 3703 3102 3707
rect 3106 3703 3109 3707
rect 3109 3703 3110 3707
rect 4114 3703 4118 3707
rect 4122 3703 4125 3707
rect 4125 3703 4126 3707
rect 382 3698 386 3702
rect 574 3698 578 3702
rect 766 3698 770 3702
rect 1038 3698 1042 3702
rect 1102 3698 1106 3702
rect 1398 3698 1402 3702
rect 1718 3698 1722 3702
rect 1910 3698 1914 3702
rect 2622 3698 2626 3702
rect 3254 3698 3258 3702
rect 3390 3698 3394 3702
rect 4262 3698 4266 3702
rect 4278 3698 4282 3702
rect 4366 3698 4370 3702
rect 4414 3698 4418 3702
rect 4702 3698 4706 3702
rect 4782 3698 4786 3702
rect 398 3688 402 3692
rect 462 3688 466 3692
rect 1582 3688 1586 3692
rect 1590 3688 1594 3692
rect 1878 3688 1882 3692
rect 2102 3688 2106 3692
rect 2262 3688 2266 3692
rect 2734 3688 2738 3692
rect 3086 3688 3090 3692
rect 3462 3688 3466 3692
rect 3646 3688 3650 3692
rect 3846 3688 3850 3692
rect 3926 3688 3930 3692
rect 3974 3688 3978 3692
rect 478 3678 482 3682
rect 998 3678 1002 3682
rect 1078 3678 1082 3682
rect 1310 3678 1314 3682
rect 1582 3678 1586 3682
rect 1694 3678 1698 3682
rect 1718 3678 1722 3682
rect 1894 3678 1898 3682
rect 2358 3678 2362 3682
rect 2462 3678 2466 3682
rect 2478 3678 2482 3682
rect 3118 3678 3122 3682
rect 3718 3678 3722 3682
rect 3734 3678 3738 3682
rect 4798 3678 4802 3682
rect 5086 3678 5090 3682
rect 478 3668 482 3672
rect 1158 3668 1162 3672
rect 1222 3668 1226 3672
rect 1470 3668 1474 3672
rect 1534 3668 1538 3672
rect 1598 3668 1602 3672
rect 1614 3668 1618 3672
rect 2046 3668 2050 3672
rect 2286 3668 2290 3672
rect 2390 3668 2394 3672
rect 2526 3668 2530 3672
rect 2750 3668 2754 3672
rect 2942 3668 2946 3672
rect 2966 3668 2970 3672
rect 3246 3668 3250 3672
rect 3390 3668 3394 3672
rect 3422 3668 3426 3672
rect 4014 3668 4018 3672
rect 4502 3668 4506 3672
rect 4846 3668 4850 3672
rect 5110 3668 5114 3672
rect 166 3658 170 3662
rect 462 3658 466 3662
rect 502 3658 506 3662
rect 942 3658 946 3662
rect 1078 3658 1082 3662
rect 1110 3658 1114 3662
rect 1142 3658 1146 3662
rect 1166 3658 1170 3662
rect 1646 3658 1650 3662
rect 1750 3658 1754 3662
rect 1790 3658 1794 3662
rect 1814 3658 1818 3662
rect 1902 3658 1906 3662
rect 1982 3658 1986 3662
rect 2422 3658 2426 3662
rect 3254 3658 3258 3662
rect 3326 3658 3330 3662
rect 3446 3658 3450 3662
rect 3454 3658 3458 3662
rect 3518 3658 3522 3662
rect 3542 3658 3546 3662
rect 3878 3658 3882 3662
rect 3998 3658 4002 3662
rect 4270 3658 4274 3662
rect 4358 3658 4362 3662
rect 4454 3658 4458 3662
rect 4702 3658 4706 3662
rect 4854 3658 4858 3662
rect 446 3648 450 3652
rect 694 3648 698 3652
rect 718 3648 722 3652
rect 1486 3648 1490 3652
rect 1582 3648 1586 3652
rect 1590 3648 1594 3652
rect 2182 3648 2186 3652
rect 2238 3648 2242 3652
rect 2406 3648 2410 3652
rect 2614 3648 2618 3652
rect 2662 3648 2666 3652
rect 3446 3648 3450 3652
rect 3686 3648 3690 3652
rect 3702 3648 3706 3652
rect 3870 3648 3874 3652
rect 4462 3648 4466 3652
rect 4622 3648 4626 3652
rect 4798 3648 4802 3652
rect 302 3638 306 3642
rect 470 3638 474 3642
rect 614 3638 618 3642
rect 766 3638 770 3642
rect 878 3638 882 3642
rect 1278 3638 1282 3642
rect 1958 3638 1962 3642
rect 2686 3638 2690 3642
rect 2726 3638 2730 3642
rect 3590 3638 3594 3642
rect 3766 3638 3770 3642
rect 3942 3638 3946 3642
rect 4206 3638 4210 3642
rect 4254 3638 4258 3642
rect 4710 3638 4714 3642
rect 390 3628 394 3632
rect 406 3628 410 3632
rect 1702 3628 1706 3632
rect 2374 3628 2378 3632
rect 4102 3628 4106 3632
rect 4182 3628 4186 3632
rect 4406 3628 4410 3632
rect 4654 3628 4658 3632
rect 4662 3628 4666 3632
rect 734 3618 738 3622
rect 1230 3618 1234 3622
rect 1590 3618 1594 3622
rect 2326 3618 2330 3622
rect 3406 3618 3410 3622
rect 3430 3618 3434 3622
rect 4318 3618 4322 3622
rect 4478 3618 4482 3622
rect 1030 3608 1034 3612
rect 1310 3608 1314 3612
rect 1998 3608 2002 3612
rect 2646 3608 2650 3612
rect 3030 3608 3034 3612
rect 538 3603 542 3607
rect 546 3603 549 3607
rect 549 3603 550 3607
rect 1562 3603 1566 3607
rect 1570 3603 1573 3607
rect 1573 3603 1574 3607
rect 2586 3603 2590 3607
rect 2594 3603 2597 3607
rect 2597 3603 2598 3607
rect 3610 3603 3614 3607
rect 3618 3603 3621 3607
rect 3621 3603 3622 3607
rect 4634 3603 4638 3607
rect 4642 3603 4645 3607
rect 4645 3603 4646 3607
rect 1486 3598 1490 3602
rect 1582 3598 1586 3602
rect 1750 3598 1754 3602
rect 1918 3598 1922 3602
rect 2710 3598 2714 3602
rect 2974 3598 2978 3602
rect 3814 3598 3818 3602
rect 3838 3598 3842 3602
rect 4686 3598 4690 3602
rect 1758 3588 1762 3592
rect 1838 3588 1842 3592
rect 1982 3588 1986 3592
rect 2230 3588 2234 3592
rect 2294 3588 2298 3592
rect 3022 3588 3026 3592
rect 3126 3588 3130 3592
rect 3510 3588 3514 3592
rect 3830 3588 3834 3592
rect 3958 3588 3962 3592
rect 4046 3588 4050 3592
rect 4214 3588 4218 3592
rect 4294 3588 4298 3592
rect 4310 3588 4314 3592
rect 1142 3578 1146 3582
rect 1302 3578 1306 3582
rect 2606 3578 2610 3582
rect 3038 3578 3042 3582
rect 3574 3578 3578 3582
rect 3718 3578 3722 3582
rect 4902 3578 4906 3582
rect 894 3568 898 3572
rect 1382 3568 1386 3572
rect 1422 3568 1426 3572
rect 1926 3568 1930 3572
rect 3502 3568 3506 3572
rect 4430 3568 4434 3572
rect 4750 3568 4754 3572
rect 422 3558 426 3562
rect 726 3558 730 3562
rect 926 3558 930 3562
rect 1166 3558 1170 3562
rect 1246 3558 1250 3562
rect 1318 3558 1322 3562
rect 1678 3558 1682 3562
rect 2958 3558 2962 3562
rect 3126 3558 3130 3562
rect 3342 3558 3346 3562
rect 3742 3558 3746 3562
rect 3918 3558 3922 3562
rect 4510 3558 4514 3562
rect 5054 3558 5058 3562
rect 6 3548 10 3552
rect 358 3548 362 3552
rect 398 3548 402 3552
rect 606 3548 610 3552
rect 678 3548 682 3552
rect 830 3548 834 3552
rect 1390 3548 1394 3552
rect 1622 3548 1626 3552
rect 2038 3548 2042 3552
rect 2054 3548 2058 3552
rect 2414 3548 2418 3552
rect 2438 3548 2442 3552
rect 270 3538 274 3542
rect 414 3538 418 3542
rect 606 3538 610 3542
rect 3078 3548 3082 3552
rect 3302 3548 3306 3552
rect 3910 3548 3914 3552
rect 4134 3548 4138 3552
rect 4406 3548 4410 3552
rect 4510 3548 4514 3552
rect 2358 3538 2362 3542
rect 2478 3538 2482 3542
rect 3454 3538 3458 3542
rect 3478 3538 3482 3542
rect 3782 3538 3786 3542
rect 4310 3538 4314 3542
rect 4502 3538 4506 3542
rect 4758 3538 4762 3542
rect 4886 3538 4890 3542
rect 5150 3538 5154 3542
rect 478 3528 482 3532
rect 598 3528 602 3532
rect 1118 3528 1122 3532
rect 1494 3528 1498 3532
rect 1590 3528 1594 3532
rect 1862 3528 1866 3532
rect 1902 3528 1906 3532
rect 2862 3528 2866 3532
rect 3134 3528 3138 3532
rect 3406 3528 3410 3532
rect 3438 3528 3442 3532
rect 3694 3528 3698 3532
rect 3750 3528 3754 3532
rect 3974 3528 3978 3532
rect 4118 3528 4122 3532
rect 4214 3528 4218 3532
rect 4534 3528 4538 3532
rect 510 3518 514 3522
rect 598 3518 602 3522
rect 1022 3518 1026 3522
rect 1038 3518 1042 3522
rect 1270 3518 1274 3522
rect 1310 3518 1314 3522
rect 1438 3518 1442 3522
rect 1774 3518 1778 3522
rect 2310 3518 2314 3522
rect 3310 3518 3314 3522
rect 3382 3518 3386 3522
rect 6 3508 10 3512
rect 1270 3508 1274 3512
rect 1334 3508 1338 3512
rect 1686 3508 1690 3512
rect 2094 3508 2098 3512
rect 2550 3508 2554 3512
rect 2670 3508 2674 3512
rect 2974 3508 2978 3512
rect 2982 3508 2986 3512
rect 3806 3508 3810 3512
rect 4518 3508 4522 3512
rect 142 3498 146 3502
rect 382 3498 386 3502
rect 1050 3503 1054 3507
rect 1058 3503 1061 3507
rect 1061 3503 1062 3507
rect 2074 3503 2078 3507
rect 2082 3503 2085 3507
rect 2085 3503 2086 3507
rect 3098 3503 3102 3507
rect 3106 3503 3109 3507
rect 3109 3503 3110 3507
rect 4114 3503 4118 3507
rect 4122 3503 4125 3507
rect 4125 3503 4126 3507
rect 1038 3498 1042 3502
rect 1414 3498 1418 3502
rect 1446 3498 1450 3502
rect 1814 3498 1818 3502
rect 2390 3498 2394 3502
rect 3294 3498 3298 3502
rect 3766 3498 3770 3502
rect 4574 3498 4578 3502
rect 1310 3488 1314 3492
rect 2614 3488 2618 3492
rect 174 3478 178 3482
rect 230 3478 234 3482
rect 774 3478 778 3482
rect 1238 3478 1242 3482
rect 1382 3478 1386 3482
rect 1598 3478 1602 3482
rect 2654 3478 2658 3482
rect 2942 3478 2946 3482
rect 3110 3478 3114 3482
rect 3766 3478 3770 3482
rect 3822 3478 3826 3482
rect 3894 3478 3898 3482
rect 4358 3478 4362 3482
rect 4622 3478 4626 3482
rect 5190 3478 5194 3482
rect 158 3468 162 3472
rect 222 3468 226 3472
rect 446 3468 450 3472
rect 494 3468 498 3472
rect 1334 3468 1338 3472
rect 1366 3468 1370 3472
rect 1406 3468 1410 3472
rect 1430 3468 1434 3472
rect 2006 3468 2010 3472
rect 2118 3468 2122 3472
rect 2614 3468 2618 3472
rect 2678 3468 2682 3472
rect 2750 3468 2754 3472
rect 3422 3468 3426 3472
rect 3534 3468 3538 3472
rect 3662 3468 3666 3472
rect 3886 3468 3890 3472
rect 4206 3468 4210 3472
rect 4398 3468 4402 3472
rect 4454 3468 4458 3472
rect 4606 3468 4610 3472
rect 4718 3468 4722 3472
rect 870 3458 874 3462
rect 982 3458 986 3462
rect 990 3458 994 3462
rect 1038 3458 1042 3462
rect 1302 3458 1306 3462
rect 1454 3458 1458 3462
rect 1630 3458 1634 3462
rect 1694 3458 1698 3462
rect 1838 3458 1842 3462
rect 1990 3458 1994 3462
rect 2014 3458 2018 3462
rect 2534 3458 2538 3462
rect 2878 3458 2882 3462
rect 3150 3458 3154 3462
rect 3182 3458 3186 3462
rect 3478 3458 3482 3462
rect 3494 3458 3498 3462
rect 4014 3458 4018 3462
rect 4198 3458 4202 3462
rect 4334 3458 4338 3462
rect 4382 3458 4386 3462
rect 4726 3458 4730 3462
rect 230 3448 234 3452
rect 262 3448 266 3452
rect 398 3448 402 3452
rect 686 3448 690 3452
rect 750 3448 754 3452
rect 806 3448 810 3452
rect 870 3448 874 3452
rect 902 3448 906 3452
rect 958 3448 962 3452
rect 1326 3448 1330 3452
rect 1390 3448 1394 3452
rect 1446 3448 1450 3452
rect 1502 3448 1506 3452
rect 1678 3448 1682 3452
rect 1734 3448 1738 3452
rect 2086 3448 2090 3452
rect 2238 3448 2242 3452
rect 2374 3448 2378 3452
rect 2502 3448 2506 3452
rect 2998 3448 3002 3452
rect 3390 3448 3394 3452
rect 3662 3448 3666 3452
rect 4566 3448 4570 3452
rect 614 3438 618 3442
rect 678 3438 682 3442
rect 1350 3438 1354 3442
rect 1486 3438 1490 3442
rect 1702 3438 1706 3442
rect 2158 3438 2162 3442
rect 2334 3438 2338 3442
rect 2622 3438 2626 3442
rect 2782 3438 2786 3442
rect 3078 3438 3082 3442
rect 3358 3438 3362 3442
rect 3446 3438 3450 3442
rect 3654 3438 3658 3442
rect 3782 3438 3786 3442
rect 3918 3438 3922 3442
rect 4166 3438 4170 3442
rect 4366 3438 4370 3442
rect 4558 3438 4562 3442
rect 4934 3438 4938 3442
rect 1358 3428 1362 3432
rect 1862 3428 1866 3432
rect 2030 3428 2034 3432
rect 2118 3428 2122 3432
rect 2654 3428 2658 3432
rect 3038 3428 3042 3432
rect 3558 3428 3562 3432
rect 4054 3428 4058 3432
rect 4174 3428 4178 3432
rect 5166 3428 5170 3432
rect 238 3418 242 3422
rect 1158 3418 1162 3422
rect 1518 3418 1522 3422
rect 2470 3418 2474 3422
rect 3006 3418 3010 3422
rect 3350 3418 3354 3422
rect 3582 3418 3586 3422
rect 1110 3408 1114 3412
rect 1198 3408 1202 3412
rect 1782 3408 1786 3412
rect 3662 3408 3666 3412
rect 3918 3408 3922 3412
rect 4174 3408 4178 3412
rect 4222 3408 4226 3412
rect 538 3403 542 3407
rect 546 3403 549 3407
rect 549 3403 550 3407
rect 1562 3403 1566 3407
rect 1570 3403 1573 3407
rect 1573 3403 1574 3407
rect 2586 3403 2590 3407
rect 2594 3403 2597 3407
rect 2597 3403 2598 3407
rect 3610 3403 3614 3407
rect 3618 3403 3621 3407
rect 3621 3403 3622 3407
rect 4634 3403 4638 3407
rect 4642 3403 4645 3407
rect 4645 3403 4646 3407
rect 902 3398 906 3402
rect 974 3398 978 3402
rect 1390 3398 1394 3402
rect 2494 3398 2498 3402
rect 2574 3398 2578 3402
rect 846 3388 850 3392
rect 2774 3388 2778 3392
rect 2822 3388 2826 3392
rect 3518 3388 3522 3392
rect 4334 3388 4338 3392
rect 830 3378 834 3382
rect 1142 3378 1146 3382
rect 1470 3378 1474 3382
rect 1678 3378 1682 3382
rect 2110 3378 2114 3382
rect 2966 3378 2970 3382
rect 3638 3378 3642 3382
rect 3974 3378 3978 3382
rect 4726 3378 4730 3382
rect 4998 3378 5002 3382
rect 494 3368 498 3372
rect 550 3368 554 3372
rect 862 3368 866 3372
rect 1254 3368 1258 3372
rect 1582 3368 1586 3372
rect 2782 3368 2786 3372
rect 3206 3368 3210 3372
rect 3966 3368 3970 3372
rect 4654 3368 4658 3372
rect 5174 3368 5178 3372
rect 558 3358 562 3362
rect 1398 3358 1402 3362
rect 1406 3358 1410 3362
rect 1494 3358 1498 3362
rect 1854 3358 1858 3362
rect 2022 3358 2026 3362
rect 2054 3358 2058 3362
rect 2454 3358 2458 3362
rect 3086 3358 3090 3362
rect 3518 3358 3522 3362
rect 3710 3358 3714 3362
rect 4038 3358 4042 3362
rect 4166 3358 4170 3362
rect 4614 3358 4618 3362
rect 4654 3358 4658 3362
rect 4766 3358 4770 3362
rect 4790 3358 4794 3362
rect 4966 3358 4970 3362
rect 4982 3358 4986 3362
rect 5126 3358 5130 3362
rect 5166 3358 5170 3362
rect 94 3348 98 3352
rect 422 3348 426 3352
rect 1422 3348 1426 3352
rect 1734 3348 1738 3352
rect 2278 3348 2282 3352
rect 2670 3348 2674 3352
rect 2686 3348 2690 3352
rect 2734 3348 2738 3352
rect 2974 3348 2978 3352
rect 3134 3348 3138 3352
rect 3622 3348 3626 3352
rect 3726 3348 3730 3352
rect 3734 3348 3738 3352
rect 3974 3348 3978 3352
rect 4142 3348 4146 3352
rect 4294 3348 4298 3352
rect 4390 3348 4394 3352
rect 4558 3348 4562 3352
rect 4574 3348 4578 3352
rect 4590 3348 4594 3352
rect 4870 3348 4874 3352
rect 4918 3348 4922 3352
rect 5006 3348 5010 3352
rect 5062 3348 5066 3352
rect 5134 3348 5138 3352
rect 518 3338 522 3342
rect 742 3338 746 3342
rect 1182 3338 1186 3342
rect 1462 3338 1466 3342
rect 1502 3338 1506 3342
rect 1710 3338 1714 3342
rect 2038 3338 2042 3342
rect 2334 3338 2338 3342
rect 2454 3338 2458 3342
rect 2630 3338 2634 3342
rect 2822 3338 2826 3342
rect 2902 3338 2906 3342
rect 3254 3338 3258 3342
rect 3494 3338 3498 3342
rect 3838 3338 3842 3342
rect 3974 3338 3978 3342
rect 4078 3338 4082 3342
rect 4094 3338 4098 3342
rect 4246 3338 4250 3342
rect 4790 3338 4794 3342
rect 5078 3338 5082 3342
rect 5086 3338 5090 3342
rect 238 3328 242 3332
rect 342 3328 346 3332
rect 422 3328 426 3332
rect 670 3328 674 3332
rect 966 3328 970 3332
rect 1214 3328 1218 3332
rect 1270 3328 1274 3332
rect 1422 3328 1426 3332
rect 2014 3328 2018 3332
rect 2550 3328 2554 3332
rect 2558 3328 2562 3332
rect 3030 3328 3034 3332
rect 3062 3328 3066 3332
rect 3078 3328 3082 3332
rect 3350 3328 3354 3332
rect 3742 3328 3746 3332
rect 4190 3328 4194 3332
rect 4526 3328 4530 3332
rect 4574 3328 4578 3332
rect 4750 3328 4754 3332
rect 5078 3328 5082 3332
rect 5158 3328 5162 3332
rect 158 3318 162 3322
rect 382 3318 386 3322
rect 478 3318 482 3322
rect 910 3318 914 3322
rect 1070 3318 1074 3322
rect 1470 3318 1474 3322
rect 2886 3318 2890 3322
rect 3150 3318 3154 3322
rect 3910 3318 3914 3322
rect 4150 3318 4154 3322
rect 4158 3318 4162 3322
rect 4614 3318 4618 3322
rect 1430 3308 1434 3312
rect 1806 3308 1810 3312
rect 3078 3308 3082 3312
rect 3398 3308 3402 3312
rect 3550 3308 3554 3312
rect 4590 3308 4594 3312
rect 4702 3308 4706 3312
rect 4918 3308 4922 3312
rect 1050 3303 1054 3307
rect 1058 3303 1061 3307
rect 1061 3303 1062 3307
rect 2074 3303 2078 3307
rect 2082 3303 2085 3307
rect 2085 3303 2086 3307
rect 3098 3303 3102 3307
rect 3106 3303 3109 3307
rect 3109 3303 3110 3307
rect 4114 3303 4118 3307
rect 4122 3303 4125 3307
rect 4125 3303 4126 3307
rect 2102 3298 2106 3302
rect 2286 3298 2290 3302
rect 2462 3298 2466 3302
rect 2790 3298 2794 3302
rect 2926 3298 2930 3302
rect 3086 3298 3090 3302
rect 3310 3298 3314 3302
rect 3326 3298 3330 3302
rect 3398 3298 3402 3302
rect 3654 3298 3658 3302
rect 4262 3298 4266 3302
rect 4430 3298 4434 3302
rect 4742 3298 4746 3302
rect 4974 3298 4978 3302
rect 1254 3288 1258 3292
rect 1502 3288 1506 3292
rect 2790 3288 2794 3292
rect 3774 3288 3778 3292
rect 4038 3288 4042 3292
rect 4182 3288 4186 3292
rect 4854 3288 4858 3292
rect 606 3278 610 3282
rect 622 3278 626 3282
rect 1534 3278 1538 3282
rect 1870 3278 1874 3282
rect 2190 3278 2194 3282
rect 3262 3278 3266 3282
rect 3558 3278 3562 3282
rect 3726 3278 3730 3282
rect 3966 3278 3970 3282
rect 4190 3278 4194 3282
rect 4766 3278 4770 3282
rect 4830 3278 4834 3282
rect 4862 3278 4866 3282
rect 4934 3278 4938 3282
rect 222 3268 226 3272
rect 446 3268 450 3272
rect 886 3268 890 3272
rect 990 3268 994 3272
rect 1182 3268 1186 3272
rect 1190 3268 1194 3272
rect 1342 3268 1346 3272
rect 1510 3268 1514 3272
rect 2142 3268 2146 3272
rect 2254 3268 2258 3272
rect 2350 3268 2354 3272
rect 2638 3268 2642 3272
rect 2662 3268 2666 3272
rect 2718 3268 2722 3272
rect 3198 3268 3202 3272
rect 3262 3268 3266 3272
rect 3550 3268 3554 3272
rect 3662 3268 3666 3272
rect 3670 3268 3674 3272
rect 3734 3268 3738 3272
rect 3982 3268 3986 3272
rect 4150 3268 4154 3272
rect 4534 3268 4538 3272
rect 126 3258 130 3262
rect 398 3258 402 3262
rect 694 3258 698 3262
rect 1086 3258 1090 3262
rect 1150 3258 1154 3262
rect 1174 3258 1178 3262
rect 1382 3258 1386 3262
rect 1670 3258 1674 3262
rect 1950 3258 1954 3262
rect 2382 3258 2386 3262
rect 2614 3258 2618 3262
rect 2814 3258 2818 3262
rect 2894 3258 2898 3262
rect 2966 3258 2970 3262
rect 3462 3258 3466 3262
rect 3470 3258 3474 3262
rect 3990 3258 3994 3262
rect 4134 3258 4138 3262
rect 4238 3258 4242 3262
rect 4406 3258 4410 3262
rect 4558 3258 4562 3262
rect 4782 3258 4786 3262
rect 6 3248 10 3252
rect 662 3248 666 3252
rect 918 3248 922 3252
rect 1006 3248 1010 3252
rect 1118 3248 1122 3252
rect 1182 3248 1186 3252
rect 1278 3248 1282 3252
rect 1470 3248 1474 3252
rect 1774 3248 1778 3252
rect 1902 3248 1906 3252
rect 2126 3248 2130 3252
rect 2310 3248 2314 3252
rect 2694 3248 2698 3252
rect 2734 3248 2738 3252
rect 2774 3248 2778 3252
rect 2798 3248 2802 3252
rect 2990 3248 2994 3252
rect 3478 3248 3482 3252
rect 3542 3248 3546 3252
rect 3558 3248 3562 3252
rect 4574 3248 4578 3252
rect 5190 3248 5194 3252
rect 1190 3238 1194 3242
rect 1966 3238 1970 3242
rect 2854 3238 2858 3242
rect 3358 3238 3362 3242
rect 4222 3238 4226 3242
rect 4470 3238 4474 3242
rect 4806 3238 4810 3242
rect 4926 3238 4930 3242
rect 550 3228 554 3232
rect 1358 3228 1362 3232
rect 1502 3228 1506 3232
rect 2046 3228 2050 3232
rect 2638 3228 2642 3232
rect 2902 3228 2906 3232
rect 3318 3228 3322 3232
rect 3590 3228 3594 3232
rect 3894 3228 3898 3232
rect 4862 3228 4866 3232
rect 326 3218 330 3222
rect 806 3218 810 3222
rect 1758 3218 1762 3222
rect 1942 3218 1946 3222
rect 2510 3218 2514 3222
rect 3718 3218 3722 3222
rect 4142 3218 4146 3222
rect 4310 3218 4314 3222
rect 4438 3218 4442 3222
rect 4782 3218 4786 3222
rect 430 3208 434 3212
rect 566 3208 570 3212
rect 934 3208 938 3212
rect 1662 3208 1666 3212
rect 1806 3208 1810 3212
rect 2638 3208 2642 3212
rect 2814 3208 2818 3212
rect 3246 3208 3250 3212
rect 3678 3208 3682 3212
rect 3790 3208 3794 3212
rect 4742 3208 4746 3212
rect 538 3203 542 3207
rect 546 3203 549 3207
rect 549 3203 550 3207
rect 1562 3203 1566 3207
rect 1570 3203 1573 3207
rect 1573 3203 1574 3207
rect 2586 3203 2590 3207
rect 2594 3203 2597 3207
rect 2597 3203 2598 3207
rect 3610 3203 3614 3207
rect 3618 3203 3621 3207
rect 3621 3203 3622 3207
rect 4634 3203 4638 3207
rect 4642 3203 4645 3207
rect 4645 3203 4646 3207
rect 1094 3198 1098 3202
rect 1902 3198 1906 3202
rect 2214 3198 2218 3202
rect 2606 3198 2610 3202
rect 3086 3198 3090 3202
rect 3694 3198 3698 3202
rect 1222 3188 1226 3192
rect 1462 3188 1466 3192
rect 1750 3188 1754 3192
rect 1998 3188 2002 3192
rect 2718 3188 2722 3192
rect 3062 3188 3066 3192
rect 3390 3188 3394 3192
rect 4190 3188 4194 3192
rect 4982 3188 4986 3192
rect 1134 3178 1138 3182
rect 1158 3178 1162 3182
rect 1638 3178 1642 3182
rect 2102 3178 2106 3182
rect 2550 3178 2554 3182
rect 2918 3178 2922 3182
rect 3422 3178 3426 3182
rect 4950 3178 4954 3182
rect 814 3168 818 3172
rect 1494 3168 1498 3172
rect 1798 3168 1802 3172
rect 1910 3168 1914 3172
rect 1990 3168 1994 3172
rect 2230 3168 2234 3172
rect 2438 3168 2442 3172
rect 2606 3168 2610 3172
rect 3694 3168 3698 3172
rect 3830 3168 3834 3172
rect 5142 3168 5146 3172
rect 334 3158 338 3162
rect 766 3158 770 3162
rect 830 3158 834 3162
rect 926 3158 930 3162
rect 982 3158 986 3162
rect 1174 3158 1178 3162
rect 1502 3158 1506 3162
rect 1678 3158 1682 3162
rect 1854 3158 1858 3162
rect 1934 3158 1938 3162
rect 1942 3158 1946 3162
rect 2862 3158 2866 3162
rect 3926 3158 3930 3162
rect 4262 3158 4266 3162
rect 4726 3158 4730 3162
rect 4806 3158 4810 3162
rect 4934 3158 4938 3162
rect 14 3148 18 3152
rect 102 3148 106 3152
rect 718 3148 722 3152
rect 950 3148 954 3152
rect 990 3148 994 3152
rect 1118 3148 1122 3152
rect 1198 3148 1202 3152
rect 1334 3148 1338 3152
rect 1550 3148 1554 3152
rect 1950 3148 1954 3152
rect 2166 3148 2170 3152
rect 2942 3148 2946 3152
rect 3374 3148 3378 3152
rect 4206 3148 4210 3152
rect 4510 3148 4514 3152
rect 4726 3148 4730 3152
rect 4990 3148 4994 3152
rect 374 3138 378 3142
rect 382 3138 386 3142
rect 390 3138 394 3142
rect 622 3138 626 3142
rect 686 3138 690 3142
rect 734 3138 738 3142
rect 758 3138 762 3142
rect 814 3138 818 3142
rect 1014 3138 1018 3142
rect 1294 3138 1298 3142
rect 1470 3138 1474 3142
rect 1526 3138 1530 3142
rect 1606 3138 1610 3142
rect 1726 3138 1730 3142
rect 1974 3138 1978 3142
rect 2358 3138 2362 3142
rect 2430 3138 2434 3142
rect 2502 3138 2506 3142
rect 2934 3138 2938 3142
rect 2966 3138 2970 3142
rect 3038 3138 3042 3142
rect 3470 3138 3474 3142
rect 3838 3138 3842 3142
rect 4062 3138 4066 3142
rect 4662 3138 4666 3142
rect 4678 3138 4682 3142
rect 4758 3138 4762 3142
rect 4910 3138 4914 3142
rect 4942 3138 4946 3142
rect 1030 3128 1034 3132
rect 1190 3128 1194 3132
rect 1326 3128 1330 3132
rect 1438 3128 1442 3132
rect 1686 3128 1690 3132
rect 1830 3128 1834 3132
rect 2094 3128 2098 3132
rect 2790 3128 2794 3132
rect 2878 3128 2882 3132
rect 2974 3128 2978 3132
rect 3142 3128 3146 3132
rect 3446 3128 3450 3132
rect 3462 3128 3466 3132
rect 3734 3128 3738 3132
rect 4102 3128 4106 3132
rect 4174 3128 4178 3132
rect 4758 3128 4762 3132
rect 894 3118 898 3122
rect 974 3118 978 3122
rect 998 3118 1002 3122
rect 1414 3118 1418 3122
rect 1710 3118 1714 3122
rect 2542 3118 2546 3122
rect 2870 3118 2874 3122
rect 3358 3118 3362 3122
rect 3806 3118 3810 3122
rect 3878 3118 3882 3122
rect 4158 3118 4162 3122
rect 4518 3118 4522 3122
rect 118 3108 122 3112
rect 1206 3108 1210 3112
rect 1278 3108 1282 3112
rect 1318 3108 1322 3112
rect 1654 3108 1658 3112
rect 1790 3108 1794 3112
rect 1798 3108 1802 3112
rect 2062 3108 2066 3112
rect 2270 3108 2274 3112
rect 2526 3108 2530 3112
rect 3030 3108 3034 3112
rect 4262 3108 4266 3112
rect 5086 3108 5090 3112
rect 430 3098 434 3102
rect 1050 3103 1054 3107
rect 1058 3103 1061 3107
rect 1061 3103 1062 3107
rect 2074 3103 2078 3107
rect 2082 3103 2085 3107
rect 2085 3103 2086 3107
rect 3098 3103 3102 3107
rect 3106 3103 3109 3107
rect 3109 3103 3110 3107
rect 4114 3103 4118 3107
rect 4122 3103 4125 3107
rect 4125 3103 4126 3107
rect 814 3098 818 3102
rect 894 3098 898 3102
rect 1598 3098 1602 3102
rect 2054 3098 2058 3102
rect 2742 3098 2746 3102
rect 2830 3098 2834 3102
rect 3182 3098 3186 3102
rect 3686 3098 3690 3102
rect 3942 3098 3946 3102
rect 4470 3098 4474 3102
rect 4774 3098 4778 3102
rect 710 3088 714 3092
rect 1110 3088 1114 3092
rect 326 3078 330 3082
rect 1678 3088 1682 3092
rect 1846 3088 1850 3092
rect 2262 3088 2266 3092
rect 2774 3088 2778 3092
rect 3078 3088 3082 3092
rect 3310 3088 3314 3092
rect 3822 3088 3826 3092
rect 4238 3088 4242 3092
rect 4894 3088 4898 3092
rect 4974 3088 4978 3092
rect 1486 3078 1490 3082
rect 1606 3078 1610 3082
rect 1702 3078 1706 3082
rect 1782 3078 1786 3082
rect 1966 3078 1970 3082
rect 342 3068 346 3072
rect 518 3068 522 3072
rect 774 3068 778 3072
rect 822 3068 826 3072
rect 942 3068 946 3072
rect 1358 3068 1362 3072
rect 1374 3068 1378 3072
rect 1454 3068 1458 3072
rect 1614 3068 1618 3072
rect 1622 3068 1626 3072
rect 1950 3068 1954 3072
rect 2518 3078 2522 3082
rect 2822 3078 2826 3082
rect 2902 3078 2906 3082
rect 3038 3078 3042 3082
rect 3686 3078 3690 3082
rect 3726 3078 3730 3082
rect 3830 3078 3834 3082
rect 3918 3078 3922 3082
rect 4038 3078 4042 3082
rect 4774 3078 4778 3082
rect 5086 3078 5090 3082
rect 2318 3068 2322 3072
rect 2334 3068 2338 3072
rect 2526 3068 2530 3072
rect 2550 3068 2554 3072
rect 2574 3068 2578 3072
rect 2862 3068 2866 3072
rect 2902 3068 2906 3072
rect 3326 3068 3330 3072
rect 3342 3068 3346 3072
rect 3918 3068 3922 3072
rect 3942 3068 3946 3072
rect 4198 3068 4202 3072
rect 4342 3068 4346 3072
rect 4350 3068 4354 3072
rect 182 3058 186 3062
rect 398 3058 402 3062
rect 574 3058 578 3062
rect 622 3058 626 3062
rect 1158 3058 1162 3062
rect 1206 3058 1210 3062
rect 1294 3058 1298 3062
rect 1470 3058 1474 3062
rect 1910 3058 1914 3062
rect 1982 3058 1986 3062
rect 2182 3058 2186 3062
rect 2422 3058 2426 3062
rect 2486 3058 2490 3062
rect 2502 3058 2506 3062
rect 3526 3058 3530 3062
rect 3958 3058 3962 3062
rect 3998 3058 4002 3062
rect 4014 3058 4018 3062
rect 4262 3058 4266 3062
rect 4486 3058 4490 3062
rect 4670 3058 4674 3062
rect 5134 3058 5138 3062
rect 686 3048 690 3052
rect 1206 3048 1210 3052
rect 1350 3048 1354 3052
rect 1358 3048 1362 3052
rect 1478 3048 1482 3052
rect 1582 3048 1586 3052
rect 1702 3048 1706 3052
rect 1782 3048 1786 3052
rect 2286 3048 2290 3052
rect 2510 3048 2514 3052
rect 2726 3048 2730 3052
rect 3246 3048 3250 3052
rect 3470 3048 3474 3052
rect 3518 3048 3522 3052
rect 3526 3048 3530 3052
rect 4134 3048 4138 3052
rect 4142 3048 4146 3052
rect 870 3038 874 3042
rect 934 3038 938 3042
rect 950 3038 954 3042
rect 4286 3048 4290 3052
rect 4614 3048 4618 3052
rect 5150 3048 5154 3052
rect 1758 3038 1762 3042
rect 2438 3038 2442 3042
rect 2718 3038 2722 3042
rect 3342 3038 3346 3042
rect 3518 3038 3522 3042
rect 4006 3038 4010 3042
rect 4070 3038 4074 3042
rect 4342 3038 4346 3042
rect 5070 3038 5074 3042
rect 5086 3038 5090 3042
rect 246 3028 250 3032
rect 958 3028 962 3032
rect 1142 3028 1146 3032
rect 1358 3028 1362 3032
rect 1398 3028 1402 3032
rect 1662 3028 1666 3032
rect 2270 3028 2274 3032
rect 2278 3028 2282 3032
rect 2438 3028 2442 3032
rect 2838 3028 2842 3032
rect 3510 3028 3514 3032
rect 4278 3028 4282 3032
rect 1486 3018 1490 3022
rect 2342 3018 2346 3022
rect 2910 3018 2914 3022
rect 4022 3018 4026 3022
rect 4094 3018 4098 3022
rect 4166 3018 4170 3022
rect 4478 3018 4482 3022
rect 1238 3008 1242 3012
rect 1582 3008 1586 3012
rect 1814 3008 1818 3012
rect 1974 3008 1978 3012
rect 2398 3008 2402 3012
rect 2534 3008 2538 3012
rect 3838 3008 3842 3012
rect 3966 3008 3970 3012
rect 4382 3008 4386 3012
rect 4462 3008 4466 3012
rect 4622 3008 4626 3012
rect 538 3003 542 3007
rect 546 3003 549 3007
rect 549 3003 550 3007
rect 1562 3003 1566 3007
rect 1570 3003 1573 3007
rect 1573 3003 1574 3007
rect 2586 3003 2590 3007
rect 2594 3003 2597 3007
rect 2597 3003 2598 3007
rect 3610 3003 3614 3007
rect 3618 3003 3621 3007
rect 3621 3003 3622 3007
rect 4634 3003 4638 3007
rect 4642 3003 4645 3007
rect 4645 3003 4646 3007
rect 1502 2998 1506 3002
rect 3406 2998 3410 3002
rect 3758 2998 3762 3002
rect 4006 2998 4010 3002
rect 4870 2998 4874 3002
rect 366 2988 370 2992
rect 918 2988 922 2992
rect 1422 2988 1426 2992
rect 1534 2988 1538 2992
rect 1758 2988 1762 2992
rect 1870 2988 1874 2992
rect 1982 2988 1986 2992
rect 2222 2988 2226 2992
rect 2838 2988 2842 2992
rect 2950 2988 2954 2992
rect 3710 2988 3714 2992
rect 3998 2988 4002 2992
rect 4206 2988 4210 2992
rect 4462 2988 4466 2992
rect 974 2978 978 2982
rect 1134 2978 1138 2982
rect 1398 2978 1402 2982
rect 1534 2978 1538 2982
rect 2166 2978 2170 2982
rect 3190 2978 3194 2982
rect 3494 2978 3498 2982
rect 3854 2978 3858 2982
rect 1014 2968 1018 2972
rect 1318 2968 1322 2972
rect 1390 2968 1394 2972
rect 2534 2968 2538 2972
rect 2678 2968 2682 2972
rect 2702 2968 2706 2972
rect 2774 2968 2778 2972
rect 3022 2968 3026 2972
rect 3286 2968 3290 2972
rect 3550 2968 3554 2972
rect 3886 2968 3890 2972
rect 4782 2968 4786 2972
rect 4950 2968 4954 2972
rect 4982 2968 4986 2972
rect 5158 2968 5162 2972
rect 646 2958 650 2962
rect 1174 2958 1178 2962
rect 1806 2958 1810 2962
rect 2486 2958 2490 2962
rect 2734 2958 2738 2962
rect 2758 2958 2762 2962
rect 3606 2958 3610 2962
rect 3718 2958 3722 2962
rect 3774 2958 3778 2962
rect 3982 2958 3986 2962
rect 4182 2958 4186 2962
rect 4590 2958 4594 2962
rect 4694 2958 4698 2962
rect 206 2948 210 2952
rect 566 2948 570 2952
rect 654 2948 658 2952
rect 678 2948 682 2952
rect 734 2948 738 2952
rect 774 2948 778 2952
rect 870 2948 874 2952
rect 1046 2948 1050 2952
rect 1142 2948 1146 2952
rect 1342 2948 1346 2952
rect 1630 2948 1634 2952
rect 1694 2948 1698 2952
rect 2014 2948 2018 2952
rect 2494 2948 2498 2952
rect 2534 2948 2538 2952
rect 2606 2948 2610 2952
rect 2630 2948 2634 2952
rect 2646 2948 2650 2952
rect 2950 2948 2954 2952
rect 3126 2948 3130 2952
rect 3358 2948 3362 2952
rect 358 2938 362 2942
rect 526 2938 530 2942
rect 750 2938 754 2942
rect 790 2938 794 2942
rect 1118 2938 1122 2942
rect 1302 2938 1306 2942
rect 1318 2938 1322 2942
rect 1438 2938 1442 2942
rect 1702 2938 1706 2942
rect 1750 2938 1754 2942
rect 2014 2938 2018 2942
rect 2166 2938 2170 2942
rect 2286 2938 2290 2942
rect 2310 2938 2314 2942
rect 2326 2938 2330 2942
rect 3662 2948 3666 2952
rect 3718 2948 3722 2952
rect 3966 2948 3970 2952
rect 4310 2948 4314 2952
rect 4630 2948 4634 2952
rect 4838 2948 4842 2952
rect 4998 2948 5002 2952
rect 5174 2948 5178 2952
rect 2622 2938 2626 2942
rect 2982 2938 2986 2942
rect 3110 2938 3114 2942
rect 3278 2938 3282 2942
rect 3318 2938 3322 2942
rect 4030 2938 4034 2942
rect 4038 2938 4042 2942
rect 4134 2938 4138 2942
rect 4182 2938 4186 2942
rect 4206 2938 4210 2942
rect 4398 2938 4402 2942
rect 4454 2938 4458 2942
rect 5118 2938 5122 2942
rect 454 2928 458 2932
rect 654 2928 658 2932
rect 982 2928 986 2932
rect 1190 2928 1194 2932
rect 1814 2928 1818 2932
rect 2150 2928 2154 2932
rect 2486 2928 2490 2932
rect 2606 2928 2610 2932
rect 3198 2928 3202 2932
rect 3238 2928 3242 2932
rect 3574 2928 3578 2932
rect 3798 2928 3802 2932
rect 3870 2928 3874 2932
rect 4030 2928 4034 2932
rect 4078 2928 4082 2932
rect 4126 2928 4130 2932
rect 4342 2928 4346 2932
rect 4398 2928 4402 2932
rect 5102 2928 5106 2932
rect 630 2918 634 2922
rect 774 2918 778 2922
rect 1014 2918 1018 2922
rect 1222 2918 1226 2922
rect 1462 2918 1466 2922
rect 1910 2918 1914 2922
rect 2046 2918 2050 2922
rect 2758 2918 2762 2922
rect 2814 2918 2818 2922
rect 3022 2918 3026 2922
rect 3150 2918 3154 2922
rect 3318 2918 3322 2922
rect 3326 2918 3330 2922
rect 3766 2918 3770 2922
rect 3830 2918 3834 2922
rect 4262 2918 4266 2922
rect 4462 2918 4466 2922
rect 4582 2918 4586 2922
rect 238 2908 242 2912
rect 958 2908 962 2912
rect 1078 2908 1082 2912
rect 1446 2908 1450 2912
rect 1542 2908 1546 2912
rect 2022 2908 2026 2912
rect 2622 2908 2626 2912
rect 2630 2908 2634 2912
rect 2782 2908 2786 2912
rect 3070 2908 3074 2912
rect 4054 2908 4058 2912
rect 4334 2908 4338 2912
rect 4814 2908 4818 2912
rect 1050 2903 1054 2907
rect 1058 2903 1061 2907
rect 1061 2903 1062 2907
rect 2074 2903 2078 2907
rect 2082 2903 2085 2907
rect 2085 2903 2086 2907
rect 3098 2903 3102 2907
rect 3106 2903 3109 2907
rect 3109 2903 3110 2907
rect 4114 2903 4118 2907
rect 4122 2903 4125 2907
rect 4125 2903 4126 2907
rect 246 2898 250 2902
rect 662 2898 666 2902
rect 1374 2898 1378 2902
rect 1782 2898 1786 2902
rect 2462 2898 2466 2902
rect 2662 2898 2666 2902
rect 2774 2898 2778 2902
rect 2886 2898 2890 2902
rect 3118 2898 3122 2902
rect 3750 2898 3754 2902
rect 3846 2898 3850 2902
rect 4846 2898 4850 2902
rect 4902 2898 4906 2902
rect 5030 2898 5034 2902
rect 822 2888 826 2892
rect 838 2888 842 2892
rect 950 2888 954 2892
rect 1030 2888 1034 2892
rect 1078 2888 1082 2892
rect 1094 2888 1098 2892
rect 1230 2888 1234 2892
rect 1318 2888 1322 2892
rect 1582 2888 1586 2892
rect 1662 2888 1666 2892
rect 1694 2888 1698 2892
rect 1830 2888 1834 2892
rect 2006 2888 2010 2892
rect 2646 2888 2650 2892
rect 2806 2888 2810 2892
rect 3630 2888 3634 2892
rect 3678 2888 3682 2892
rect 4702 2888 4706 2892
rect 5062 2888 5066 2892
rect 902 2878 906 2882
rect 934 2878 938 2882
rect 1582 2878 1586 2882
rect 1630 2878 1634 2882
rect 1662 2878 1666 2882
rect 3278 2878 3282 2882
rect 3678 2878 3682 2882
rect 4190 2878 4194 2882
rect 4454 2878 4458 2882
rect 4622 2878 4626 2882
rect 102 2868 106 2872
rect 766 2868 770 2872
rect 894 2868 898 2872
rect 1086 2868 1090 2872
rect 1214 2868 1218 2872
rect 1326 2868 1330 2872
rect 1494 2868 1498 2872
rect 1510 2868 1514 2872
rect 1542 2868 1546 2872
rect 1630 2868 1634 2872
rect 1678 2868 1682 2872
rect 1862 2868 1866 2872
rect 1902 2868 1906 2872
rect 1942 2868 1946 2872
rect 2038 2868 2042 2872
rect 2222 2868 2226 2872
rect 2470 2868 2474 2872
rect 2550 2868 2554 2872
rect 2646 2868 2650 2872
rect 2670 2868 2674 2872
rect 2838 2868 2842 2872
rect 3350 2868 3354 2872
rect 3870 2868 3874 2872
rect 4526 2868 4530 2872
rect 4598 2868 4602 2872
rect 4750 2868 4754 2872
rect 398 2858 402 2862
rect 574 2858 578 2862
rect 1094 2858 1098 2862
rect 1110 2858 1114 2862
rect 1182 2858 1186 2862
rect 1270 2858 1274 2862
rect 1670 2858 1674 2862
rect 1774 2858 1778 2862
rect 2798 2858 2802 2862
rect 2974 2858 2978 2862
rect 3174 2858 3178 2862
rect 3390 2858 3394 2862
rect 3398 2858 3402 2862
rect 3510 2858 3514 2862
rect 3614 2858 3618 2862
rect 4142 2858 4146 2862
rect 4166 2858 4170 2862
rect 4518 2858 4522 2862
rect 4542 2858 4546 2862
rect 4622 2858 4626 2862
rect 4734 2858 4738 2862
rect 870 2848 874 2852
rect 1590 2848 1594 2852
rect 1606 2848 1610 2852
rect 1750 2848 1754 2852
rect 1758 2848 1762 2852
rect 2014 2848 2018 2852
rect 2054 2848 2058 2852
rect 2142 2848 2146 2852
rect 2166 2848 2170 2852
rect 2310 2848 2314 2852
rect 2470 2848 2474 2852
rect 2478 2848 2482 2852
rect 3022 2848 3026 2852
rect 3118 2848 3122 2852
rect 3254 2848 3258 2852
rect 3550 2848 3554 2852
rect 3678 2848 3682 2852
rect 3758 2848 3762 2852
rect 3846 2848 3850 2852
rect 3910 2848 3914 2852
rect 4454 2848 4458 2852
rect 4526 2848 4530 2852
rect 4710 2848 4714 2852
rect 4790 2848 4794 2852
rect 1110 2838 1114 2842
rect 1270 2838 1274 2842
rect 1342 2838 1346 2842
rect 2382 2838 2386 2842
rect 2830 2838 2834 2842
rect 3334 2838 3338 2842
rect 3342 2838 3346 2842
rect 3414 2838 3418 2842
rect 3566 2838 3570 2842
rect 3806 2838 3810 2842
rect 4622 2838 4626 2842
rect 1334 2828 1338 2832
rect 1358 2828 1362 2832
rect 1550 2828 1554 2832
rect 1678 2828 1682 2832
rect 1878 2828 1882 2832
rect 2118 2828 2122 2832
rect 2678 2828 2682 2832
rect 2750 2828 2754 2832
rect 2878 2828 2882 2832
rect 3166 2828 3170 2832
rect 3302 2828 3306 2832
rect 4334 2828 4338 2832
rect 4422 2828 4426 2832
rect 4974 2828 4978 2832
rect 774 2818 778 2822
rect 2206 2818 2210 2822
rect 3086 2818 3090 2822
rect 3326 2818 3330 2822
rect 3646 2818 3650 2822
rect 4222 2818 4226 2822
rect 4350 2818 4354 2822
rect 5014 2818 5018 2822
rect 1454 2808 1458 2812
rect 1678 2808 1682 2812
rect 2414 2808 2418 2812
rect 2510 2808 2514 2812
rect 2790 2808 2794 2812
rect 3358 2808 3362 2812
rect 3678 2808 3682 2812
rect 4086 2808 4090 2812
rect 4198 2808 4202 2812
rect 538 2803 542 2807
rect 546 2803 549 2807
rect 549 2803 550 2807
rect 1562 2803 1566 2807
rect 1570 2803 1573 2807
rect 1573 2803 1574 2807
rect 2586 2803 2590 2807
rect 2594 2803 2597 2807
rect 2597 2803 2598 2807
rect 838 2798 842 2802
rect 1198 2798 1202 2802
rect 1438 2798 1442 2802
rect 1478 2798 1482 2802
rect 1782 2798 1786 2802
rect 1966 2798 1970 2802
rect 2046 2798 2050 2802
rect 2102 2798 2106 2802
rect 3610 2803 3614 2807
rect 3618 2803 3621 2807
rect 3621 2803 3622 2807
rect 4634 2803 4638 2807
rect 4642 2803 4645 2807
rect 4645 2803 4646 2807
rect 3390 2798 3394 2802
rect 3766 2798 3770 2802
rect 3934 2798 3938 2802
rect 406 2788 410 2792
rect 1118 2788 1122 2792
rect 1702 2788 1706 2792
rect 1806 2788 1810 2792
rect 2406 2788 2410 2792
rect 2814 2788 2818 2792
rect 2838 2788 2842 2792
rect 3246 2788 3250 2792
rect 3310 2788 3314 2792
rect 3502 2788 3506 2792
rect 1782 2778 1786 2782
rect 2134 2778 2138 2782
rect 2518 2778 2522 2782
rect 2854 2778 2858 2782
rect 3102 2778 3106 2782
rect 3278 2778 3282 2782
rect 4566 2778 4570 2782
rect 502 2768 506 2772
rect 742 2768 746 2772
rect 1126 2768 1130 2772
rect 1494 2768 1498 2772
rect 1854 2768 1858 2772
rect 1990 2768 1994 2772
rect 2454 2768 2458 2772
rect 3478 2768 3482 2772
rect 3558 2768 3562 2772
rect 3614 2768 3618 2772
rect 3878 2768 3882 2772
rect 3894 2768 3898 2772
rect 4350 2768 4354 2772
rect 4462 2768 4466 2772
rect 4758 2768 4762 2772
rect 5190 2768 5194 2772
rect 382 2758 386 2762
rect 654 2758 658 2762
rect 1198 2758 1202 2762
rect 1422 2758 1426 2762
rect 1678 2758 1682 2762
rect 2086 2758 2090 2762
rect 2158 2758 2162 2762
rect 2838 2758 2842 2762
rect 3038 2758 3042 2762
rect 3854 2758 3858 2762
rect 4182 2758 4186 2762
rect 4278 2758 4282 2762
rect 4902 2758 4906 2762
rect 5014 2758 5018 2762
rect 5110 2758 5114 2762
rect 6 2738 10 2742
rect 582 2748 586 2752
rect 854 2748 858 2752
rect 950 2748 954 2752
rect 1006 2748 1010 2752
rect 1142 2748 1146 2752
rect 1542 2748 1546 2752
rect 1798 2748 1802 2752
rect 1830 2748 1834 2752
rect 1862 2748 1866 2752
rect 814 2738 818 2742
rect 1942 2748 1946 2752
rect 2102 2748 2106 2752
rect 2198 2748 2202 2752
rect 2358 2748 2362 2752
rect 2550 2748 2554 2752
rect 3390 2748 3394 2752
rect 3502 2748 3506 2752
rect 3550 2748 3554 2752
rect 1406 2738 1410 2742
rect 1622 2738 1626 2742
rect 1718 2738 1722 2742
rect 1750 2738 1754 2742
rect 1774 2738 1778 2742
rect 2142 2738 2146 2742
rect 2158 2738 2162 2742
rect 3806 2748 3810 2752
rect 3830 2748 3834 2752
rect 3894 2748 3898 2752
rect 3942 2748 3946 2752
rect 4062 2748 4066 2752
rect 4086 2748 4090 2752
rect 4678 2748 4682 2752
rect 4758 2748 4762 2752
rect 4830 2748 4834 2752
rect 2870 2738 2874 2742
rect 2942 2738 2946 2742
rect 3782 2738 3786 2742
rect 3798 2738 3802 2742
rect 3902 2738 3906 2742
rect 4398 2738 4402 2742
rect 4742 2738 4746 2742
rect 4958 2738 4962 2742
rect 5014 2738 5018 2742
rect 798 2728 802 2732
rect 822 2728 826 2732
rect 1422 2728 1426 2732
rect 1502 2728 1506 2732
rect 1774 2728 1778 2732
rect 1878 2728 1882 2732
rect 2038 2728 2042 2732
rect 2222 2728 2226 2732
rect 2270 2728 2274 2732
rect 2350 2728 2354 2732
rect 2542 2728 2546 2732
rect 2702 2728 2706 2732
rect 2718 2728 2722 2732
rect 3006 2728 3010 2732
rect 3118 2728 3122 2732
rect 3126 2728 3130 2732
rect 3214 2728 3218 2732
rect 3286 2728 3290 2732
rect 3630 2728 3634 2732
rect 3646 2728 3650 2732
rect 3726 2728 3730 2732
rect 3806 2728 3810 2732
rect 3894 2728 3898 2732
rect 4006 2728 4010 2732
rect 4182 2728 4186 2732
rect 4414 2728 4418 2732
rect 4462 2728 4466 2732
rect 4574 2728 4578 2732
rect 4822 2728 4826 2732
rect 4902 2728 4906 2732
rect 1430 2718 1434 2722
rect 1710 2718 1714 2722
rect 1934 2718 1938 2722
rect 2118 2718 2122 2722
rect 2838 2718 2842 2722
rect 2846 2718 2850 2722
rect 3070 2718 3074 2722
rect 3518 2718 3522 2722
rect 3838 2718 3842 2722
rect 3918 2718 3922 2722
rect 4398 2718 4402 2722
rect 4454 2718 4458 2722
rect 4702 2718 4706 2722
rect 854 2708 858 2712
rect 998 2708 1002 2712
rect 1350 2708 1354 2712
rect 2206 2708 2210 2712
rect 2838 2708 2842 2712
rect 3006 2708 3010 2712
rect 3142 2708 3146 2712
rect 3406 2708 3410 2712
rect 3894 2708 3898 2712
rect 4102 2708 4106 2712
rect 1050 2703 1054 2707
rect 1058 2703 1061 2707
rect 1061 2703 1062 2707
rect 1030 2698 1034 2702
rect 1582 2698 1586 2702
rect 2074 2703 2078 2707
rect 2082 2703 2085 2707
rect 2085 2703 2086 2707
rect 3098 2703 3102 2707
rect 3106 2703 3109 2707
rect 3109 2703 3110 2707
rect 4114 2703 4118 2707
rect 4122 2703 4125 2707
rect 4125 2703 4126 2707
rect 2054 2698 2058 2702
rect 2262 2698 2266 2702
rect 2350 2698 2354 2702
rect 2374 2698 2378 2702
rect 2614 2698 2618 2702
rect 3078 2698 3082 2702
rect 3118 2698 3122 2702
rect 3582 2698 3586 2702
rect 358 2688 362 2692
rect 582 2688 586 2692
rect 1838 2688 1842 2692
rect 2974 2688 2978 2692
rect 3662 2688 3666 2692
rect 4286 2688 4290 2692
rect 4326 2688 4330 2692
rect 4774 2688 4778 2692
rect 4998 2688 5002 2692
rect 206 2678 210 2682
rect 702 2678 706 2682
rect 1086 2678 1090 2682
rect 1366 2678 1370 2682
rect 1414 2678 1418 2682
rect 1446 2678 1450 2682
rect 1502 2678 1506 2682
rect 1750 2678 1754 2682
rect 1822 2678 1826 2682
rect 1838 2678 1842 2682
rect 1934 2678 1938 2682
rect 2246 2678 2250 2682
rect 2374 2678 2378 2682
rect 2494 2678 2498 2682
rect 2766 2678 2770 2682
rect 3054 2678 3058 2682
rect 3310 2678 3314 2682
rect 3534 2678 3538 2682
rect 3806 2678 3810 2682
rect 4366 2678 4370 2682
rect 4686 2678 4690 2682
rect 4982 2678 4986 2682
rect 270 2668 274 2672
rect 678 2668 682 2672
rect 1030 2668 1034 2672
rect 1246 2668 1250 2672
rect 1398 2668 1402 2672
rect 1510 2668 1514 2672
rect 1654 2668 1658 2672
rect 1998 2668 2002 2672
rect 2102 2668 2106 2672
rect 2374 2668 2378 2672
rect 2854 2668 2858 2672
rect 2878 2668 2882 2672
rect 3686 2668 3690 2672
rect 3886 2668 3890 2672
rect 3926 2668 3930 2672
rect 4566 2668 4570 2672
rect 4646 2668 4650 2672
rect 4670 2668 4674 2672
rect 4878 2668 4882 2672
rect 5070 2668 5074 2672
rect 190 2658 194 2662
rect 814 2658 818 2662
rect 830 2658 834 2662
rect 1166 2658 1170 2662
rect 1294 2658 1298 2662
rect 1382 2658 1386 2662
rect 1430 2658 1434 2662
rect 1798 2658 1802 2662
rect 1966 2658 1970 2662
rect 2078 2658 2082 2662
rect 2142 2658 2146 2662
rect 2278 2658 2282 2662
rect 2334 2658 2338 2662
rect 2358 2658 2362 2662
rect 2382 2658 2386 2662
rect 2702 2658 2706 2662
rect 2902 2658 2906 2662
rect 3038 2658 3042 2662
rect 3566 2658 3570 2662
rect 3590 2658 3594 2662
rect 3678 2658 3682 2662
rect 3942 2658 3946 2662
rect 4014 2658 4018 2662
rect 4286 2658 4290 2662
rect 5014 2658 5018 2662
rect 5142 2658 5146 2662
rect 5166 2658 5170 2662
rect 326 2648 330 2652
rect 582 2648 586 2652
rect 654 2648 658 2652
rect 894 2648 898 2652
rect 1150 2648 1154 2652
rect 1414 2648 1418 2652
rect 1462 2648 1466 2652
rect 2254 2648 2258 2652
rect 2294 2648 2298 2652
rect 2542 2648 2546 2652
rect 2782 2648 2786 2652
rect 3086 2648 3090 2652
rect 3174 2648 3178 2652
rect 3350 2648 3354 2652
rect 3542 2648 3546 2652
rect 3694 2648 3698 2652
rect 4014 2648 4018 2652
rect 4686 2648 4690 2652
rect 5166 2648 5170 2652
rect 5190 2648 5194 2652
rect 678 2638 682 2642
rect 2702 2638 2706 2642
rect 3318 2638 3322 2642
rect 3478 2638 3482 2642
rect 3566 2638 3570 2642
rect 3678 2638 3682 2642
rect 4182 2638 4186 2642
rect 4326 2638 4330 2642
rect 5110 2638 5114 2642
rect 670 2628 674 2632
rect 934 2628 938 2632
rect 998 2628 1002 2632
rect 1878 2628 1882 2632
rect 2070 2628 2074 2632
rect 2390 2628 2394 2632
rect 3550 2628 3554 2632
rect 3574 2628 3578 2632
rect 270 2618 274 2622
rect 590 2618 594 2622
rect 694 2618 698 2622
rect 918 2618 922 2622
rect 1214 2618 1218 2622
rect 1574 2618 1578 2622
rect 1606 2618 1610 2622
rect 2046 2618 2050 2622
rect 2454 2618 2458 2622
rect 2862 2618 2866 2622
rect 2878 2618 2882 2622
rect 3134 2618 3138 2622
rect 3478 2618 3482 2622
rect 3550 2618 3554 2622
rect 3782 2618 3786 2622
rect 4694 2618 4698 2622
rect 4934 2618 4938 2622
rect 5078 2618 5082 2622
rect 998 2608 1002 2612
rect 1174 2608 1178 2612
rect 1990 2608 1994 2612
rect 2054 2608 2058 2612
rect 2958 2608 2962 2612
rect 3230 2608 3234 2612
rect 3742 2608 3746 2612
rect 3790 2608 3794 2612
rect 4278 2608 4282 2612
rect 4446 2608 4450 2612
rect 4654 2608 4658 2612
rect 538 2603 542 2607
rect 546 2603 549 2607
rect 549 2603 550 2607
rect 1562 2603 1566 2607
rect 1570 2603 1573 2607
rect 1573 2603 1574 2607
rect 782 2598 786 2602
rect 1542 2598 1546 2602
rect 1710 2598 1714 2602
rect 2586 2603 2590 2607
rect 2594 2603 2597 2607
rect 2597 2603 2598 2607
rect 3610 2603 3614 2607
rect 3618 2603 3621 2607
rect 3621 2603 3622 2607
rect 4634 2603 4638 2607
rect 4642 2603 4645 2607
rect 4645 2603 4646 2607
rect 1862 2598 1866 2602
rect 1950 2598 1954 2602
rect 1974 2598 1978 2602
rect 2030 2598 2034 2602
rect 3350 2598 3354 2602
rect 3630 2598 3634 2602
rect 4862 2598 4866 2602
rect 1022 2588 1026 2592
rect 1846 2588 1850 2592
rect 1894 2588 1898 2592
rect 1934 2588 1938 2592
rect 2230 2588 2234 2592
rect 2334 2588 2338 2592
rect 2510 2588 2514 2592
rect 2534 2588 2538 2592
rect 3606 2588 3610 2592
rect 4222 2588 4226 2592
rect 1070 2578 1074 2582
rect 1158 2578 1162 2582
rect 1190 2578 1194 2582
rect 1846 2578 1850 2582
rect 2022 2578 2026 2582
rect 2246 2578 2250 2582
rect 2294 2578 2298 2582
rect 3534 2578 3538 2582
rect 3590 2578 3594 2582
rect 4742 2578 4746 2582
rect 5006 2578 5010 2582
rect 502 2568 506 2572
rect 574 2568 578 2572
rect 742 2568 746 2572
rect 782 2568 786 2572
rect 1134 2568 1138 2572
rect 1486 2568 1490 2572
rect 2566 2568 2570 2572
rect 2686 2568 2690 2572
rect 2814 2568 2818 2572
rect 2854 2568 2858 2572
rect 2918 2568 2922 2572
rect 3014 2568 3018 2572
rect 3206 2568 3210 2572
rect 3526 2568 3530 2572
rect 3558 2568 3562 2572
rect 3958 2568 3962 2572
rect 4494 2568 4498 2572
rect 4846 2568 4850 2572
rect 5118 2568 5122 2572
rect 142 2558 146 2562
rect 606 2558 610 2562
rect 1406 2558 1410 2562
rect 1526 2558 1530 2562
rect 1670 2558 1674 2562
rect 1838 2558 1842 2562
rect 2326 2558 2330 2562
rect 2886 2558 2890 2562
rect 2926 2558 2930 2562
rect 3334 2558 3338 2562
rect 3358 2558 3362 2562
rect 3454 2558 3458 2562
rect 3686 2558 3690 2562
rect 3750 2558 3754 2562
rect 3838 2558 3842 2562
rect 4150 2558 4154 2562
rect 4390 2558 4394 2562
rect 4598 2558 4602 2562
rect 5126 2558 5130 2562
rect 6 2548 10 2552
rect 422 2548 426 2552
rect 638 2548 642 2552
rect 790 2548 794 2552
rect 806 2548 810 2552
rect 846 2548 850 2552
rect 1158 2548 1162 2552
rect 1238 2548 1242 2552
rect 1422 2548 1426 2552
rect 1470 2548 1474 2552
rect 1486 2548 1490 2552
rect 1510 2548 1514 2552
rect 1670 2548 1674 2552
rect 1830 2548 1834 2552
rect 1854 2548 1858 2552
rect 1934 2548 1938 2552
rect 2014 2548 2018 2552
rect 2062 2548 2066 2552
rect 2086 2548 2090 2552
rect 2150 2548 2154 2552
rect 2334 2548 2338 2552
rect 2350 2548 2354 2552
rect 2398 2548 2402 2552
rect 2710 2548 2714 2552
rect 2742 2548 2746 2552
rect 2846 2548 2850 2552
rect 518 2538 522 2542
rect 582 2538 586 2542
rect 622 2538 626 2542
rect 1150 2538 1154 2542
rect 1198 2538 1202 2542
rect 1230 2538 1234 2542
rect 1430 2538 1434 2542
rect 1446 2538 1450 2542
rect 1494 2538 1498 2542
rect 1526 2538 1530 2542
rect 1662 2538 1666 2542
rect 1838 2538 1842 2542
rect 1894 2538 1898 2542
rect 1990 2538 1994 2542
rect 3630 2548 3634 2552
rect 4070 2548 4074 2552
rect 4126 2548 4130 2552
rect 4158 2548 4162 2552
rect 4526 2548 4530 2552
rect 4598 2548 4602 2552
rect 4766 2548 4770 2552
rect 5158 2548 5162 2552
rect 2110 2538 2114 2542
rect 2678 2538 2682 2542
rect 2702 2538 2706 2542
rect 3230 2538 3234 2542
rect 3286 2538 3290 2542
rect 3382 2538 3386 2542
rect 3454 2538 3458 2542
rect 3462 2538 3466 2542
rect 3846 2538 3850 2542
rect 4334 2538 4338 2542
rect 4358 2538 4362 2542
rect 4574 2538 4578 2542
rect 4974 2538 4978 2542
rect 5102 2538 5106 2542
rect 5126 2538 5130 2542
rect 502 2528 506 2532
rect 686 2528 690 2532
rect 1182 2528 1186 2532
rect 1238 2528 1242 2532
rect 1318 2528 1322 2532
rect 1822 2528 1826 2532
rect 1958 2528 1962 2532
rect 2150 2528 2154 2532
rect 2350 2528 2354 2532
rect 2694 2528 2698 2532
rect 2862 2528 2866 2532
rect 3006 2528 3010 2532
rect 3086 2528 3090 2532
rect 3206 2528 3210 2532
rect 3478 2528 3482 2532
rect 3582 2528 3586 2532
rect 3814 2528 3818 2532
rect 3950 2528 3954 2532
rect 4054 2528 4058 2532
rect 4366 2528 4370 2532
rect 4774 2528 4778 2532
rect 4790 2528 4794 2532
rect 5158 2528 5162 2532
rect 478 2518 482 2522
rect 518 2518 522 2522
rect 902 2518 906 2522
rect 918 2518 922 2522
rect 1934 2518 1938 2522
rect 1950 2518 1954 2522
rect 2046 2518 2050 2522
rect 2206 2518 2210 2522
rect 2342 2518 2346 2522
rect 2822 2518 2826 2522
rect 2902 2518 2906 2522
rect 3334 2518 3338 2522
rect 3526 2518 3530 2522
rect 4342 2518 4346 2522
rect 4998 2518 5002 2522
rect 14 2508 18 2512
rect 134 2508 138 2512
rect 630 2508 634 2512
rect 1118 2508 1122 2512
rect 1374 2508 1378 2512
rect 1398 2508 1402 2512
rect 1686 2508 1690 2512
rect 1726 2508 1730 2512
rect 1750 2508 1754 2512
rect 2030 2508 2034 2512
rect 2150 2508 2154 2512
rect 2382 2508 2386 2512
rect 2742 2508 2746 2512
rect 2806 2508 2810 2512
rect 3862 2508 3866 2512
rect 4158 2508 4162 2512
rect 4190 2508 4194 2512
rect 5038 2508 5042 2512
rect 1050 2503 1054 2507
rect 1058 2503 1061 2507
rect 1061 2503 1062 2507
rect 2074 2503 2078 2507
rect 2082 2503 2085 2507
rect 2085 2503 2086 2507
rect 3098 2503 3102 2507
rect 3106 2503 3109 2507
rect 3109 2503 3110 2507
rect 4114 2503 4118 2507
rect 4122 2503 4125 2507
rect 4125 2503 4126 2507
rect 2046 2498 2050 2502
rect 2214 2498 2218 2502
rect 2518 2498 2522 2502
rect 2934 2498 2938 2502
rect 3134 2498 3138 2502
rect 3310 2498 3314 2502
rect 3366 2498 3370 2502
rect 3430 2498 3434 2502
rect 6 2488 10 2492
rect 806 2488 810 2492
rect 1262 2488 1266 2492
rect 1542 2488 1546 2492
rect 1558 2488 1562 2492
rect 1742 2488 1746 2492
rect 1782 2488 1786 2492
rect 1806 2488 1810 2492
rect 3006 2488 3010 2492
rect 3062 2488 3066 2492
rect 3078 2488 3082 2492
rect 3214 2488 3218 2492
rect 3366 2488 3370 2492
rect 3382 2488 3386 2492
rect 3582 2488 3586 2492
rect 3670 2498 3674 2502
rect 3750 2498 3754 2502
rect 3974 2498 3978 2502
rect 4102 2498 4106 2502
rect 4430 2498 4434 2502
rect 4526 2498 4530 2502
rect 4534 2498 4538 2502
rect 4566 2498 4570 2502
rect 3702 2488 3706 2492
rect 3934 2488 3938 2492
rect 4086 2488 4090 2492
rect 4342 2488 4346 2492
rect 4454 2488 4458 2492
rect 4550 2488 4554 2492
rect 4742 2488 4746 2492
rect 5182 2488 5186 2492
rect 422 2478 426 2482
rect 550 2478 554 2482
rect 846 2478 850 2482
rect 854 2478 858 2482
rect 1158 2478 1162 2482
rect 1182 2478 1186 2482
rect 1654 2478 1658 2482
rect 1838 2478 1842 2482
rect 1886 2478 1890 2482
rect 1950 2478 1954 2482
rect 2182 2478 2186 2482
rect 2510 2478 2514 2482
rect 2646 2478 2650 2482
rect 2822 2478 2826 2482
rect 4270 2478 4274 2482
rect 4566 2478 4570 2482
rect 4838 2478 4842 2482
rect 4974 2478 4978 2482
rect 470 2468 474 2472
rect 118 2458 122 2462
rect 862 2468 866 2472
rect 958 2468 962 2472
rect 966 2468 970 2472
rect 1230 2468 1234 2472
rect 1318 2468 1322 2472
rect 1398 2468 1402 2472
rect 2246 2468 2250 2472
rect 2398 2468 2402 2472
rect 2422 2468 2426 2472
rect 2646 2468 2650 2472
rect 2710 2468 2714 2472
rect 2742 2468 2746 2472
rect 2846 2468 2850 2472
rect 3054 2468 3058 2472
rect 3134 2468 3138 2472
rect 3190 2468 3194 2472
rect 3238 2468 3242 2472
rect 3318 2468 3322 2472
rect 3950 2468 3954 2472
rect 3982 2468 3986 2472
rect 4038 2468 4042 2472
rect 4262 2468 4266 2472
rect 4358 2468 4362 2472
rect 4414 2468 4418 2472
rect 4430 2468 4434 2472
rect 4750 2468 4754 2472
rect 4854 2468 4858 2472
rect 4862 2468 4866 2472
rect 5110 2468 5114 2472
rect 406 2458 410 2462
rect 430 2458 434 2462
rect 598 2458 602 2462
rect 806 2458 810 2462
rect 838 2458 842 2462
rect 1254 2458 1258 2462
rect 1614 2458 1618 2462
rect 1790 2458 1794 2462
rect 1870 2458 1874 2462
rect 1878 2458 1882 2462
rect 1902 2458 1906 2462
rect 1942 2458 1946 2462
rect 2006 2458 2010 2462
rect 2198 2458 2202 2462
rect 2270 2458 2274 2462
rect 2334 2458 2338 2462
rect 2478 2458 2482 2462
rect 2614 2458 2618 2462
rect 2694 2458 2698 2462
rect 2766 2458 2770 2462
rect 702 2448 706 2452
rect 830 2448 834 2452
rect 1158 2448 1162 2452
rect 1262 2448 1266 2452
rect 1454 2448 1458 2452
rect 1806 2448 1810 2452
rect 1830 2448 1834 2452
rect 1966 2448 1970 2452
rect 2294 2448 2298 2452
rect 2318 2448 2322 2452
rect 2462 2448 2466 2452
rect 2798 2458 2802 2462
rect 3022 2458 3026 2462
rect 3262 2458 3266 2462
rect 3302 2458 3306 2462
rect 3390 2458 3394 2462
rect 3406 2458 3410 2462
rect 3462 2458 3466 2462
rect 3526 2458 3530 2462
rect 3622 2458 3626 2462
rect 3670 2458 3674 2462
rect 3982 2458 3986 2462
rect 4006 2458 4010 2462
rect 4094 2458 4098 2462
rect 4206 2458 4210 2462
rect 4438 2458 4442 2462
rect 4518 2458 4522 2462
rect 4734 2458 4738 2462
rect 4894 2458 4898 2462
rect 2606 2448 2610 2452
rect 2614 2448 2618 2452
rect 2838 2448 2842 2452
rect 3254 2448 3258 2452
rect 3614 2448 3618 2452
rect 3862 2448 3866 2452
rect 3950 2448 3954 2452
rect 4342 2448 4346 2452
rect 4550 2448 4554 2452
rect 4702 2448 4706 2452
rect 5022 2448 5026 2452
rect 5174 2448 5178 2452
rect 1214 2438 1218 2442
rect 1238 2438 1242 2442
rect 1262 2438 1266 2442
rect 1558 2438 1562 2442
rect 1878 2438 1882 2442
rect 1902 2438 1906 2442
rect 1990 2438 1994 2442
rect 2238 2438 2242 2442
rect 2398 2438 2402 2442
rect 2406 2438 2410 2442
rect 3302 2438 3306 2442
rect 3350 2438 3354 2442
rect 3382 2438 3386 2442
rect 3422 2438 3426 2442
rect 3614 2438 3618 2442
rect 3718 2438 3722 2442
rect 3766 2438 3770 2442
rect 3790 2438 3794 2442
rect 3910 2438 3914 2442
rect 4486 2438 4490 2442
rect 5126 2438 5130 2442
rect 630 2428 634 2432
rect 846 2428 850 2432
rect 1374 2428 1378 2432
rect 1390 2428 1394 2432
rect 1750 2428 1754 2432
rect 1782 2428 1786 2432
rect 1966 2428 1970 2432
rect 2174 2428 2178 2432
rect 2182 2428 2186 2432
rect 2614 2428 2618 2432
rect 3950 2428 3954 2432
rect 3974 2428 3978 2432
rect 3990 2428 3994 2432
rect 4942 2428 4946 2432
rect 5094 2428 5098 2432
rect 718 2418 722 2422
rect 1374 2418 1378 2422
rect 1646 2418 1650 2422
rect 1870 2418 1874 2422
rect 3126 2418 3130 2422
rect 3414 2418 3418 2422
rect 3422 2418 3426 2422
rect 3486 2418 3490 2422
rect 3590 2418 3594 2422
rect 3606 2418 3610 2422
rect 3638 2418 3642 2422
rect 3694 2418 3698 2422
rect 3790 2418 3794 2422
rect 4222 2418 4226 2422
rect 5182 2418 5186 2422
rect 798 2408 802 2412
rect 998 2408 1002 2412
rect 1110 2408 1114 2412
rect 1254 2408 1258 2412
rect 1414 2408 1418 2412
rect 1686 2408 1690 2412
rect 1838 2408 1842 2412
rect 2382 2408 2386 2412
rect 2550 2408 2554 2412
rect 2654 2408 2658 2412
rect 3030 2408 3034 2412
rect 3110 2408 3114 2412
rect 3158 2408 3162 2412
rect 3446 2408 3450 2412
rect 4182 2408 4186 2412
rect 4654 2408 4658 2412
rect 538 2403 542 2407
rect 546 2403 549 2407
rect 549 2403 550 2407
rect 1562 2403 1566 2407
rect 1570 2403 1573 2407
rect 1573 2403 1574 2407
rect 2586 2403 2590 2407
rect 2594 2403 2597 2407
rect 2597 2403 2598 2407
rect 3610 2403 3614 2407
rect 3618 2403 3621 2407
rect 3621 2403 3622 2407
rect 4634 2403 4638 2407
rect 4642 2403 4645 2407
rect 4645 2403 4646 2407
rect 622 2398 626 2402
rect 630 2398 634 2402
rect 1806 2398 1810 2402
rect 2262 2398 2266 2402
rect 2286 2398 2290 2402
rect 3182 2398 3186 2402
rect 3198 2398 3202 2402
rect 3302 2398 3306 2402
rect 3806 2398 3810 2402
rect 4070 2398 4074 2402
rect 5030 2398 5034 2402
rect 470 2388 474 2392
rect 846 2388 850 2392
rect 1174 2388 1178 2392
rect 1606 2388 1610 2392
rect 1750 2388 1754 2392
rect 1918 2388 1922 2392
rect 2142 2388 2146 2392
rect 2182 2388 2186 2392
rect 3494 2388 3498 2392
rect 3806 2388 3810 2392
rect 3950 2388 3954 2392
rect 4886 2388 4890 2392
rect 742 2378 746 2382
rect 1278 2378 1282 2382
rect 1318 2378 1322 2382
rect 1350 2378 1354 2382
rect 1502 2378 1506 2382
rect 2174 2378 2178 2382
rect 3790 2378 3794 2382
rect 4238 2378 4242 2382
rect 902 2368 906 2372
rect 1262 2368 1266 2372
rect 1366 2368 1370 2372
rect 1878 2368 1882 2372
rect 1910 2368 1914 2372
rect 1934 2368 1938 2372
rect 2006 2368 2010 2372
rect 2046 2368 2050 2372
rect 2086 2368 2090 2372
rect 2166 2368 2170 2372
rect 2246 2368 2250 2372
rect 2502 2368 2506 2372
rect 2566 2368 2570 2372
rect 2630 2368 2634 2372
rect 2710 2368 2714 2372
rect 3118 2368 3122 2372
rect 3230 2368 3234 2372
rect 4182 2368 4186 2372
rect 5046 2368 5050 2372
rect 5094 2368 5098 2372
rect 598 2358 602 2362
rect 894 2358 898 2362
rect 958 2358 962 2362
rect 1126 2358 1130 2362
rect 1166 2358 1170 2362
rect 1230 2358 1234 2362
rect 2142 2358 2146 2362
rect 2390 2358 2394 2362
rect 2510 2358 2514 2362
rect 2822 2358 2826 2362
rect 2934 2358 2938 2362
rect 3190 2358 3194 2362
rect 3198 2358 3202 2362
rect 3246 2358 3250 2362
rect 3358 2358 3362 2362
rect 3470 2358 3474 2362
rect 3766 2358 3770 2362
rect 3806 2358 3810 2362
rect 4534 2358 4538 2362
rect 4942 2358 4946 2362
rect 6 2348 10 2352
rect 94 2348 98 2352
rect 526 2348 530 2352
rect 646 2348 650 2352
rect 934 2348 938 2352
rect 1222 2348 1226 2352
rect 1342 2348 1346 2352
rect 1510 2348 1514 2352
rect 1718 2348 1722 2352
rect 1750 2348 1754 2352
rect 1838 2348 1842 2352
rect 2302 2348 2306 2352
rect 2318 2348 2322 2352
rect 2454 2348 2458 2352
rect 3174 2348 3178 2352
rect 3294 2348 3298 2352
rect 3398 2348 3402 2352
rect 3414 2348 3418 2352
rect 3598 2348 3602 2352
rect 3830 2348 3834 2352
rect 4134 2348 4138 2352
rect 4182 2348 4186 2352
rect 4198 2348 4202 2352
rect 4374 2348 4378 2352
rect 4470 2348 4474 2352
rect 4766 2348 4770 2352
rect 4902 2348 4906 2352
rect 4926 2348 4930 2352
rect 5054 2348 5058 2352
rect 470 2338 474 2342
rect 510 2338 514 2342
rect 582 2338 586 2342
rect 814 2338 818 2342
rect 870 2338 874 2342
rect 1486 2338 1490 2342
rect 1798 2338 1802 2342
rect 1846 2338 1850 2342
rect 2134 2338 2138 2342
rect 2310 2338 2314 2342
rect 2374 2338 2378 2342
rect 2582 2338 2586 2342
rect 2622 2338 2626 2342
rect 2670 2338 2674 2342
rect 2878 2338 2882 2342
rect 3054 2338 3058 2342
rect 3318 2338 3322 2342
rect 3502 2338 3506 2342
rect 3518 2338 3522 2342
rect 3726 2338 3730 2342
rect 3950 2338 3954 2342
rect 4030 2338 4034 2342
rect 4414 2338 4418 2342
rect 4702 2338 4706 2342
rect 5110 2338 5114 2342
rect 5126 2338 5130 2342
rect 6 2328 10 2332
rect 502 2328 506 2332
rect 934 2328 938 2332
rect 1382 2328 1386 2332
rect 1406 2328 1410 2332
rect 1694 2328 1698 2332
rect 1822 2328 1826 2332
rect 1838 2328 1842 2332
rect 1902 2328 1906 2332
rect 1918 2328 1922 2332
rect 2238 2328 2242 2332
rect 2542 2328 2546 2332
rect 2822 2328 2826 2332
rect 3134 2328 3138 2332
rect 3414 2328 3418 2332
rect 3454 2328 3458 2332
rect 3550 2328 3554 2332
rect 3758 2328 3762 2332
rect 4262 2328 4266 2332
rect 4302 2328 4306 2332
rect 382 2318 386 2322
rect 782 2318 786 2322
rect 806 2318 810 2322
rect 814 2318 818 2322
rect 1838 2318 1842 2322
rect 1934 2318 1938 2322
rect 2006 2318 2010 2322
rect 2334 2318 2338 2322
rect 2814 2318 2818 2322
rect 3278 2318 3282 2322
rect 3422 2318 3426 2322
rect 4246 2318 4250 2322
rect 4310 2318 4314 2322
rect 4326 2318 4330 2322
rect 4358 2318 4362 2322
rect 4382 2318 4386 2322
rect 4638 2318 4642 2322
rect 4822 2318 4826 2322
rect 4942 2318 4946 2322
rect 5030 2318 5034 2322
rect 798 2308 802 2312
rect 1166 2308 1170 2312
rect 1262 2308 1266 2312
rect 1526 2308 1530 2312
rect 1598 2308 1602 2312
rect 1638 2308 1642 2312
rect 1662 2308 1666 2312
rect 1878 2308 1882 2312
rect 2782 2308 2786 2312
rect 2910 2308 2914 2312
rect 2942 2308 2946 2312
rect 3070 2308 3074 2312
rect 3478 2308 3482 2312
rect 3614 2308 3618 2312
rect 4238 2308 4242 2312
rect 4390 2308 4394 2312
rect 4694 2308 4698 2312
rect 1050 2303 1054 2307
rect 1058 2303 1061 2307
rect 1061 2303 1062 2307
rect 2074 2303 2078 2307
rect 2082 2303 2085 2307
rect 2085 2303 2086 2307
rect 3098 2303 3102 2307
rect 3106 2303 3109 2307
rect 3109 2303 3110 2307
rect 4114 2303 4118 2307
rect 4122 2303 4125 2307
rect 4125 2303 4126 2307
rect 902 2298 906 2302
rect 1350 2298 1354 2302
rect 1406 2298 1410 2302
rect 1854 2298 1858 2302
rect 2134 2298 2138 2302
rect 2158 2298 2162 2302
rect 2198 2298 2202 2302
rect 2206 2298 2210 2302
rect 2446 2298 2450 2302
rect 2814 2298 2818 2302
rect 3150 2298 3154 2302
rect 3342 2298 3346 2302
rect 3494 2298 3498 2302
rect 3526 2298 3530 2302
rect 3558 2298 3562 2302
rect 3686 2298 3690 2302
rect 4662 2298 4666 2302
rect 5062 2298 5066 2302
rect 982 2288 986 2292
rect 1654 2288 1658 2292
rect 1886 2288 1890 2292
rect 2102 2288 2106 2292
rect 2270 2288 2274 2292
rect 2286 2288 2290 2292
rect 2934 2288 2938 2292
rect 2958 2288 2962 2292
rect 3758 2288 3762 2292
rect 4158 2288 4162 2292
rect 4206 2288 4210 2292
rect 4350 2288 4354 2292
rect 4534 2288 4538 2292
rect 5142 2288 5146 2292
rect 214 2278 218 2282
rect 1118 2278 1122 2282
rect 1254 2278 1258 2282
rect 1334 2278 1338 2282
rect 1678 2278 1682 2282
rect 1918 2278 1922 2282
rect 1998 2278 2002 2282
rect 2238 2278 2242 2282
rect 2542 2278 2546 2282
rect 2742 2278 2746 2282
rect 2910 2278 2914 2282
rect 2998 2278 3002 2282
rect 3222 2278 3226 2282
rect 3238 2278 3242 2282
rect 3334 2278 3338 2282
rect 4598 2278 4602 2282
rect 4646 2278 4650 2282
rect 4838 2278 4842 2282
rect 4886 2278 4890 2282
rect 5134 2278 5138 2282
rect 302 2268 306 2272
rect 870 2268 874 2272
rect 1302 2268 1306 2272
rect 1534 2268 1538 2272
rect 1614 2268 1618 2272
rect 1670 2268 1674 2272
rect 1726 2268 1730 2272
rect 1750 2268 1754 2272
rect 1790 2268 1794 2272
rect 1958 2268 1962 2272
rect 1966 2268 1970 2272
rect 2150 2268 2154 2272
rect 2270 2268 2274 2272
rect 2422 2268 2426 2272
rect 2950 2268 2954 2272
rect 2966 2268 2970 2272
rect 3046 2268 3050 2272
rect 3326 2268 3330 2272
rect 3374 2268 3378 2272
rect 4926 2268 4930 2272
rect 5150 2268 5154 2272
rect 590 2258 594 2262
rect 622 2258 626 2262
rect 654 2258 658 2262
rect 862 2258 866 2262
rect 942 2258 946 2262
rect 1190 2258 1194 2262
rect 1198 2258 1202 2262
rect 1222 2258 1226 2262
rect 1502 2258 1506 2262
rect 1734 2258 1738 2262
rect 1894 2258 1898 2262
rect 2062 2258 2066 2262
rect 2142 2258 2146 2262
rect 2454 2258 2458 2262
rect 2694 2258 2698 2262
rect 3078 2258 3082 2262
rect 3102 2258 3106 2262
rect 3414 2258 3418 2262
rect 3750 2258 3754 2262
rect 4102 2258 4106 2262
rect 4358 2258 4362 2262
rect 4462 2258 4466 2262
rect 4558 2258 4562 2262
rect 4702 2258 4706 2262
rect 4886 2258 4890 2262
rect 5158 2258 5162 2262
rect 446 2248 450 2252
rect 1814 2248 1818 2252
rect 2070 2248 2074 2252
rect 2102 2248 2106 2252
rect 2150 2248 2154 2252
rect 2230 2248 2234 2252
rect 2350 2248 2354 2252
rect 3174 2248 3178 2252
rect 3630 2248 3634 2252
rect 3710 2248 3714 2252
rect 3782 2248 3786 2252
rect 3982 2248 3986 2252
rect 4118 2248 4122 2252
rect 4286 2248 4290 2252
rect 4702 2248 4706 2252
rect 4750 2248 4754 2252
rect 1350 2238 1354 2242
rect 1606 2238 1610 2242
rect 1750 2238 1754 2242
rect 2094 2238 2098 2242
rect 2118 2238 2122 2242
rect 2166 2238 2170 2242
rect 3046 2238 3050 2242
rect 3366 2238 3370 2242
rect 3510 2238 3514 2242
rect 3758 2238 3762 2242
rect 3806 2238 3810 2242
rect 3870 2238 3874 2242
rect 3902 2238 3906 2242
rect 870 2228 874 2232
rect 910 2228 914 2232
rect 958 2228 962 2232
rect 2078 2228 2082 2232
rect 2206 2228 2210 2232
rect 2494 2228 2498 2232
rect 2846 2228 2850 2232
rect 3102 2228 3106 2232
rect 3118 2228 3122 2232
rect 3286 2228 3290 2232
rect 3734 2228 3738 2232
rect 3862 2228 3866 2232
rect 3942 2228 3946 2232
rect 4230 2228 4234 2232
rect 4414 2228 4418 2232
rect 438 2218 442 2222
rect 830 2218 834 2222
rect 1822 2218 1826 2222
rect 1830 2218 1834 2222
rect 1886 2218 1890 2222
rect 1926 2218 1930 2222
rect 1990 2218 1994 2222
rect 2054 2218 2058 2222
rect 2118 2218 2122 2222
rect 2150 2218 2154 2222
rect 2358 2218 2362 2222
rect 2654 2218 2658 2222
rect 2742 2218 2746 2222
rect 2790 2218 2794 2222
rect 3014 2218 3018 2222
rect 3470 2218 3474 2222
rect 3806 2218 3810 2222
rect 4598 2218 4602 2222
rect 446 2208 450 2212
rect 694 2208 698 2212
rect 1542 2208 1546 2212
rect 1718 2208 1722 2212
rect 1950 2208 1954 2212
rect 1966 2208 1970 2212
rect 2486 2208 2490 2212
rect 3126 2208 3130 2212
rect 3158 2208 3162 2212
rect 3462 2208 3466 2212
rect 3582 2208 3586 2212
rect 3886 2208 3890 2212
rect 4206 2208 4210 2212
rect 4838 2208 4842 2212
rect 538 2203 542 2207
rect 546 2203 549 2207
rect 549 2203 550 2207
rect 1562 2203 1566 2207
rect 1570 2203 1573 2207
rect 1573 2203 1574 2207
rect 2586 2203 2590 2207
rect 2594 2203 2597 2207
rect 2597 2203 2598 2207
rect 3610 2203 3614 2207
rect 3618 2203 3621 2207
rect 3621 2203 3622 2207
rect 4634 2203 4638 2207
rect 4642 2203 4645 2207
rect 4645 2203 4646 2207
rect 814 2198 818 2202
rect 1246 2198 1250 2202
rect 1582 2198 1586 2202
rect 1814 2198 1818 2202
rect 1918 2198 1922 2202
rect 1990 2198 1994 2202
rect 2206 2198 2210 2202
rect 2486 2198 2490 2202
rect 3310 2198 3314 2202
rect 3470 2198 3474 2202
rect 4030 2198 4034 2202
rect 4038 2198 4042 2202
rect 4294 2198 4298 2202
rect 4830 2198 4834 2202
rect 838 2188 842 2192
rect 862 2188 866 2192
rect 1958 2188 1962 2192
rect 2070 2188 2074 2192
rect 2078 2188 2082 2192
rect 2270 2188 2274 2192
rect 2582 2188 2586 2192
rect 3214 2188 3218 2192
rect 3510 2188 3514 2192
rect 3822 2188 3826 2192
rect 3926 2188 3930 2192
rect 4726 2188 4730 2192
rect 4774 2188 4778 2192
rect 718 2178 722 2182
rect 1838 2178 1842 2182
rect 1910 2178 1914 2182
rect 1934 2178 1938 2182
rect 2030 2178 2034 2182
rect 2158 2178 2162 2182
rect 2230 2178 2234 2182
rect 3774 2178 3778 2182
rect 4742 2178 4746 2182
rect 382 2168 386 2172
rect 1430 2168 1434 2172
rect 1790 2168 1794 2172
rect 1934 2168 1938 2172
rect 2046 2168 2050 2172
rect 2286 2168 2290 2172
rect 2294 2168 2298 2172
rect 2342 2168 2346 2172
rect 2462 2168 2466 2172
rect 2526 2168 2530 2172
rect 2806 2168 2810 2172
rect 2990 2168 2994 2172
rect 3582 2168 3586 2172
rect 3694 2168 3698 2172
rect 3822 2168 3826 2172
rect 4246 2168 4250 2172
rect 4318 2168 4322 2172
rect 4486 2168 4490 2172
rect 4550 2168 4554 2172
rect 4854 2168 4858 2172
rect 438 2158 442 2162
rect 606 2158 610 2162
rect 630 2158 634 2162
rect 646 2158 650 2162
rect 846 2158 850 2162
rect 1126 2158 1130 2162
rect 1318 2158 1322 2162
rect 1390 2158 1394 2162
rect 1414 2158 1418 2162
rect 1430 2158 1434 2162
rect 1662 2158 1666 2162
rect 1790 2158 1794 2162
rect 1990 2158 1994 2162
rect 2062 2158 2066 2162
rect 2150 2158 2154 2162
rect 2182 2158 2186 2162
rect 2198 2158 2202 2162
rect 2302 2158 2306 2162
rect 2446 2158 2450 2162
rect 2470 2158 2474 2162
rect 2838 2158 2842 2162
rect 3038 2158 3042 2162
rect 3110 2158 3114 2162
rect 3246 2158 3250 2162
rect 3270 2158 3274 2162
rect 3342 2158 3346 2162
rect 3558 2158 3562 2162
rect 3566 2158 3570 2162
rect 3630 2158 3634 2162
rect 3654 2158 3658 2162
rect 3758 2158 3762 2162
rect 4742 2158 4746 2162
rect 4798 2158 4802 2162
rect 4862 2158 4866 2162
rect 4902 2158 4906 2162
rect 94 2148 98 2152
rect 286 2148 290 2152
rect 694 2148 698 2152
rect 710 2148 714 2152
rect 958 2148 962 2152
rect 1286 2148 1290 2152
rect 1366 2148 1370 2152
rect 1406 2148 1410 2152
rect 1718 2148 1722 2152
rect 2174 2148 2178 2152
rect 2270 2148 2274 2152
rect 2414 2148 2418 2152
rect 2926 2148 2930 2152
rect 3350 2148 3354 2152
rect 3534 2148 3538 2152
rect 3598 2148 3602 2152
rect 3694 2148 3698 2152
rect 3742 2148 3746 2152
rect 3990 2148 3994 2152
rect 4022 2148 4026 2152
rect 4078 2148 4082 2152
rect 4150 2148 4154 2152
rect 4222 2148 4226 2152
rect 4350 2148 4354 2152
rect 4726 2148 4730 2152
rect 4790 2148 4794 2152
rect 4822 2148 4826 2152
rect 4934 2148 4938 2152
rect 878 2138 882 2142
rect 910 2138 914 2142
rect 934 2138 938 2142
rect 1126 2138 1130 2142
rect 1366 2138 1370 2142
rect 1662 2138 1666 2142
rect 1798 2138 1802 2142
rect 1942 2138 1946 2142
rect 1950 2138 1954 2142
rect 2102 2138 2106 2142
rect 2446 2138 2450 2142
rect 3038 2138 3042 2142
rect 3046 2138 3050 2142
rect 3526 2138 3530 2142
rect 3654 2138 3658 2142
rect 3854 2138 3858 2142
rect 3942 2138 3946 2142
rect 4174 2138 4178 2142
rect 4646 2138 4650 2142
rect 4854 2138 4858 2142
rect 638 2128 642 2132
rect 782 2128 786 2132
rect 830 2128 834 2132
rect 1270 2128 1274 2132
rect 1718 2128 1722 2132
rect 1742 2128 1746 2132
rect 1926 2128 1930 2132
rect 1974 2128 1978 2132
rect 2094 2128 2098 2132
rect 2534 2128 2538 2132
rect 2950 2128 2954 2132
rect 3054 2128 3058 2132
rect 3958 2128 3962 2132
rect 4038 2128 4042 2132
rect 4374 2128 4378 2132
rect 4526 2128 4530 2132
rect 4566 2128 4570 2132
rect 4790 2128 4794 2132
rect 5070 2128 5074 2132
rect 286 2118 290 2122
rect 566 2118 570 2122
rect 758 2118 762 2122
rect 870 2118 874 2122
rect 1470 2118 1474 2122
rect 1558 2118 1562 2122
rect 1726 2118 1730 2122
rect 1814 2118 1818 2122
rect 1878 2118 1882 2122
rect 1910 2118 1914 2122
rect 2142 2118 2146 2122
rect 2670 2118 2674 2122
rect 3014 2118 3018 2122
rect 3078 2118 3082 2122
rect 3134 2118 3138 2122
rect 3302 2118 3306 2122
rect 3318 2118 3322 2122
rect 3582 2118 3586 2122
rect 4382 2118 4386 2122
rect 4950 2118 4954 2122
rect 222 2108 226 2112
rect 446 2108 450 2112
rect 502 2108 506 2112
rect 806 2108 810 2112
rect 1126 2108 1130 2112
rect 1174 2108 1178 2112
rect 1334 2108 1338 2112
rect 1398 2108 1402 2112
rect 1630 2108 1634 2112
rect 1678 2108 1682 2112
rect 1702 2108 1706 2112
rect 2254 2108 2258 2112
rect 2310 2108 2314 2112
rect 3126 2108 3130 2112
rect 3150 2108 3154 2112
rect 3198 2108 3202 2112
rect 3286 2108 3290 2112
rect 3486 2108 3490 2112
rect 3710 2108 3714 2112
rect 1050 2103 1054 2107
rect 1058 2103 1061 2107
rect 1061 2103 1062 2107
rect 2074 2103 2078 2107
rect 2082 2103 2085 2107
rect 2085 2103 2086 2107
rect 302 2098 306 2102
rect 1078 2098 1082 2102
rect 1870 2098 1874 2102
rect 1934 2098 1938 2102
rect 1942 2098 1946 2102
rect 2182 2098 2186 2102
rect 2278 2098 2282 2102
rect 3098 2103 3102 2107
rect 3106 2103 3109 2107
rect 3109 2103 3110 2107
rect 4114 2103 4118 2107
rect 4122 2103 4125 2107
rect 4125 2103 4126 2107
rect 2998 2098 3002 2102
rect 3646 2098 3650 2102
rect 4342 2098 4346 2102
rect 4494 2098 4498 2102
rect 4934 2098 4938 2102
rect 5174 2098 5178 2102
rect 70 2088 74 2092
rect 214 2088 218 2092
rect 974 2088 978 2092
rect 1190 2088 1194 2092
rect 1470 2088 1474 2092
rect 1894 2088 1898 2092
rect 1926 2088 1930 2092
rect 2038 2088 2042 2092
rect 2390 2088 2394 2092
rect 3414 2088 3418 2092
rect 3534 2088 3538 2092
rect 4902 2088 4906 2092
rect 166 2078 170 2082
rect 742 2078 746 2082
rect 1038 2078 1042 2082
rect 1102 2078 1106 2082
rect 1454 2078 1458 2082
rect 1638 2078 1642 2082
rect 1910 2078 1914 2082
rect 2110 2078 2114 2082
rect 2118 2078 2122 2082
rect 2254 2078 2258 2082
rect 2350 2078 2354 2082
rect 3126 2078 3130 2082
rect 3462 2078 3466 2082
rect 3502 2078 3506 2082
rect 3910 2078 3914 2082
rect 3942 2078 3946 2082
rect 4134 2078 4138 2082
rect 4478 2078 4482 2082
rect 4814 2078 4818 2082
rect 5174 2078 5178 2082
rect 1302 2068 1306 2072
rect 1342 2068 1346 2072
rect 1486 2068 1490 2072
rect 1502 2068 1506 2072
rect 1582 2068 1586 2072
rect 1974 2068 1978 2072
rect 2006 2068 2010 2072
rect 2102 2068 2106 2072
rect 2150 2068 2154 2072
rect 2318 2068 2322 2072
rect 2622 2068 2626 2072
rect 2790 2068 2794 2072
rect 2894 2068 2898 2072
rect 3446 2068 3450 2072
rect 3518 2068 3522 2072
rect 4062 2068 4066 2072
rect 4198 2068 4202 2072
rect 4526 2068 4530 2072
rect 4742 2068 4746 2072
rect 4798 2068 4802 2072
rect 5006 2068 5010 2072
rect 5062 2068 5066 2072
rect 5094 2068 5098 2072
rect 5110 2068 5114 2072
rect 134 2058 138 2062
rect 438 2058 442 2062
rect 750 2058 754 2062
rect 982 2058 986 2062
rect 998 2058 1002 2062
rect 1118 2058 1122 2062
rect 1174 2058 1178 2062
rect 1566 2058 1570 2062
rect 1614 2058 1618 2062
rect 1686 2058 1690 2062
rect 1894 2058 1898 2062
rect 2710 2058 2714 2062
rect 2934 2058 2938 2062
rect 3038 2058 3042 2062
rect 3174 2058 3178 2062
rect 3398 2058 3402 2062
rect 3430 2058 3434 2062
rect 3470 2058 3474 2062
rect 4406 2058 4410 2062
rect 4782 2058 4786 2062
rect 5038 2058 5042 2062
rect 5190 2058 5194 2062
rect 374 2048 378 2052
rect 486 2048 490 2052
rect 934 2048 938 2052
rect 1742 2048 1746 2052
rect 1830 2048 1834 2052
rect 2078 2048 2082 2052
rect 2270 2048 2274 2052
rect 2662 2048 2666 2052
rect 2830 2048 2834 2052
rect 3118 2048 3122 2052
rect 3262 2048 3266 2052
rect 3294 2048 3298 2052
rect 3486 2048 3490 2052
rect 4390 2048 4394 2052
rect 4462 2048 4466 2052
rect 4574 2048 4578 2052
rect 5070 2048 5074 2052
rect 5166 2048 5170 2052
rect 526 2038 530 2042
rect 958 2038 962 2042
rect 1078 2038 1082 2042
rect 1094 2038 1098 2042
rect 1166 2038 1170 2042
rect 1190 2038 1194 2042
rect 1278 2038 1282 2042
rect 1630 2038 1634 2042
rect 1758 2038 1762 2042
rect 2734 2038 2738 2042
rect 2854 2038 2858 2042
rect 3318 2038 3322 2042
rect 3422 2038 3426 2042
rect 3478 2038 3482 2042
rect 3854 2038 3858 2042
rect 3982 2038 3986 2042
rect 4110 2038 4114 2042
rect 4118 2038 4122 2042
rect 5166 2038 5170 2042
rect 814 2028 818 2032
rect 1182 2028 1186 2032
rect 1206 2028 1210 2032
rect 1270 2028 1274 2032
rect 2030 2028 2034 2032
rect 2102 2028 2106 2032
rect 3678 2028 3682 2032
rect 4006 2028 4010 2032
rect 4190 2028 4194 2032
rect 4238 2028 4242 2032
rect 5086 2028 5090 2032
rect 1094 2018 1098 2022
rect 1110 2018 1114 2022
rect 1270 2018 1274 2022
rect 1686 2018 1690 2022
rect 2358 2018 2362 2022
rect 2822 2018 2826 2022
rect 2862 2018 2866 2022
rect 3286 2018 3290 2022
rect 3766 2018 3770 2022
rect 4086 2018 4090 2022
rect 4134 2018 4138 2022
rect 4166 2018 4170 2022
rect 966 2008 970 2012
rect 990 2008 994 2012
rect 1550 2008 1554 2012
rect 1798 2008 1802 2012
rect 2118 2008 2122 2012
rect 2334 2008 2338 2012
rect 2494 2008 2498 2012
rect 2550 2008 2554 2012
rect 2790 2008 2794 2012
rect 3342 2008 3346 2012
rect 3598 2008 3602 2012
rect 4086 2008 4090 2012
rect 4406 2008 4410 2012
rect 4478 2008 4482 2012
rect 5102 2008 5106 2012
rect 538 2003 542 2007
rect 546 2003 549 2007
rect 549 2003 550 2007
rect 1562 2003 1566 2007
rect 1570 2003 1573 2007
rect 1573 2003 1574 2007
rect 2586 2003 2590 2007
rect 2594 2003 2597 2007
rect 2597 2003 2598 2007
rect 3610 2003 3614 2007
rect 3618 2003 3621 2007
rect 3621 2003 3622 2007
rect 4634 2003 4638 2007
rect 4642 2003 4645 2007
rect 4645 2003 4646 2007
rect 822 1998 826 2002
rect 1950 1998 1954 2002
rect 1966 1998 1970 2002
rect 2310 1998 2314 2002
rect 2574 1998 2578 2002
rect 3454 1998 3458 2002
rect 3462 1998 3466 2002
rect 4022 1998 4026 2002
rect 4134 1998 4138 2002
rect 4302 1998 4306 2002
rect 4534 1998 4538 2002
rect 4542 1998 4546 2002
rect 5022 1998 5026 2002
rect 1342 1988 1346 1992
rect 1606 1988 1610 1992
rect 1710 1988 1714 1992
rect 1990 1988 1994 1992
rect 2014 1988 2018 1992
rect 2118 1988 2122 1992
rect 2262 1988 2266 1992
rect 2406 1988 2410 1992
rect 2430 1988 2434 1992
rect 2694 1988 2698 1992
rect 2798 1988 2802 1992
rect 4326 1988 4330 1992
rect 1550 1978 1554 1982
rect 1742 1978 1746 1982
rect 1894 1978 1898 1982
rect 2006 1978 2010 1982
rect 2246 1978 2250 1982
rect 2278 1978 2282 1982
rect 2870 1978 2874 1982
rect 3774 1978 3778 1982
rect 5174 1978 5178 1982
rect 878 1968 882 1972
rect 1502 1968 1506 1972
rect 1534 1968 1538 1972
rect 2062 1968 2066 1972
rect 2534 1968 2538 1972
rect 2630 1968 2634 1972
rect 2982 1968 2986 1972
rect 3014 1968 3018 1972
rect 3198 1968 3202 1972
rect 3222 1968 3226 1972
rect 3862 1968 3866 1972
rect 4182 1968 4186 1972
rect 4318 1968 4322 1972
rect 4494 1968 4498 1972
rect 5086 1968 5090 1972
rect 294 1958 298 1962
rect 302 1958 306 1962
rect 462 1958 466 1962
rect 894 1958 898 1962
rect 942 1958 946 1962
rect 966 1958 970 1962
rect 1102 1958 1106 1962
rect 1150 1958 1154 1962
rect 1302 1958 1306 1962
rect 1350 1958 1354 1962
rect 1838 1958 1842 1962
rect 2502 1958 2506 1962
rect 2958 1958 2962 1962
rect 3326 1958 3330 1962
rect 3430 1958 3434 1962
rect 3462 1958 3466 1962
rect 3574 1958 3578 1962
rect 3758 1958 3762 1962
rect 3854 1958 3858 1962
rect 4078 1958 4082 1962
rect 4150 1958 4154 1962
rect 4454 1958 4458 1962
rect 4494 1958 4498 1962
rect 4750 1958 4754 1962
rect 5166 1958 5170 1962
rect 478 1948 482 1952
rect 614 1948 618 1952
rect 774 1948 778 1952
rect 974 1948 978 1952
rect 1030 1948 1034 1952
rect 1046 1948 1050 1952
rect 1086 1948 1090 1952
rect 1142 1948 1146 1952
rect 1310 1948 1314 1952
rect 1334 1948 1338 1952
rect 1774 1948 1778 1952
rect 2022 1948 2026 1952
rect 2078 1948 2082 1952
rect 2198 1948 2202 1952
rect 2238 1948 2242 1952
rect 2310 1948 2314 1952
rect 2470 1948 2474 1952
rect 2494 1948 2498 1952
rect 2566 1948 2570 1952
rect 2702 1948 2706 1952
rect 3566 1948 3570 1952
rect 3662 1948 3666 1952
rect 3670 1948 3674 1952
rect 3782 1948 3786 1952
rect 3878 1948 3882 1952
rect 4030 1948 4034 1952
rect 4086 1948 4090 1952
rect 4262 1948 4266 1952
rect 4646 1948 4650 1952
rect 4702 1948 4706 1952
rect 4742 1948 4746 1952
rect 4814 1948 4818 1952
rect 558 1938 562 1942
rect 1086 1938 1090 1942
rect 1134 1938 1138 1942
rect 1158 1938 1162 1942
rect 1342 1938 1346 1942
rect 1766 1938 1770 1942
rect 1886 1938 1890 1942
rect 1894 1938 1898 1942
rect 2094 1938 2098 1942
rect 2614 1938 2618 1942
rect 2982 1938 2986 1942
rect 3302 1938 3306 1942
rect 3358 1938 3362 1942
rect 3374 1938 3378 1942
rect 3390 1938 3394 1942
rect 3422 1938 3426 1942
rect 3534 1938 3538 1942
rect 3678 1938 3682 1942
rect 4590 1938 4594 1942
rect 5174 1938 5178 1942
rect 758 1928 762 1932
rect 1646 1928 1650 1932
rect 2422 1928 2426 1932
rect 2710 1928 2714 1932
rect 3350 1928 3354 1932
rect 3526 1928 3530 1932
rect 3790 1928 3794 1932
rect 3838 1928 3842 1932
rect 3982 1928 3986 1932
rect 4014 1928 4018 1932
rect 4390 1928 4394 1932
rect 4614 1928 4618 1932
rect 4878 1928 4882 1932
rect 5062 1928 5066 1932
rect 5150 1928 5154 1932
rect 486 1918 490 1922
rect 814 1918 818 1922
rect 942 1918 946 1922
rect 958 1918 962 1922
rect 1102 1918 1106 1922
rect 1606 1918 1610 1922
rect 1622 1918 1626 1922
rect 1990 1918 1994 1922
rect 2422 1918 2426 1922
rect 2534 1918 2538 1922
rect 2790 1918 2794 1922
rect 3174 1918 3178 1922
rect 4038 1918 4042 1922
rect 4382 1918 4386 1922
rect 4574 1918 4578 1922
rect 558 1908 562 1912
rect 1222 1908 1226 1912
rect 1526 1908 1530 1912
rect 2022 1908 2026 1912
rect 2286 1908 2290 1912
rect 2806 1908 2810 1912
rect 3006 1908 3010 1912
rect 3078 1908 3082 1912
rect 3150 1908 3154 1912
rect 3262 1908 3266 1912
rect 3606 1908 3610 1912
rect 4390 1908 4394 1912
rect 4670 1908 4674 1912
rect 4710 1908 4714 1912
rect 5142 1908 5146 1912
rect 1050 1903 1054 1907
rect 1058 1903 1061 1907
rect 1061 1903 1062 1907
rect 2074 1903 2078 1907
rect 2082 1903 2085 1907
rect 2085 1903 2086 1907
rect 686 1898 690 1902
rect 1214 1898 1218 1902
rect 1734 1898 1738 1902
rect 1894 1898 1898 1902
rect 2318 1898 2322 1902
rect 3098 1903 3102 1907
rect 3106 1903 3109 1907
rect 3109 1903 3110 1907
rect 4114 1903 4118 1907
rect 4122 1903 4125 1907
rect 4125 1903 4126 1907
rect 3086 1898 3090 1902
rect 3134 1898 3138 1902
rect 3262 1898 3266 1902
rect 3486 1898 3490 1902
rect 3494 1898 3498 1902
rect 3822 1898 3826 1902
rect 4094 1898 4098 1902
rect 4462 1898 4466 1902
rect 1734 1888 1738 1892
rect 1966 1888 1970 1892
rect 2006 1888 2010 1892
rect 2350 1888 2354 1892
rect 2374 1888 2378 1892
rect 2430 1888 2434 1892
rect 2446 1888 2450 1892
rect 3078 1888 3082 1892
rect 3366 1888 3370 1892
rect 3414 1888 3418 1892
rect 4342 1888 4346 1892
rect 4438 1888 4442 1892
rect 4822 1888 4826 1892
rect 494 1878 498 1882
rect 574 1868 578 1872
rect 766 1868 770 1872
rect 1158 1878 1162 1882
rect 1374 1878 1378 1882
rect 1582 1878 1586 1882
rect 1590 1878 1594 1882
rect 2094 1878 2098 1882
rect 2918 1878 2922 1882
rect 3030 1878 3034 1882
rect 3798 1878 3802 1882
rect 3822 1878 3826 1882
rect 3902 1878 3906 1882
rect 4238 1878 4242 1882
rect 4326 1878 4330 1882
rect 4406 1878 4410 1882
rect 4854 1878 4858 1882
rect 5014 1878 5018 1882
rect 5142 1878 5146 1882
rect 1174 1868 1178 1872
rect 1230 1868 1234 1872
rect 1470 1868 1474 1872
rect 1806 1868 1810 1872
rect 1846 1868 1850 1872
rect 2086 1868 2090 1872
rect 2134 1868 2138 1872
rect 2566 1868 2570 1872
rect 2806 1868 2810 1872
rect 3182 1868 3186 1872
rect 3254 1868 3258 1872
rect 3582 1868 3586 1872
rect 3894 1868 3898 1872
rect 4062 1868 4066 1872
rect 4174 1868 4178 1872
rect 4286 1868 4290 1872
rect 4478 1868 4482 1872
rect 4710 1868 4714 1872
rect 4718 1868 4722 1872
rect 5118 1868 5122 1872
rect 398 1858 402 1862
rect 470 1858 474 1862
rect 1006 1858 1010 1862
rect 1654 1858 1658 1862
rect 1774 1858 1778 1862
rect 1830 1858 1834 1862
rect 1846 1858 1850 1862
rect 1854 1858 1858 1862
rect 1918 1858 1922 1862
rect 2142 1858 2146 1862
rect 2206 1858 2210 1862
rect 2326 1858 2330 1862
rect 2350 1858 2354 1862
rect 3118 1858 3122 1862
rect 3158 1858 3162 1862
rect 3166 1858 3170 1862
rect 3494 1858 3498 1862
rect 3782 1858 3786 1862
rect 4510 1858 4514 1862
rect 4814 1858 4818 1862
rect 4846 1858 4850 1862
rect 446 1848 450 1852
rect 478 1848 482 1852
rect 694 1848 698 1852
rect 1518 1848 1522 1852
rect 1774 1848 1778 1852
rect 1918 1848 1922 1852
rect 2126 1848 2130 1852
rect 2334 1848 2338 1852
rect 2430 1848 2434 1852
rect 2862 1848 2866 1852
rect 3142 1848 3146 1852
rect 3326 1848 3330 1852
rect 3446 1848 3450 1852
rect 3494 1848 3498 1852
rect 3862 1848 3866 1852
rect 4158 1848 4162 1852
rect 4182 1848 4186 1852
rect 4206 1848 4210 1852
rect 4478 1848 4482 1852
rect 4558 1848 4562 1852
rect 4742 1848 4746 1852
rect 4806 1848 4810 1852
rect 4862 1848 4866 1852
rect 4910 1848 4914 1852
rect 4966 1848 4970 1852
rect 126 1838 130 1842
rect 774 1838 778 1842
rect 1214 1838 1218 1842
rect 2086 1838 2090 1842
rect 2422 1838 2426 1842
rect 3374 1838 3378 1842
rect 3678 1838 3682 1842
rect 4454 1838 4458 1842
rect 1038 1828 1042 1832
rect 1126 1828 1130 1832
rect 1910 1828 1914 1832
rect 2038 1828 2042 1832
rect 2070 1828 2074 1832
rect 3182 1828 3186 1832
rect 3190 1828 3194 1832
rect 4094 1828 4098 1832
rect 4374 1828 4378 1832
rect 4438 1828 4442 1832
rect 446 1818 450 1822
rect 1078 1818 1082 1822
rect 1414 1818 1418 1822
rect 1478 1818 1482 1822
rect 1486 1818 1490 1822
rect 3174 1818 3178 1822
rect 3422 1818 3426 1822
rect 3646 1818 3650 1822
rect 3934 1818 3938 1822
rect 4542 1818 4546 1822
rect 4702 1818 4706 1822
rect 1190 1808 1194 1812
rect 1526 1808 1530 1812
rect 2502 1808 2506 1812
rect 3030 1808 3034 1812
rect 3542 1808 3546 1812
rect 3694 1808 3698 1812
rect 538 1803 542 1807
rect 546 1803 549 1807
rect 549 1803 550 1807
rect 1562 1803 1566 1807
rect 1570 1803 1573 1807
rect 1573 1803 1574 1807
rect 2586 1803 2590 1807
rect 2594 1803 2597 1807
rect 2597 1803 2598 1807
rect 3610 1803 3614 1807
rect 3618 1803 3621 1807
rect 3621 1803 3622 1807
rect 4634 1803 4638 1807
rect 4642 1803 4645 1807
rect 4645 1803 4646 1807
rect 1238 1798 1242 1802
rect 1494 1798 1498 1802
rect 1990 1798 1994 1802
rect 2062 1798 2066 1802
rect 2526 1798 2530 1802
rect 2854 1798 2858 1802
rect 2934 1798 2938 1802
rect 3678 1798 3682 1802
rect 3958 1798 3962 1802
rect 4222 1798 4226 1802
rect 4582 1798 4586 1802
rect 1294 1788 1298 1792
rect 1318 1788 1322 1792
rect 1510 1788 1514 1792
rect 2654 1788 2658 1792
rect 3598 1788 3602 1792
rect 4070 1788 4074 1792
rect 4294 1788 4298 1792
rect 4574 1788 4578 1792
rect 4742 1788 4746 1792
rect 870 1778 874 1782
rect 1190 1778 1194 1782
rect 1254 1778 1258 1782
rect 1294 1778 1298 1782
rect 1366 1778 1370 1782
rect 1542 1778 1546 1782
rect 1710 1778 1714 1782
rect 1870 1778 1874 1782
rect 2078 1778 2082 1782
rect 2430 1778 2434 1782
rect 2622 1778 2626 1782
rect 2638 1778 2642 1782
rect 4374 1778 4378 1782
rect 1350 1768 1354 1772
rect 2782 1768 2786 1772
rect 2990 1768 2994 1772
rect 2998 1768 3002 1772
rect 3054 1768 3058 1772
rect 3758 1768 3762 1772
rect 3982 1768 3986 1772
rect 4062 1768 4066 1772
rect 4918 1768 4922 1772
rect 654 1758 658 1762
rect 3454 1758 3458 1762
rect 3502 1758 3506 1762
rect 3574 1758 3578 1762
rect 3582 1758 3586 1762
rect 4006 1758 4010 1762
rect 4078 1758 4082 1762
rect 4222 1758 4226 1762
rect 4262 1758 4266 1762
rect 4590 1758 4594 1762
rect 5182 1758 5186 1762
rect 702 1748 706 1752
rect 710 1748 714 1752
rect 734 1748 738 1752
rect 1182 1748 1186 1752
rect 1206 1748 1210 1752
rect 1478 1748 1482 1752
rect 382 1738 386 1742
rect 478 1738 482 1742
rect 574 1738 578 1742
rect 1110 1738 1114 1742
rect 1278 1738 1282 1742
rect 1870 1748 1874 1752
rect 1886 1748 1890 1752
rect 2198 1748 2202 1752
rect 2238 1748 2242 1752
rect 2414 1748 2418 1752
rect 2430 1748 2434 1752
rect 2494 1748 2498 1752
rect 2654 1748 2658 1752
rect 2734 1748 2738 1752
rect 2958 1748 2962 1752
rect 2982 1748 2986 1752
rect 2998 1748 3002 1752
rect 3062 1748 3066 1752
rect 3070 1748 3074 1752
rect 3190 1748 3194 1752
rect 3270 1748 3274 1752
rect 3406 1748 3410 1752
rect 3542 1748 3546 1752
rect 3646 1748 3650 1752
rect 3654 1748 3658 1752
rect 3814 1748 3818 1752
rect 3822 1748 3826 1752
rect 4302 1748 4306 1752
rect 4382 1748 4386 1752
rect 4430 1748 4434 1752
rect 4470 1748 4474 1752
rect 4590 1748 4594 1752
rect 1750 1738 1754 1742
rect 2222 1738 2226 1742
rect 2278 1738 2282 1742
rect 2646 1738 2650 1742
rect 2702 1738 2706 1742
rect 2958 1738 2962 1742
rect 3534 1738 3538 1742
rect 4806 1738 4810 1742
rect 5078 1738 5082 1742
rect 1502 1728 1506 1732
rect 1998 1728 2002 1732
rect 2190 1728 2194 1732
rect 3214 1728 3218 1732
rect 3462 1728 3466 1732
rect 3494 1728 3498 1732
rect 4582 1728 4586 1732
rect 4918 1728 4922 1732
rect 910 1718 914 1722
rect 1102 1718 1106 1722
rect 1374 1718 1378 1722
rect 2374 1718 2378 1722
rect 2422 1718 2426 1722
rect 3278 1718 3282 1722
rect 3382 1718 3386 1722
rect 3750 1718 3754 1722
rect 3790 1718 3794 1722
rect 4078 1718 4082 1722
rect 4118 1718 4122 1722
rect 758 1708 762 1712
rect 982 1708 986 1712
rect 1302 1708 1306 1712
rect 1478 1708 1482 1712
rect 1790 1708 1794 1712
rect 1886 1708 1890 1712
rect 2134 1708 2138 1712
rect 2774 1708 2778 1712
rect 2870 1708 2874 1712
rect 3038 1708 3042 1712
rect 3758 1708 3762 1712
rect 3814 1708 3818 1712
rect 4222 1708 4226 1712
rect 4302 1708 4306 1712
rect 1050 1703 1054 1707
rect 1058 1703 1061 1707
rect 1061 1703 1062 1707
rect 2074 1703 2078 1707
rect 2082 1703 2085 1707
rect 2085 1703 2086 1707
rect 3098 1703 3102 1707
rect 3106 1703 3109 1707
rect 3109 1703 3110 1707
rect 4114 1703 4118 1707
rect 4122 1703 4125 1707
rect 4125 1703 4126 1707
rect 670 1698 674 1702
rect 814 1698 818 1702
rect 1030 1698 1034 1702
rect 1326 1698 1330 1702
rect 1662 1698 1666 1702
rect 1798 1698 1802 1702
rect 1862 1698 1866 1702
rect 1966 1698 1970 1702
rect 2846 1698 2850 1702
rect 3230 1698 3234 1702
rect 3454 1698 3458 1702
rect 3510 1698 3514 1702
rect 3766 1698 3770 1702
rect 3966 1698 3970 1702
rect 3990 1698 3994 1702
rect 3998 1698 4002 1702
rect 4782 1698 4786 1702
rect 5022 1698 5026 1702
rect 838 1688 842 1692
rect 950 1688 954 1692
rect 1198 1688 1202 1692
rect 2086 1688 2090 1692
rect 2102 1688 2106 1692
rect 2190 1688 2194 1692
rect 2966 1688 2970 1692
rect 3086 1688 3090 1692
rect 3126 1688 3130 1692
rect 3174 1688 3178 1692
rect 3262 1688 3266 1692
rect 3654 1688 3658 1692
rect 3742 1688 3746 1692
rect 3798 1688 3802 1692
rect 3854 1688 3858 1692
rect 3990 1688 3994 1692
rect 4006 1688 4010 1692
rect 4150 1688 4154 1692
rect 4214 1688 4218 1692
rect 4222 1688 4226 1692
rect 4278 1688 4282 1692
rect 4686 1688 4690 1692
rect 4854 1688 4858 1692
rect 4862 1688 4866 1692
rect 438 1678 442 1682
rect 766 1678 770 1682
rect 1102 1678 1106 1682
rect 1206 1678 1210 1682
rect 1462 1678 1466 1682
rect 1894 1678 1898 1682
rect 1902 1678 1906 1682
rect 2126 1678 2130 1682
rect 2150 1678 2154 1682
rect 2190 1678 2194 1682
rect 2390 1678 2394 1682
rect 2766 1678 2770 1682
rect 3022 1678 3026 1682
rect 3134 1678 3138 1682
rect 3206 1678 3210 1682
rect 3854 1678 3858 1682
rect 4334 1678 4338 1682
rect 4422 1678 4426 1682
rect 4734 1678 4738 1682
rect 358 1668 362 1672
rect 582 1668 586 1672
rect 782 1668 786 1672
rect 1094 1668 1098 1672
rect 1230 1668 1234 1672
rect 1286 1668 1290 1672
rect 1750 1668 1754 1672
rect 1774 1668 1778 1672
rect 2094 1668 2098 1672
rect 2254 1668 2258 1672
rect 2398 1668 2402 1672
rect 2446 1668 2450 1672
rect 2574 1668 2578 1672
rect 2782 1668 2786 1672
rect 3086 1668 3090 1672
rect 3494 1668 3498 1672
rect 3718 1668 3722 1672
rect 3846 1668 3850 1672
rect 4294 1668 4298 1672
rect 4406 1668 4410 1672
rect 4550 1668 4554 1672
rect 4630 1668 4634 1672
rect 4718 1668 4722 1672
rect 4782 1668 4786 1672
rect 5062 1668 5066 1672
rect 646 1658 650 1662
rect 702 1658 706 1662
rect 766 1658 770 1662
rect 910 1658 914 1662
rect 926 1658 930 1662
rect 1246 1658 1250 1662
rect 1366 1658 1370 1662
rect 1486 1658 1490 1662
rect 1814 1658 1818 1662
rect 1886 1658 1890 1662
rect 2950 1658 2954 1662
rect 2966 1658 2970 1662
rect 3374 1658 3378 1662
rect 3382 1658 3386 1662
rect 3838 1658 3842 1662
rect 4366 1658 4370 1662
rect 4438 1658 4442 1662
rect 4446 1658 4450 1662
rect 4470 1658 4474 1662
rect 4574 1658 4578 1662
rect 4670 1658 4674 1662
rect 614 1648 618 1652
rect 1070 1648 1074 1652
rect 1174 1648 1178 1652
rect 1726 1648 1730 1652
rect 1878 1648 1882 1652
rect 2150 1648 2154 1652
rect 2294 1648 2298 1652
rect 2374 1648 2378 1652
rect 2422 1648 2426 1652
rect 2470 1648 2474 1652
rect 3030 1648 3034 1652
rect 3278 1648 3282 1652
rect 3430 1648 3434 1652
rect 3630 1648 3634 1652
rect 3766 1648 3770 1652
rect 4198 1648 4202 1652
rect 4350 1648 4354 1652
rect 4678 1648 4682 1652
rect 5070 1648 5074 1652
rect 358 1638 362 1642
rect 374 1638 378 1642
rect 694 1638 698 1642
rect 950 1638 954 1642
rect 1438 1638 1442 1642
rect 1662 1638 1666 1642
rect 2142 1638 2146 1642
rect 3174 1638 3178 1642
rect 3278 1638 3282 1642
rect 3558 1638 3562 1642
rect 4726 1638 4730 1642
rect 518 1628 522 1632
rect 670 1628 674 1632
rect 702 1628 706 1632
rect 1262 1628 1266 1632
rect 2414 1628 2418 1632
rect 3910 1628 3914 1632
rect 4070 1628 4074 1632
rect 4078 1628 4082 1632
rect 4654 1628 4658 1632
rect 1166 1618 1170 1622
rect 2158 1618 2162 1622
rect 2742 1618 2746 1622
rect 3070 1618 3074 1622
rect 3414 1618 3418 1622
rect 3942 1618 3946 1622
rect 5150 1618 5154 1622
rect 422 1608 426 1612
rect 622 1608 626 1612
rect 1734 1608 1738 1612
rect 3070 1608 3074 1612
rect 3118 1608 3122 1612
rect 4022 1608 4026 1612
rect 4654 1608 4658 1612
rect 538 1603 542 1607
rect 546 1603 549 1607
rect 549 1603 550 1607
rect 1562 1603 1566 1607
rect 1570 1603 1573 1607
rect 1573 1603 1574 1607
rect 2586 1603 2590 1607
rect 2594 1603 2597 1607
rect 2597 1603 2598 1607
rect 3610 1603 3614 1607
rect 3618 1603 3621 1607
rect 3621 1603 3622 1607
rect 4634 1603 4638 1607
rect 4642 1603 4645 1607
rect 4645 1603 4646 1607
rect 734 1598 738 1602
rect 1070 1598 1074 1602
rect 1422 1598 1426 1602
rect 1702 1598 1706 1602
rect 1726 1598 1730 1602
rect 1974 1598 1978 1602
rect 2342 1598 2346 1602
rect 2998 1598 3002 1602
rect 3006 1598 3010 1602
rect 3630 1598 3634 1602
rect 4374 1598 4378 1602
rect 4606 1598 4610 1602
rect 1014 1588 1018 1592
rect 1046 1588 1050 1592
rect 1318 1588 1322 1592
rect 1774 1588 1778 1592
rect 2030 1588 2034 1592
rect 2982 1588 2986 1592
rect 3118 1588 3122 1592
rect 4006 1588 4010 1592
rect 4030 1588 4034 1592
rect 4038 1588 4042 1592
rect 4102 1588 4106 1592
rect 4342 1588 4346 1592
rect 4806 1588 4810 1592
rect 734 1578 738 1582
rect 1078 1578 1082 1582
rect 1198 1578 1202 1582
rect 1542 1578 1546 1582
rect 1910 1578 1914 1582
rect 1926 1578 1930 1582
rect 2206 1578 2210 1582
rect 2230 1578 2234 1582
rect 2238 1578 2242 1582
rect 2302 1578 2306 1582
rect 2310 1578 2314 1582
rect 2910 1578 2914 1582
rect 3350 1578 3354 1582
rect 3414 1578 3418 1582
rect 3750 1578 3754 1582
rect 734 1568 738 1572
rect 942 1568 946 1572
rect 1014 1568 1018 1572
rect 1046 1568 1050 1572
rect 3166 1568 3170 1572
rect 3174 1568 3178 1572
rect 4390 1568 4394 1572
rect 4798 1568 4802 1572
rect 5046 1568 5050 1572
rect 462 1558 466 1562
rect 614 1558 618 1562
rect 998 1558 1002 1562
rect 1142 1558 1146 1562
rect 1318 1558 1322 1562
rect 1566 1558 1570 1562
rect 1598 1558 1602 1562
rect 1782 1558 1786 1562
rect 1926 1558 1930 1562
rect 2102 1558 2106 1562
rect 2190 1558 2194 1562
rect 2518 1558 2522 1562
rect 2886 1558 2890 1562
rect 3030 1558 3034 1562
rect 3142 1558 3146 1562
rect 3622 1558 3626 1562
rect 3958 1558 3962 1562
rect 358 1548 362 1552
rect 606 1548 610 1552
rect 774 1548 778 1552
rect 990 1548 994 1552
rect 1022 1548 1026 1552
rect 1030 1548 1034 1552
rect 1086 1548 1090 1552
rect 1150 1548 1154 1552
rect 1158 1548 1162 1552
rect 1214 1548 1218 1552
rect 1390 1548 1394 1552
rect 1414 1548 1418 1552
rect 1494 1548 1498 1552
rect 1558 1548 1562 1552
rect 1566 1548 1570 1552
rect 1590 1548 1594 1552
rect 1702 1548 1706 1552
rect 1734 1548 1738 1552
rect 1838 1548 1842 1552
rect 1950 1548 1954 1552
rect 1982 1548 1986 1552
rect 2054 1548 2058 1552
rect 2198 1548 2202 1552
rect 2206 1548 2210 1552
rect 2238 1548 2242 1552
rect 2286 1548 2290 1552
rect 2310 1548 2314 1552
rect 2734 1548 2738 1552
rect 2846 1548 2850 1552
rect 2862 1548 2866 1552
rect 2878 1548 2882 1552
rect 2910 1548 2914 1552
rect 3054 1548 3058 1552
rect 3246 1548 3250 1552
rect 3542 1548 3546 1552
rect 3814 1548 3818 1552
rect 3846 1548 3850 1552
rect 4054 1558 4058 1562
rect 4830 1558 4834 1562
rect 5046 1558 5050 1562
rect 5166 1558 5170 1562
rect 3966 1548 3970 1552
rect 3990 1548 3994 1552
rect 4078 1548 4082 1552
rect 222 1538 226 1542
rect 406 1538 410 1542
rect 526 1538 530 1542
rect 790 1538 794 1542
rect 950 1538 954 1542
rect 1470 1538 1474 1542
rect 1766 1538 1770 1542
rect 2238 1538 2242 1542
rect 2390 1538 2394 1542
rect 2998 1538 3002 1542
rect 3006 1538 3010 1542
rect 3022 1538 3026 1542
rect 3062 1538 3066 1542
rect 3342 1538 3346 1542
rect 3350 1538 3354 1542
rect 3718 1538 3722 1542
rect 3902 1538 3906 1542
rect 5014 1538 5018 1542
rect 326 1528 330 1532
rect 670 1528 674 1532
rect 1126 1528 1130 1532
rect 1198 1528 1202 1532
rect 1502 1528 1506 1532
rect 1518 1528 1522 1532
rect 1534 1528 1538 1532
rect 1566 1528 1570 1532
rect 1710 1528 1714 1532
rect 1958 1528 1962 1532
rect 2094 1528 2098 1532
rect 2222 1528 2226 1532
rect 2286 1528 2290 1532
rect 2750 1528 2754 1532
rect 2854 1528 2858 1532
rect 2894 1528 2898 1532
rect 2942 1528 2946 1532
rect 2958 1528 2962 1532
rect 3214 1528 3218 1532
rect 3238 1528 3242 1532
rect 3534 1528 3538 1532
rect 3686 1528 3690 1532
rect 3894 1528 3898 1532
rect 4158 1528 4162 1532
rect 4854 1528 4858 1532
rect 5038 1528 5042 1532
rect 5102 1528 5106 1532
rect 286 1518 290 1522
rect 718 1518 722 1522
rect 1022 1518 1026 1522
rect 1318 1518 1322 1522
rect 1782 1518 1786 1522
rect 1918 1518 1922 1522
rect 2694 1518 2698 1522
rect 2814 1518 2818 1522
rect 2846 1518 2850 1522
rect 3646 1518 3650 1522
rect 3862 1518 3866 1522
rect 4150 1518 4154 1522
rect 654 1508 658 1512
rect 1166 1508 1170 1512
rect 1342 1508 1346 1512
rect 2094 1508 2098 1512
rect 2262 1508 2266 1512
rect 4102 1508 4106 1512
rect 4166 1508 4170 1512
rect 1050 1503 1054 1507
rect 1058 1503 1061 1507
rect 1061 1503 1062 1507
rect 2074 1503 2078 1507
rect 2082 1503 2085 1507
rect 2085 1503 2086 1507
rect 3098 1503 3102 1507
rect 3106 1503 3109 1507
rect 3109 1503 3110 1507
rect 4114 1503 4118 1507
rect 4122 1503 4125 1507
rect 4125 1503 4126 1507
rect 942 1498 946 1502
rect 1390 1498 1394 1502
rect 2126 1498 2130 1502
rect 2150 1498 2154 1502
rect 2342 1498 2346 1502
rect 2462 1498 2466 1502
rect 2790 1498 2794 1502
rect 2982 1498 2986 1502
rect 3134 1498 3138 1502
rect 3574 1498 3578 1502
rect 4158 1498 4162 1502
rect 4870 1498 4874 1502
rect 5086 1498 5090 1502
rect 670 1488 674 1492
rect 934 1488 938 1492
rect 1302 1488 1306 1492
rect 1422 1488 1426 1492
rect 1486 1488 1490 1492
rect 1510 1488 1514 1492
rect 1550 1488 1554 1492
rect 1678 1488 1682 1492
rect 2438 1488 2442 1492
rect 2750 1488 2754 1492
rect 2782 1488 2786 1492
rect 2798 1488 2802 1492
rect 3142 1488 3146 1492
rect 3318 1488 3322 1492
rect 3590 1488 3594 1492
rect 3686 1488 3690 1492
rect 3734 1488 3738 1492
rect 3918 1488 3922 1492
rect 3926 1488 3930 1492
rect 4126 1488 4130 1492
rect 4942 1488 4946 1492
rect 1598 1478 1602 1482
rect 2182 1478 2186 1482
rect 2198 1478 2202 1482
rect 2326 1478 2330 1482
rect 3854 1478 3858 1482
rect 3974 1478 3978 1482
rect 4742 1478 4746 1482
rect 4766 1478 4770 1482
rect 4934 1478 4938 1482
rect 414 1468 418 1472
rect 430 1468 434 1472
rect 630 1468 634 1472
rect 662 1468 666 1472
rect 742 1468 746 1472
rect 758 1468 762 1472
rect 766 1468 770 1472
rect 926 1468 930 1472
rect 318 1458 322 1462
rect 446 1458 450 1462
rect 558 1458 562 1462
rect 958 1468 962 1472
rect 1038 1468 1042 1472
rect 1646 1468 1650 1472
rect 1678 1468 1682 1472
rect 1798 1468 1802 1472
rect 1942 1468 1946 1472
rect 2086 1468 2090 1472
rect 2166 1468 2170 1472
rect 2614 1468 2618 1472
rect 2686 1468 2690 1472
rect 3038 1468 3042 1472
rect 3054 1468 3058 1472
rect 3190 1468 3194 1472
rect 3438 1468 3442 1472
rect 3462 1468 3466 1472
rect 4246 1468 4250 1472
rect 4318 1468 4322 1472
rect 4358 1468 4362 1472
rect 4854 1468 4858 1472
rect 4910 1468 4914 1472
rect 1134 1458 1138 1462
rect 1198 1458 1202 1462
rect 1326 1458 1330 1462
rect 1350 1458 1354 1462
rect 1774 1458 1778 1462
rect 1974 1458 1978 1462
rect 2038 1458 2042 1462
rect 2462 1458 2466 1462
rect 2934 1458 2938 1462
rect 3206 1458 3210 1462
rect 3566 1458 3570 1462
rect 3630 1458 3634 1462
rect 3902 1458 3906 1462
rect 3990 1458 3994 1462
rect 438 1448 442 1452
rect 638 1448 642 1452
rect 1030 1448 1034 1452
rect 1526 1448 1530 1452
rect 1758 1448 1762 1452
rect 2198 1448 2202 1452
rect 2254 1448 2258 1452
rect 2686 1448 2690 1452
rect 3350 1448 3354 1452
rect 3870 1448 3874 1452
rect 4254 1448 4258 1452
rect 5110 1448 5114 1452
rect 798 1438 802 1442
rect 2094 1438 2098 1442
rect 2102 1438 2106 1442
rect 2190 1438 2194 1442
rect 2422 1438 2426 1442
rect 2798 1438 2802 1442
rect 3014 1438 3018 1442
rect 3918 1438 3922 1442
rect 3934 1438 3938 1442
rect 4710 1438 4714 1442
rect 374 1428 378 1432
rect 438 1428 442 1432
rect 782 1428 786 1432
rect 990 1428 994 1432
rect 1198 1428 1202 1432
rect 1222 1428 1226 1432
rect 1366 1428 1370 1432
rect 1550 1428 1554 1432
rect 1742 1428 1746 1432
rect 1750 1428 1754 1432
rect 2134 1428 2138 1432
rect 2182 1428 2186 1432
rect 2918 1428 2922 1432
rect 4046 1428 4050 1432
rect 4750 1428 4754 1432
rect 374 1418 378 1422
rect 1110 1418 1114 1422
rect 2046 1418 2050 1422
rect 2086 1418 2090 1422
rect 2166 1418 2170 1422
rect 2422 1418 2426 1422
rect 3070 1418 3074 1422
rect 3126 1418 3130 1422
rect 3158 1418 3162 1422
rect 3254 1418 3258 1422
rect 3406 1418 3410 1422
rect 4142 1418 4146 1422
rect 4446 1418 4450 1422
rect 662 1408 666 1412
rect 742 1408 746 1412
rect 1422 1408 1426 1412
rect 1638 1408 1642 1412
rect 2054 1408 2058 1412
rect 2086 1408 2090 1412
rect 2742 1408 2746 1412
rect 3422 1408 3426 1412
rect 3950 1408 3954 1412
rect 4014 1408 4018 1412
rect 4246 1408 4250 1412
rect 4694 1408 4698 1412
rect 4782 1408 4786 1412
rect 4854 1408 4858 1412
rect 538 1403 542 1407
rect 546 1403 549 1407
rect 549 1403 550 1407
rect 1562 1403 1566 1407
rect 1570 1403 1573 1407
rect 1573 1403 1574 1407
rect 2586 1403 2590 1407
rect 2594 1403 2597 1407
rect 2597 1403 2598 1407
rect 3610 1403 3614 1407
rect 3618 1403 3621 1407
rect 3621 1403 3622 1407
rect 4634 1403 4638 1407
rect 4642 1403 4645 1407
rect 4645 1403 4646 1407
rect 126 1398 130 1402
rect 526 1398 530 1402
rect 686 1398 690 1402
rect 806 1398 810 1402
rect 1238 1398 1242 1402
rect 1742 1398 1746 1402
rect 2118 1398 2122 1402
rect 2246 1398 2250 1402
rect 2574 1398 2578 1402
rect 3966 1398 3970 1402
rect 414 1388 418 1392
rect 654 1388 658 1392
rect 998 1388 1002 1392
rect 1214 1388 1218 1392
rect 2150 1388 2154 1392
rect 2302 1388 2306 1392
rect 2558 1388 2562 1392
rect 2838 1388 2842 1392
rect 3022 1388 3026 1392
rect 3286 1388 3290 1392
rect 3454 1388 3458 1392
rect 4134 1388 4138 1392
rect 502 1378 506 1382
rect 526 1378 530 1382
rect 1638 1378 1642 1382
rect 1902 1378 1906 1382
rect 2478 1378 2482 1382
rect 2574 1378 2578 1382
rect 2918 1378 2922 1382
rect 3390 1378 3394 1382
rect 4862 1378 4866 1382
rect 4926 1378 4930 1382
rect 638 1368 642 1372
rect 1390 1368 1394 1372
rect 1710 1368 1714 1372
rect 2550 1368 2554 1372
rect 2678 1368 2682 1372
rect 2886 1368 2890 1372
rect 3382 1368 3386 1372
rect 3630 1368 3634 1372
rect 3814 1368 3818 1372
rect 4230 1368 4234 1372
rect 4846 1368 4850 1372
rect 838 1358 842 1362
rect 846 1358 850 1362
rect 942 1358 946 1362
rect 1094 1358 1098 1362
rect 1102 1358 1106 1362
rect 1350 1358 1354 1362
rect 1374 1358 1378 1362
rect 1406 1358 1410 1362
rect 1502 1358 1506 1362
rect 1606 1358 1610 1362
rect 1646 1358 1650 1362
rect 2310 1358 2314 1362
rect 2326 1358 2330 1362
rect 2630 1358 2634 1362
rect 2646 1358 2650 1362
rect 2654 1358 2658 1362
rect 3294 1358 3298 1362
rect 3534 1358 3538 1362
rect 3654 1358 3658 1362
rect 3766 1358 3770 1362
rect 4054 1358 4058 1362
rect 4982 1358 4986 1362
rect 5054 1358 5058 1362
rect 414 1348 418 1352
rect 566 1348 570 1352
rect 598 1348 602 1352
rect 854 1348 858 1352
rect 886 1348 890 1352
rect 918 1348 922 1352
rect 942 1348 946 1352
rect 974 1348 978 1352
rect 1222 1348 1226 1352
rect 1390 1348 1394 1352
rect 1542 1348 1546 1352
rect 1766 1348 1770 1352
rect 2006 1348 2010 1352
rect 2062 1348 2066 1352
rect 2110 1348 2114 1352
rect 2382 1348 2386 1352
rect 2390 1348 2394 1352
rect 2486 1348 2490 1352
rect 2758 1348 2762 1352
rect 2822 1348 2826 1352
rect 3006 1348 3010 1352
rect 3166 1348 3170 1352
rect 3662 1348 3666 1352
rect 3670 1348 3674 1352
rect 3830 1348 3834 1352
rect 4014 1348 4018 1352
rect 4046 1348 4050 1352
rect 4078 1348 4082 1352
rect 4190 1348 4194 1352
rect 4982 1348 4986 1352
rect 342 1338 346 1342
rect 558 1338 562 1342
rect 678 1338 682 1342
rect 878 1338 882 1342
rect 1198 1338 1202 1342
rect 1334 1338 1338 1342
rect 1366 1338 1370 1342
rect 1494 1338 1498 1342
rect 1558 1338 1562 1342
rect 1614 1338 1618 1342
rect 2094 1338 2098 1342
rect 2534 1338 2538 1342
rect 2574 1338 2578 1342
rect 2742 1338 2746 1342
rect 3214 1338 3218 1342
rect 3318 1338 3322 1342
rect 3894 1338 3898 1342
rect 4286 1338 4290 1342
rect 4390 1338 4394 1342
rect 422 1328 426 1332
rect 462 1328 466 1332
rect 806 1328 810 1332
rect 862 1328 866 1332
rect 1254 1328 1258 1332
rect 2158 1328 2162 1332
rect 2270 1328 2274 1332
rect 2550 1328 2554 1332
rect 2870 1328 2874 1332
rect 2934 1328 2938 1332
rect 3110 1328 3114 1332
rect 3134 1328 3138 1332
rect 3246 1328 3250 1332
rect 3614 1328 3618 1332
rect 3878 1328 3882 1332
rect 4886 1328 4890 1332
rect 278 1318 282 1322
rect 590 1318 594 1322
rect 830 1318 834 1322
rect 1166 1318 1170 1322
rect 1542 1318 1546 1322
rect 1590 1318 1594 1322
rect 2862 1318 2866 1322
rect 2870 1318 2874 1322
rect 3022 1318 3026 1322
rect 3246 1318 3250 1322
rect 3294 1318 3298 1322
rect 3710 1318 3714 1322
rect 4070 1318 4074 1322
rect 4302 1318 4306 1322
rect 4334 1318 4338 1322
rect 1222 1308 1226 1312
rect 1238 1308 1242 1312
rect 1334 1308 1338 1312
rect 1742 1308 1746 1312
rect 2398 1308 2402 1312
rect 3222 1308 3226 1312
rect 3230 1308 3234 1312
rect 4022 1308 4026 1312
rect 4422 1308 4426 1312
rect 1050 1303 1054 1307
rect 1058 1303 1061 1307
rect 1061 1303 1062 1307
rect 2074 1303 2078 1307
rect 2082 1303 2085 1307
rect 2085 1303 2086 1307
rect 3098 1303 3102 1307
rect 3106 1303 3109 1307
rect 3109 1303 3110 1307
rect 4114 1303 4118 1307
rect 4122 1303 4125 1307
rect 4125 1303 4126 1307
rect 1038 1298 1042 1302
rect 1550 1298 1554 1302
rect 2422 1298 2426 1302
rect 2518 1298 2522 1302
rect 2854 1298 2858 1302
rect 3446 1298 3450 1302
rect 4310 1298 4314 1302
rect 4678 1298 4682 1302
rect 4782 1298 4786 1302
rect 334 1288 338 1292
rect 750 1288 754 1292
rect 1222 1288 1226 1292
rect 1598 1288 1602 1292
rect 1710 1288 1714 1292
rect 1942 1288 1946 1292
rect 2206 1288 2210 1292
rect 2982 1288 2986 1292
rect 3150 1288 3154 1292
rect 3246 1288 3250 1292
rect 3358 1288 3362 1292
rect 3438 1288 3442 1292
rect 3454 1288 3458 1292
rect 4702 1288 4706 1292
rect 302 1278 306 1282
rect 358 1278 362 1282
rect 710 1278 714 1282
rect 1454 1278 1458 1282
rect 1582 1278 1586 1282
rect 1942 1278 1946 1282
rect 2742 1278 2746 1282
rect 3166 1278 3170 1282
rect 3182 1278 3186 1282
rect 3398 1278 3402 1282
rect 3414 1278 3418 1282
rect 3830 1278 3834 1282
rect 3902 1278 3906 1282
rect 4598 1278 4602 1282
rect 4766 1278 4770 1282
rect 4774 1278 4778 1282
rect 102 1268 106 1272
rect 222 1268 226 1272
rect 446 1268 450 1272
rect 470 1268 474 1272
rect 590 1268 594 1272
rect 670 1268 674 1272
rect 1006 1268 1010 1272
rect 1086 1268 1090 1272
rect 1198 1268 1202 1272
rect 1326 1268 1330 1272
rect 1382 1268 1386 1272
rect 1398 1268 1402 1272
rect 1950 1268 1954 1272
rect 1982 1268 1986 1272
rect 2022 1268 2026 1272
rect 2078 1268 2082 1272
rect 2294 1268 2298 1272
rect 2958 1268 2962 1272
rect 3158 1268 3162 1272
rect 3214 1268 3218 1272
rect 3222 1268 3226 1272
rect 3678 1268 3682 1272
rect 3734 1268 3738 1272
rect 3814 1268 3818 1272
rect 4582 1268 4586 1272
rect 4662 1268 4666 1272
rect 5054 1268 5058 1272
rect 358 1258 362 1262
rect 390 1258 394 1262
rect 710 1258 714 1262
rect 846 1258 850 1262
rect 982 1258 986 1262
rect 1006 1258 1010 1262
rect 1110 1258 1114 1262
rect 1126 1258 1130 1262
rect 1214 1258 1218 1262
rect 1358 1258 1362 1262
rect 1406 1258 1410 1262
rect 1606 1258 1610 1262
rect 1638 1258 1642 1262
rect 1662 1258 1666 1262
rect 2086 1258 2090 1262
rect 2166 1258 2170 1262
rect 2422 1258 2426 1262
rect 2646 1258 2650 1262
rect 2806 1258 2810 1262
rect 3038 1258 3042 1262
rect 3254 1258 3258 1262
rect 3558 1258 3562 1262
rect 3622 1258 3626 1262
rect 4046 1258 4050 1262
rect 4238 1258 4242 1262
rect 4350 1258 4354 1262
rect 4366 1258 4370 1262
rect 4374 1258 4378 1262
rect 4574 1258 4578 1262
rect 4678 1258 4682 1262
rect 4774 1258 4778 1262
rect 5030 1258 5034 1262
rect 238 1248 242 1252
rect 1198 1248 1202 1252
rect 2142 1248 2146 1252
rect 2206 1248 2210 1252
rect 2414 1248 2418 1252
rect 2582 1248 2586 1252
rect 3150 1248 3154 1252
rect 3190 1248 3194 1252
rect 3454 1248 3458 1252
rect 1262 1238 1266 1242
rect 1406 1238 1410 1242
rect 3158 1238 3162 1242
rect 3718 1248 3722 1252
rect 3790 1248 3794 1252
rect 3830 1248 3834 1252
rect 3838 1248 3842 1252
rect 4254 1248 4258 1252
rect 4718 1248 4722 1252
rect 5014 1248 5018 1252
rect 3526 1238 3530 1242
rect 3630 1238 3634 1242
rect 3790 1238 3794 1242
rect 3878 1238 3882 1242
rect 3886 1238 3890 1242
rect 4350 1238 4354 1242
rect 4438 1238 4442 1242
rect 4750 1238 4754 1242
rect 4806 1238 4810 1242
rect 830 1228 834 1232
rect 1766 1228 1770 1232
rect 2214 1228 2218 1232
rect 3158 1228 3162 1232
rect 3702 1228 3706 1232
rect 3750 1228 3754 1232
rect 4710 1228 4714 1232
rect 5054 1228 5058 1232
rect 166 1218 170 1222
rect 454 1218 458 1222
rect 1310 1218 1314 1222
rect 1734 1218 1738 1222
rect 1974 1218 1978 1222
rect 2102 1218 2106 1222
rect 2710 1218 2714 1222
rect 4086 1218 4090 1222
rect 374 1208 378 1212
rect 398 1208 402 1212
rect 630 1208 634 1212
rect 686 1208 690 1212
rect 1294 1208 1298 1212
rect 2038 1208 2042 1212
rect 2102 1208 2106 1212
rect 2262 1208 2266 1212
rect 2542 1208 2546 1212
rect 2622 1208 2626 1212
rect 3150 1208 3154 1212
rect 3302 1208 3306 1212
rect 3462 1208 3466 1212
rect 3966 1208 3970 1212
rect 3998 1208 4002 1212
rect 4462 1208 4466 1212
rect 538 1203 542 1207
rect 546 1203 549 1207
rect 549 1203 550 1207
rect 1562 1203 1566 1207
rect 1570 1203 1573 1207
rect 1573 1203 1574 1207
rect 2586 1203 2590 1207
rect 2594 1203 2597 1207
rect 2597 1203 2598 1207
rect 902 1198 906 1202
rect 1182 1198 1186 1202
rect 3610 1203 3614 1207
rect 3618 1203 3621 1207
rect 3621 1203 3622 1207
rect 4634 1203 4638 1207
rect 4642 1203 4645 1207
rect 4645 1203 4646 1207
rect 3358 1198 3362 1202
rect 3454 1198 3458 1202
rect 3950 1198 3954 1202
rect 2614 1188 2618 1192
rect 2622 1188 2626 1192
rect 3214 1188 3218 1192
rect 3278 1188 3282 1192
rect 3310 1188 3314 1192
rect 4254 1188 4258 1192
rect 4518 1188 4522 1192
rect 2014 1178 2018 1182
rect 3022 1178 3026 1182
rect 3998 1178 4002 1182
rect 4070 1178 4074 1182
rect 926 1168 930 1172
rect 1526 1168 1530 1172
rect 2294 1168 2298 1172
rect 2630 1168 2634 1172
rect 2998 1168 3002 1172
rect 3286 1168 3290 1172
rect 3854 1168 3858 1172
rect 3870 1168 3874 1172
rect 3910 1168 3914 1172
rect 4158 1168 4162 1172
rect 222 1158 226 1162
rect 1174 1158 1178 1162
rect 1414 1158 1418 1162
rect 1446 1158 1450 1162
rect 1518 1158 1522 1162
rect 2014 1158 2018 1162
rect 2046 1158 2050 1162
rect 2678 1158 2682 1162
rect 2766 1158 2770 1162
rect 3230 1158 3234 1162
rect 3638 1158 3642 1162
rect 3798 1158 3802 1162
rect 3830 1158 3834 1162
rect 4054 1158 4058 1162
rect 4174 1158 4178 1162
rect 4342 1158 4346 1162
rect 4358 1158 4362 1162
rect 4478 1158 4482 1162
rect 4502 1158 4506 1162
rect 4526 1158 4530 1162
rect 4566 1158 4570 1162
rect 134 1148 138 1152
rect 470 1148 474 1152
rect 558 1148 562 1152
rect 582 1148 586 1152
rect 782 1148 786 1152
rect 830 1148 834 1152
rect 894 1148 898 1152
rect 958 1148 962 1152
rect 1022 1148 1026 1152
rect 1046 1148 1050 1152
rect 1238 1148 1242 1152
rect 1342 1148 1346 1152
rect 1494 1148 1498 1152
rect 1558 1148 1562 1152
rect 1710 1148 1714 1152
rect 2254 1148 2258 1152
rect 2526 1148 2530 1152
rect 2710 1148 2714 1152
rect 2926 1148 2930 1152
rect 3110 1148 3114 1152
rect 3318 1148 3322 1152
rect 3342 1148 3346 1152
rect 3382 1148 3386 1152
rect 3518 1148 3522 1152
rect 3526 1148 3530 1152
rect 3678 1148 3682 1152
rect 3806 1148 3810 1152
rect 3902 1148 3906 1152
rect 4102 1148 4106 1152
rect 4390 1148 4394 1152
rect 4542 1148 4546 1152
rect 4638 1148 4642 1152
rect 4694 1148 4698 1152
rect 734 1138 738 1142
rect 822 1138 826 1142
rect 998 1138 1002 1142
rect 1078 1138 1082 1142
rect 1174 1138 1178 1142
rect 1614 1138 1618 1142
rect 1678 1138 1682 1142
rect 1718 1138 1722 1142
rect 2014 1138 2018 1142
rect 2046 1138 2050 1142
rect 2062 1138 2066 1142
rect 2198 1138 2202 1142
rect 2702 1138 2706 1142
rect 3126 1138 3130 1142
rect 3294 1138 3298 1142
rect 4382 1138 4386 1142
rect 4422 1138 4426 1142
rect 4486 1138 4490 1142
rect 4662 1138 4666 1142
rect 4862 1138 4866 1142
rect 246 1128 250 1132
rect 462 1128 466 1132
rect 614 1128 618 1132
rect 654 1128 658 1132
rect 742 1128 746 1132
rect 766 1128 770 1132
rect 2190 1128 2194 1132
rect 2606 1128 2610 1132
rect 3494 1128 3498 1132
rect 3886 1128 3890 1132
rect 3942 1128 3946 1132
rect 4110 1128 4114 1132
rect 358 1118 362 1122
rect 902 1118 906 1122
rect 1702 1118 1706 1122
rect 3518 1118 3522 1122
rect 3558 1118 3562 1122
rect 3678 1118 3682 1122
rect 3742 1118 3746 1122
rect 4054 1118 4058 1122
rect 4526 1118 4530 1122
rect 4926 1118 4930 1122
rect 398 1108 402 1112
rect 798 1108 802 1112
rect 870 1108 874 1112
rect 1150 1108 1154 1112
rect 1758 1108 1762 1112
rect 1806 1108 1810 1112
rect 1990 1108 1994 1112
rect 2654 1108 2658 1112
rect 1050 1103 1054 1107
rect 1058 1103 1061 1107
rect 1061 1103 1062 1107
rect 2074 1103 2078 1107
rect 2082 1103 2085 1107
rect 2085 1103 2086 1107
rect 3098 1103 3102 1107
rect 3106 1103 3109 1107
rect 3109 1103 3110 1107
rect 4114 1103 4118 1107
rect 4122 1103 4125 1107
rect 4125 1103 4126 1107
rect 990 1098 994 1102
rect 1174 1098 1178 1102
rect 1654 1098 1658 1102
rect 2110 1098 2114 1102
rect 2182 1098 2186 1102
rect 2246 1098 2250 1102
rect 2574 1098 2578 1102
rect 2734 1098 2738 1102
rect 3174 1098 3178 1102
rect 3598 1098 3602 1102
rect 3694 1098 3698 1102
rect 478 1088 482 1092
rect 742 1088 746 1092
rect 1398 1088 1402 1092
rect 1878 1088 1882 1092
rect 2734 1088 2738 1092
rect 3206 1088 3210 1092
rect 3662 1088 3666 1092
rect 862 1078 866 1082
rect 1078 1078 1082 1082
rect 1494 1078 1498 1082
rect 1966 1078 1970 1082
rect 2230 1078 2234 1082
rect 3006 1078 3010 1082
rect 3070 1078 3074 1082
rect 3134 1078 3138 1082
rect 3182 1078 3186 1082
rect 3654 1078 3658 1082
rect 3766 1078 3770 1082
rect 4030 1078 4034 1082
rect 222 1068 226 1072
rect 710 1068 714 1072
rect 862 1068 866 1072
rect 894 1068 898 1072
rect 1070 1068 1074 1072
rect 1094 1068 1098 1072
rect 1102 1068 1106 1072
rect 1446 1068 1450 1072
rect 1710 1068 1714 1072
rect 1774 1068 1778 1072
rect 1846 1068 1850 1072
rect 1878 1068 1882 1072
rect 1902 1068 1906 1072
rect 1910 1068 1914 1072
rect 2150 1068 2154 1072
rect 2238 1068 2242 1072
rect 2678 1068 2682 1072
rect 2726 1068 2730 1072
rect 2758 1068 2762 1072
rect 3078 1068 3082 1072
rect 3334 1068 3338 1072
rect 3342 1068 3346 1072
rect 3462 1068 3466 1072
rect 3486 1068 3490 1072
rect 3502 1068 3506 1072
rect 3934 1068 3938 1072
rect 4094 1068 4098 1072
rect 4550 1068 4554 1072
rect 422 1058 426 1062
rect 926 1058 930 1062
rect 958 1058 962 1062
rect 1054 1058 1058 1062
rect 1614 1058 1618 1062
rect 1654 1058 1658 1062
rect 2014 1058 2018 1062
rect 2206 1058 2210 1062
rect 2270 1058 2274 1062
rect 2510 1058 2514 1062
rect 2590 1058 2594 1062
rect 2630 1058 2634 1062
rect 2694 1058 2698 1062
rect 2726 1058 2730 1062
rect 3310 1058 3314 1062
rect 3742 1058 3746 1062
rect 3758 1058 3762 1062
rect 3870 1058 3874 1062
rect 4526 1058 4530 1062
rect 4710 1058 4714 1062
rect 4758 1058 4762 1062
rect 4814 1058 4818 1062
rect 1302 1048 1306 1052
rect 1558 1048 1562 1052
rect 414 1038 418 1042
rect 558 1038 562 1042
rect 894 1038 898 1042
rect 1134 1038 1138 1042
rect 2158 1048 2162 1052
rect 2966 1048 2970 1052
rect 3182 1048 3186 1052
rect 3446 1048 3450 1052
rect 3462 1048 3466 1052
rect 3766 1048 3770 1052
rect 3782 1048 3786 1052
rect 4054 1048 4058 1052
rect 4190 1048 4194 1052
rect 1286 1038 1290 1042
rect 2222 1038 2226 1042
rect 3366 1038 3370 1042
rect 3382 1038 3386 1042
rect 3558 1038 3562 1042
rect 3750 1038 3754 1042
rect 910 1028 914 1032
rect 1598 1028 1602 1032
rect 2134 1028 2138 1032
rect 2142 1028 2146 1032
rect 2430 1028 2434 1032
rect 3782 1028 3786 1032
rect 1102 1018 1106 1022
rect 1246 1018 1250 1022
rect 2014 1018 2018 1022
rect 2830 1018 2834 1022
rect 3030 1018 3034 1022
rect 3814 1018 3818 1022
rect 4742 1018 4746 1022
rect 494 1008 498 1012
rect 2006 1008 2010 1012
rect 2614 1008 2618 1012
rect 3078 1008 3082 1012
rect 3510 1008 3514 1012
rect 3766 1008 3770 1012
rect 4198 1008 4202 1012
rect 4678 1008 4682 1012
rect 538 1003 542 1007
rect 546 1003 549 1007
rect 549 1003 550 1007
rect 1562 1003 1566 1007
rect 1570 1003 1573 1007
rect 1573 1003 1574 1007
rect 2586 1003 2590 1007
rect 2594 1003 2597 1007
rect 2597 1003 2598 1007
rect 3610 1003 3614 1007
rect 3618 1003 3621 1007
rect 3621 1003 3622 1007
rect 4634 1003 4638 1007
rect 4642 1003 4645 1007
rect 4645 1003 4646 1007
rect 2574 998 2578 1002
rect 2902 998 2906 1002
rect 3238 998 3242 1002
rect 4142 998 4146 1002
rect 4694 998 4698 1002
rect 238 988 242 992
rect 462 988 466 992
rect 1422 988 1426 992
rect 1806 988 1810 992
rect 1830 988 1834 992
rect 2118 988 2122 992
rect 2678 988 2682 992
rect 3062 988 3066 992
rect 3990 988 3994 992
rect 4574 988 4578 992
rect 662 978 666 982
rect 1134 978 1138 982
rect 1318 978 1322 982
rect 1606 978 1610 982
rect 2054 978 2058 982
rect 2814 978 2818 982
rect 3118 978 3122 982
rect 3270 978 3274 982
rect 5062 978 5066 982
rect 102 968 106 972
rect 406 968 410 972
rect 830 968 834 972
rect 1182 968 1186 972
rect 1662 968 1666 972
rect 1830 968 1834 972
rect 2094 968 2098 972
rect 2542 968 2546 972
rect 3470 968 3474 972
rect 3942 968 3946 972
rect 4414 968 4418 972
rect 342 958 346 962
rect 1462 958 1466 962
rect 1550 958 1554 962
rect 2558 958 2562 962
rect 2758 958 2762 962
rect 3126 958 3130 962
rect 3142 958 3146 962
rect 3422 958 3426 962
rect 3918 958 3922 962
rect 3990 958 3994 962
rect 4390 958 4394 962
rect 4886 958 4890 962
rect 366 948 370 952
rect 654 948 658 952
rect 1390 948 1394 952
rect 1478 948 1482 952
rect 1502 948 1506 952
rect 1662 948 1666 952
rect 1774 948 1778 952
rect 2086 948 2090 952
rect 2222 948 2226 952
rect 2486 948 2490 952
rect 606 938 610 942
rect 702 938 706 942
rect 726 938 730 942
rect 814 938 818 942
rect 998 938 1002 942
rect 1174 938 1178 942
rect 1350 938 1354 942
rect 1526 938 1530 942
rect 2062 938 2066 942
rect 2198 938 2202 942
rect 2214 938 2218 942
rect 2646 948 2650 952
rect 2662 948 2666 952
rect 2782 948 2786 952
rect 2974 948 2978 952
rect 3526 948 3530 952
rect 4006 948 4010 952
rect 2526 938 2530 942
rect 3030 938 3034 942
rect 3278 938 3282 942
rect 3414 938 3418 942
rect 3790 938 3794 942
rect 3830 938 3834 942
rect 3918 938 3922 942
rect 4670 948 4674 952
rect 4694 948 4698 952
rect 4710 948 4714 952
rect 4774 948 4778 952
rect 4902 948 4906 952
rect 4198 938 4202 942
rect 4510 938 4514 942
rect 4782 938 4786 942
rect 5006 938 5010 942
rect 5166 938 5170 942
rect 246 928 250 932
rect 262 928 266 932
rect 646 928 650 932
rect 1086 928 1090 932
rect 1486 928 1490 932
rect 1678 928 1682 932
rect 2350 928 2354 932
rect 2382 928 2386 932
rect 2654 928 2658 932
rect 2966 928 2970 932
rect 3470 928 3474 932
rect 3806 928 3810 932
rect 4038 928 4042 932
rect 4150 928 4154 932
rect 4358 928 4362 932
rect 5062 928 5066 932
rect 5126 928 5130 932
rect 806 918 810 922
rect 1158 918 1162 922
rect 1726 918 1730 922
rect 2150 918 2154 922
rect 2838 918 2842 922
rect 3358 918 3362 922
rect 886 908 890 912
rect 894 908 898 912
rect 1198 908 1202 912
rect 1278 908 1282 912
rect 1342 908 1346 912
rect 1774 908 1778 912
rect 2206 908 2210 912
rect 2478 908 2482 912
rect 3078 908 3082 912
rect 3206 908 3210 912
rect 4102 908 4106 912
rect 4198 908 4202 912
rect 4470 908 4474 912
rect 4502 908 4506 912
rect 4718 908 4722 912
rect 1050 903 1054 907
rect 1058 903 1061 907
rect 1061 903 1062 907
rect 2074 903 2078 907
rect 2082 903 2085 907
rect 2085 903 2086 907
rect 3098 903 3102 907
rect 3106 903 3109 907
rect 3109 903 3110 907
rect 4114 903 4118 907
rect 4122 903 4125 907
rect 4125 903 4126 907
rect 558 898 562 902
rect 1230 898 1234 902
rect 1390 898 1394 902
rect 1526 898 1530 902
rect 2310 898 2314 902
rect 2630 898 2634 902
rect 2870 898 2874 902
rect 3030 898 3034 902
rect 3710 898 3714 902
rect 358 888 362 892
rect 422 888 426 892
rect 1206 888 1210 892
rect 2086 888 2090 892
rect 2110 888 2114 892
rect 2462 888 2466 892
rect 2638 888 2642 892
rect 3246 888 3250 892
rect 3510 888 3514 892
rect 4246 888 4250 892
rect 4478 888 4482 892
rect 4486 888 4490 892
rect 206 878 210 882
rect 326 878 330 882
rect 974 878 978 882
rect 1102 878 1106 882
rect 1254 878 1258 882
rect 1638 878 1642 882
rect 2150 878 2154 882
rect 2366 878 2370 882
rect 2814 878 2818 882
rect 3926 878 3930 882
rect 4206 878 4210 882
rect 4454 878 4458 882
rect 4694 878 4698 882
rect 4726 878 4730 882
rect 126 868 130 872
rect 606 868 610 872
rect 814 868 818 872
rect 1702 868 1706 872
rect 1718 868 1722 872
rect 1798 868 1802 872
rect 1822 868 1826 872
rect 2134 868 2138 872
rect 2894 868 2898 872
rect 2950 868 2954 872
rect 3006 868 3010 872
rect 3302 868 3306 872
rect 3342 868 3346 872
rect 3374 868 3378 872
rect 3734 868 3738 872
rect 3950 868 3954 872
rect 3982 868 3986 872
rect 590 858 594 862
rect 790 858 794 862
rect 958 858 962 862
rect 1086 858 1090 862
rect 1238 858 1242 862
rect 1422 858 1426 862
rect 1702 858 1706 862
rect 1838 858 1842 862
rect 1950 858 1954 862
rect 2534 858 2538 862
rect 2630 858 2634 862
rect 3166 858 3170 862
rect 3262 858 3266 862
rect 3270 858 3274 862
rect 3294 858 3298 862
rect 3438 858 3442 862
rect 3926 858 3930 862
rect 3974 858 3978 862
rect 4366 858 4370 862
rect 4558 858 4562 862
rect 4854 858 4858 862
rect 798 848 802 852
rect 886 848 890 852
rect 1550 848 1554 852
rect 1598 848 1602 852
rect 1606 848 1610 852
rect 1638 848 1642 852
rect 1766 848 1770 852
rect 2022 848 2026 852
rect 2214 848 2218 852
rect 2334 848 2338 852
rect 2518 848 2522 852
rect 2606 848 2610 852
rect 2646 848 2650 852
rect 3238 848 3242 852
rect 3870 848 3874 852
rect 4062 848 4066 852
rect 4694 848 4698 852
rect 5182 848 5186 852
rect 406 838 410 842
rect 1630 838 1634 842
rect 2062 838 2066 842
rect 2766 838 2770 842
rect 3278 838 3282 842
rect 3694 838 3698 842
rect 3830 838 3834 842
rect 4246 838 4250 842
rect 4470 838 4474 842
rect 454 828 458 832
rect 918 828 922 832
rect 1414 828 1418 832
rect 1726 828 1730 832
rect 1822 828 1826 832
rect 1846 828 1850 832
rect 2702 828 2706 832
rect 2822 828 2826 832
rect 3446 828 3450 832
rect 3454 828 3458 832
rect 3542 828 3546 832
rect 4486 828 4490 832
rect 4622 828 4626 832
rect 4790 828 4794 832
rect 190 818 194 822
rect 366 818 370 822
rect 614 818 618 822
rect 934 818 938 822
rect 1438 818 1442 822
rect 2270 818 2274 822
rect 2502 818 2506 822
rect 4022 818 4026 822
rect 4270 818 4274 822
rect 438 808 442 812
rect 830 808 834 812
rect 1542 808 1546 812
rect 2350 808 2354 812
rect 2606 808 2610 812
rect 3542 808 3546 812
rect 3630 808 3634 812
rect 3854 808 3858 812
rect 4294 808 4298 812
rect 4302 808 4306 812
rect 538 803 542 807
rect 546 803 549 807
rect 549 803 550 807
rect 1562 803 1566 807
rect 1570 803 1573 807
rect 1573 803 1574 807
rect 2586 803 2590 807
rect 2594 803 2597 807
rect 2597 803 2598 807
rect 3610 803 3614 807
rect 3618 803 3621 807
rect 3621 803 3622 807
rect 4634 803 4638 807
rect 4642 803 4645 807
rect 4645 803 4646 807
rect 366 798 370 802
rect 950 798 954 802
rect 1182 798 1186 802
rect 2126 798 2130 802
rect 2502 798 2506 802
rect 2950 798 2954 802
rect 3774 798 3778 802
rect 3782 798 3786 802
rect 4518 798 4522 802
rect 918 788 922 792
rect 1238 788 1242 792
rect 1478 788 1482 792
rect 3182 788 3186 792
rect 4302 788 4306 792
rect 4654 788 4658 792
rect 4806 788 4810 792
rect 5022 788 5026 792
rect 214 778 218 782
rect 910 778 914 782
rect 1286 778 1290 782
rect 1662 778 1666 782
rect 2286 778 2290 782
rect 2334 778 2338 782
rect 3070 778 3074 782
rect 3518 778 3522 782
rect 510 768 514 772
rect 902 768 906 772
rect 1422 768 1426 772
rect 1430 768 1434 772
rect 3174 768 3178 772
rect 3438 768 3442 772
rect 4430 768 4434 772
rect 822 758 826 762
rect 998 758 1002 762
rect 1070 758 1074 762
rect 1638 758 1642 762
rect 2438 758 2442 762
rect 2806 758 2810 762
rect 3134 758 3138 762
rect 3158 758 3162 762
rect 3246 758 3250 762
rect 3822 758 3826 762
rect 4326 758 4330 762
rect 4390 758 4394 762
rect 4518 758 4522 762
rect 230 748 234 752
rect 238 748 242 752
rect 702 748 706 752
rect 750 748 754 752
rect 774 748 778 752
rect 1094 748 1098 752
rect 1254 748 1258 752
rect 1670 748 1674 752
rect 1694 748 1698 752
rect 2118 748 2122 752
rect 2302 748 2306 752
rect 2518 748 2522 752
rect 2614 748 2618 752
rect 2790 748 2794 752
rect 2950 748 2954 752
rect 3206 748 3210 752
rect 3262 748 3266 752
rect 3294 748 3298 752
rect 3718 748 3722 752
rect 3774 748 3778 752
rect 3830 748 3834 752
rect 3934 748 3938 752
rect 3958 748 3962 752
rect 4006 748 4010 752
rect 4014 748 4018 752
rect 4310 748 4314 752
rect 4366 748 4370 752
rect 4518 748 4522 752
rect 4806 748 4810 752
rect 310 738 314 742
rect 462 738 466 742
rect 630 738 634 742
rect 662 738 666 742
rect 998 738 1002 742
rect 1054 738 1058 742
rect 1110 738 1114 742
rect 1118 738 1122 742
rect 1174 738 1178 742
rect 1358 738 1362 742
rect 1814 738 1818 742
rect 2246 738 2250 742
rect 2358 738 2362 742
rect 2622 738 2626 742
rect 3070 738 3074 742
rect 3366 738 3370 742
rect 3726 738 3730 742
rect 3838 738 3842 742
rect 4662 738 4666 742
rect 5062 738 5066 742
rect 270 728 274 732
rect 590 728 594 732
rect 678 728 682 732
rect 782 728 786 732
rect 1134 728 1138 732
rect 1398 728 1402 732
rect 1406 728 1410 732
rect 2270 728 2274 732
rect 3022 728 3026 732
rect 4278 728 4282 732
rect 4350 728 4354 732
rect 4558 728 4562 732
rect 5038 728 5042 732
rect 878 718 882 722
rect 1342 718 1346 722
rect 1494 718 1498 722
rect 2422 718 2426 722
rect 2686 718 2690 722
rect 2870 718 2874 722
rect 3102 718 3106 722
rect 4190 718 4194 722
rect 4374 718 4378 722
rect 102 708 106 712
rect 966 708 970 712
rect 974 708 978 712
rect 1086 708 1090 712
rect 1278 708 1282 712
rect 1390 708 1394 712
rect 1622 708 1626 712
rect 1854 708 1858 712
rect 2302 708 2306 712
rect 2902 708 2906 712
rect 3150 708 3154 712
rect 3814 708 3818 712
rect 4286 708 4290 712
rect 4766 708 4770 712
rect 4886 708 4890 712
rect 262 698 266 702
rect 1050 703 1054 707
rect 1058 703 1061 707
rect 1061 703 1062 707
rect 2074 703 2078 707
rect 2082 703 2085 707
rect 2085 703 2086 707
rect 3098 703 3102 707
rect 3106 703 3109 707
rect 3109 703 3110 707
rect 4114 703 4118 707
rect 4122 703 4125 707
rect 4125 703 4126 707
rect 1342 698 1346 702
rect 1446 698 1450 702
rect 1622 698 1626 702
rect 1638 698 1642 702
rect 1758 698 1762 702
rect 2062 698 2066 702
rect 2110 698 2114 702
rect 2318 698 2322 702
rect 2910 698 2914 702
rect 3086 698 3090 702
rect 3494 698 3498 702
rect 4590 698 4594 702
rect 4750 698 4754 702
rect 4918 698 4922 702
rect 222 688 226 692
rect 1078 688 1082 692
rect 1774 688 1778 692
rect 2174 688 2178 692
rect 2918 688 2922 692
rect 4014 688 4018 692
rect 4030 688 4034 692
rect 4062 688 4066 692
rect 398 678 402 682
rect 446 678 450 682
rect 982 678 986 682
rect 1222 678 1226 682
rect 1422 678 1426 682
rect 1998 678 2002 682
rect 2014 678 2018 682
rect 2206 678 2210 682
rect 2758 678 2762 682
rect 3182 678 3186 682
rect 4614 678 4618 682
rect 294 668 298 672
rect 398 668 402 672
rect 582 668 586 672
rect 790 668 794 672
rect 830 668 834 672
rect 910 668 914 672
rect 1174 668 1178 672
rect 1686 668 1690 672
rect 1766 668 1770 672
rect 2038 668 2042 672
rect 2374 668 2378 672
rect 2654 668 2658 672
rect 2902 668 2906 672
rect 2934 668 2938 672
rect 3006 668 3010 672
rect 3062 668 3066 672
rect 3158 668 3162 672
rect 3214 668 3218 672
rect 4046 668 4050 672
rect 4630 668 4634 672
rect 214 658 218 662
rect 414 658 418 662
rect 478 658 482 662
rect 710 658 714 662
rect 1022 658 1026 662
rect 1414 658 1418 662
rect 1454 658 1458 662
rect 1670 658 1674 662
rect 1758 658 1762 662
rect 1862 658 1866 662
rect 2366 658 2370 662
rect 2630 658 2634 662
rect 2926 658 2930 662
rect 3166 658 3170 662
rect 3198 658 3202 662
rect 3318 658 3322 662
rect 3950 658 3954 662
rect 4046 658 4050 662
rect 4446 658 4450 662
rect 4750 658 4754 662
rect 4982 658 4986 662
rect 966 648 970 652
rect 1630 648 1634 652
rect 1998 648 2002 652
rect 2142 648 2146 652
rect 2262 648 2266 652
rect 3254 648 3258 652
rect 3518 648 3522 652
rect 4070 648 4074 652
rect 4598 648 4602 652
rect 478 638 482 642
rect 870 638 874 642
rect 1518 638 1522 642
rect 3190 638 3194 642
rect 3254 638 3258 642
rect 3502 638 3506 642
rect 822 628 826 632
rect 1990 628 1994 632
rect 2622 628 2626 632
rect 2750 628 2754 632
rect 3014 628 3018 632
rect 3862 628 3866 632
rect 422 618 426 622
rect 1366 618 1370 622
rect 1814 618 1818 622
rect 2846 618 2850 622
rect 3950 618 3954 622
rect 4022 618 4026 622
rect 4622 618 4626 622
rect 4654 618 4658 622
rect 998 608 1002 612
rect 3566 608 3570 612
rect 3726 608 3730 612
rect 3790 608 3794 612
rect 3926 608 3930 612
rect 4454 608 4458 612
rect 538 603 542 607
rect 546 603 549 607
rect 549 603 550 607
rect 1562 603 1566 607
rect 1570 603 1573 607
rect 1573 603 1574 607
rect 2586 603 2590 607
rect 2594 603 2597 607
rect 2597 603 2598 607
rect 3610 603 3614 607
rect 3618 603 3621 607
rect 3621 603 3622 607
rect 4634 603 4638 607
rect 4642 603 4645 607
rect 4645 603 4646 607
rect 1678 598 1682 602
rect 4094 598 4098 602
rect 1014 588 1018 592
rect 1974 588 1978 592
rect 2030 588 2034 592
rect 2990 588 2994 592
rect 3566 588 3570 592
rect 3838 588 3842 592
rect 3846 588 3850 592
rect 3950 588 3954 592
rect 4926 588 4930 592
rect 622 578 626 582
rect 2062 578 2066 582
rect 2726 578 2730 582
rect 2974 578 2978 582
rect 4766 578 4770 582
rect 454 568 458 572
rect 1190 568 1194 572
rect 3582 568 3586 572
rect 3646 568 3650 572
rect 3806 568 3810 572
rect 262 558 266 562
rect 886 558 890 562
rect 910 558 914 562
rect 934 558 938 562
rect 950 558 954 562
rect 1030 558 1034 562
rect 1486 558 1490 562
rect 2022 558 2026 562
rect 2966 558 2970 562
rect 3470 558 3474 562
rect 3574 558 3578 562
rect 4094 558 4098 562
rect 94 548 98 552
rect 190 548 194 552
rect 206 548 210 552
rect 614 548 618 552
rect 870 548 874 552
rect 1014 548 1018 552
rect 1070 548 1074 552
rect 1142 548 1146 552
rect 1270 548 1274 552
rect 1550 548 1554 552
rect 1622 548 1626 552
rect 1702 548 1706 552
rect 1734 548 1738 552
rect 2246 548 2250 552
rect 126 538 130 542
rect 566 538 570 542
rect 630 538 634 542
rect 686 538 690 542
rect 718 538 722 542
rect 854 538 858 542
rect 862 538 866 542
rect 934 538 938 542
rect 1014 538 1018 542
rect 1030 538 1034 542
rect 1070 538 1074 542
rect 1958 538 1962 542
rect 2126 538 2130 542
rect 2806 548 2810 552
rect 2854 548 2858 552
rect 2958 548 2962 552
rect 3182 548 3186 552
rect 3422 548 3426 552
rect 3518 548 3522 552
rect 3558 548 3562 552
rect 3662 548 3666 552
rect 4030 548 4034 552
rect 4054 548 4058 552
rect 4102 548 4106 552
rect 4182 548 4186 552
rect 4414 548 4418 552
rect 4518 548 4522 552
rect 4598 548 4602 552
rect 2294 538 2298 542
rect 3254 538 3258 542
rect 3310 538 3314 542
rect 3342 538 3346 542
rect 3438 538 3442 542
rect 3446 538 3450 542
rect 3998 538 4002 542
rect 4206 538 4210 542
rect 4294 538 4298 542
rect 4422 538 4426 542
rect 4446 538 4450 542
rect 4622 538 4626 542
rect 4654 538 4658 542
rect 4742 538 4746 542
rect 4862 538 4866 542
rect 5054 538 5058 542
rect 86 528 90 532
rect 158 528 162 532
rect 1198 528 1202 532
rect 1302 528 1306 532
rect 3582 528 3586 532
rect 4478 528 4482 532
rect 766 518 770 522
rect 846 518 850 522
rect 886 518 890 522
rect 1758 518 1762 522
rect 2310 518 2314 522
rect 2814 518 2818 522
rect 2934 518 2938 522
rect 2990 518 2994 522
rect 3526 518 3530 522
rect 4134 518 4138 522
rect 4494 518 4498 522
rect 4750 518 4754 522
rect 638 508 642 512
rect 646 508 650 512
rect 1230 508 1234 512
rect 1806 508 1810 512
rect 3414 508 3418 512
rect 3454 508 3458 512
rect 3478 508 3482 512
rect 3686 508 3690 512
rect 1050 503 1054 507
rect 1058 503 1061 507
rect 1061 503 1062 507
rect 2074 503 2078 507
rect 2082 503 2085 507
rect 2085 503 2086 507
rect 3098 503 3102 507
rect 3106 503 3109 507
rect 3109 503 3110 507
rect 4114 503 4118 507
rect 4122 503 4125 507
rect 4125 503 4126 507
rect 590 498 594 502
rect 774 498 778 502
rect 3174 498 3178 502
rect 4358 498 4362 502
rect 1190 488 1194 492
rect 1438 488 1442 492
rect 1494 488 1498 492
rect 1734 488 1738 492
rect 2270 488 2274 492
rect 2350 488 2354 492
rect 2998 488 3002 492
rect 3574 488 3578 492
rect 3870 488 3874 492
rect 4470 488 4474 492
rect 4486 488 4490 492
rect 822 478 826 482
rect 926 478 930 482
rect 1470 478 1474 482
rect 1782 478 1786 482
rect 1822 478 1826 482
rect 2046 478 2050 482
rect 2342 478 2346 482
rect 2646 478 2650 482
rect 2670 478 2674 482
rect 2718 478 2722 482
rect 3406 478 3410 482
rect 4734 478 4738 482
rect 358 468 362 472
rect 406 468 410 472
rect 430 468 434 472
rect 486 468 490 472
rect 694 468 698 472
rect 782 468 786 472
rect 926 468 930 472
rect 1038 468 1042 472
rect 1134 468 1138 472
rect 1214 468 1218 472
rect 1278 468 1282 472
rect 1510 468 1514 472
rect 1766 468 1770 472
rect 2398 468 2402 472
rect 2422 468 2426 472
rect 2654 468 2658 472
rect 2830 468 2834 472
rect 2878 468 2882 472
rect 2966 468 2970 472
rect 3430 468 3434 472
rect 4086 468 4090 472
rect 4182 468 4186 472
rect 4198 468 4202 472
rect 4318 468 4322 472
rect 4326 468 4330 472
rect 4390 468 4394 472
rect 182 458 186 462
rect 398 458 402 462
rect 454 458 458 462
rect 614 458 618 462
rect 814 458 818 462
rect 958 458 962 462
rect 1006 458 1010 462
rect 1694 458 1698 462
rect 1726 458 1730 462
rect 2022 458 2026 462
rect 2278 458 2282 462
rect 3310 458 3314 462
rect 4014 458 4018 462
rect 4806 458 4810 462
rect 238 448 242 452
rect 342 448 346 452
rect 638 448 642 452
rect 182 438 186 442
rect 1030 448 1034 452
rect 2382 448 2386 452
rect 2494 448 2498 452
rect 3718 448 3722 452
rect 3878 448 3882 452
rect 4414 448 4418 452
rect 4526 448 4530 452
rect 4534 448 4538 452
rect 678 438 682 442
rect 1518 438 1522 442
rect 2790 438 2794 442
rect 3438 438 3442 442
rect 4366 438 4370 442
rect 774 428 778 432
rect 1422 428 1426 432
rect 1454 428 1458 432
rect 3134 428 3138 432
rect 2054 418 2058 422
rect 2094 418 2098 422
rect 3798 418 3802 422
rect 4406 418 4410 422
rect 4742 418 4746 422
rect 766 408 770 412
rect 798 408 802 412
rect 1430 408 1434 412
rect 1910 408 1914 412
rect 2334 408 2338 412
rect 2654 408 2658 412
rect 2702 408 2706 412
rect 2846 408 2850 412
rect 2998 408 3002 412
rect 538 403 542 407
rect 546 403 549 407
rect 549 403 550 407
rect 1562 403 1566 407
rect 1570 403 1573 407
rect 1573 403 1574 407
rect 2586 403 2590 407
rect 2594 403 2597 407
rect 2597 403 2598 407
rect 3610 403 3614 407
rect 3618 403 3621 407
rect 3621 403 3622 407
rect 4634 403 4638 407
rect 4642 403 4645 407
rect 4645 403 4646 407
rect 1014 398 1018 402
rect 1174 398 1178 402
rect 1230 398 1234 402
rect 1254 398 1258 402
rect 2110 398 2114 402
rect 2774 398 2778 402
rect 2846 398 2850 402
rect 3470 398 3474 402
rect 3646 398 3650 402
rect 3678 398 3682 402
rect 3846 398 3850 402
rect 4382 398 4386 402
rect 158 388 162 392
rect 174 388 178 392
rect 1086 388 1090 392
rect 1462 388 1466 392
rect 2350 388 2354 392
rect 2718 388 2722 392
rect 3006 388 3010 392
rect 3118 388 3122 392
rect 3294 388 3298 392
rect 4422 388 4426 392
rect 1270 378 1274 382
rect 1758 378 1762 382
rect 3454 378 3458 382
rect 3982 378 3986 382
rect 4686 378 4690 382
rect 414 368 418 372
rect 814 368 818 372
rect 974 368 978 372
rect 1078 368 1082 372
rect 1222 368 1226 372
rect 1238 368 1242 372
rect 1294 368 1298 372
rect 1334 368 1338 372
rect 1422 368 1426 372
rect 1734 368 1738 372
rect 2262 368 2266 372
rect 1534 358 1538 362
rect 1702 358 1706 362
rect 2862 368 2866 372
rect 3022 368 3026 372
rect 3334 368 3338 372
rect 3678 368 3682 372
rect 3854 368 3858 372
rect 2718 358 2722 362
rect 2950 358 2954 362
rect 3902 358 3906 362
rect 4030 358 4034 362
rect 4070 358 4074 362
rect 4566 368 4570 372
rect 4854 368 4858 372
rect 4918 368 4922 372
rect 4358 358 4362 362
rect 4518 358 4522 362
rect 206 348 210 352
rect 342 348 346 352
rect 606 348 610 352
rect 1438 348 1442 352
rect 1502 348 1506 352
rect 1934 348 1938 352
rect 2014 348 2018 352
rect 2678 348 2682 352
rect 102 338 106 342
rect 406 338 410 342
rect 3310 348 3314 352
rect 3462 348 3466 352
rect 3798 348 3802 352
rect 3878 348 3882 352
rect 3966 348 3970 352
rect 4134 348 4138 352
rect 4206 348 4210 352
rect 4478 348 4482 352
rect 4534 348 4538 352
rect 4558 348 4562 352
rect 574 338 578 342
rect 670 338 674 342
rect 862 338 866 342
rect 1118 338 1122 342
rect 2286 338 2290 342
rect 2982 338 2986 342
rect 3254 338 3258 342
rect 3366 338 3370 342
rect 3870 338 3874 342
rect 4198 338 4202 342
rect 4470 338 4474 342
rect 4758 338 4762 342
rect 166 328 170 332
rect 182 328 186 332
rect 1086 328 1090 332
rect 2734 328 2738 332
rect 2894 328 2898 332
rect 3326 328 3330 332
rect 3334 328 3338 332
rect 3838 328 3842 332
rect 574 318 578 322
rect 598 318 602 322
rect 1446 318 1450 322
rect 1470 318 1474 322
rect 1726 318 1730 322
rect 4814 318 4818 322
rect 1270 308 1274 312
rect 1958 308 1962 312
rect 2870 308 2874 312
rect 3126 308 3130 312
rect 3662 308 3666 312
rect 1050 303 1054 307
rect 1058 303 1061 307
rect 1061 303 1062 307
rect 2074 303 2078 307
rect 2082 303 2085 307
rect 2085 303 2086 307
rect 3098 303 3102 307
rect 3106 303 3109 307
rect 3109 303 3110 307
rect 4114 303 4118 307
rect 4122 303 4125 307
rect 4125 303 4126 307
rect 174 298 178 302
rect 1302 298 1306 302
rect 1950 298 1954 302
rect 2438 298 2442 302
rect 2870 298 2874 302
rect 4694 298 4698 302
rect 750 288 754 292
rect 1270 288 1274 292
rect 1534 288 1538 292
rect 1718 288 1722 292
rect 2182 288 2186 292
rect 3294 288 3298 292
rect 3750 288 3754 292
rect 5190 288 5194 292
rect 750 278 754 282
rect 1310 278 1314 282
rect 1358 278 1362 282
rect 1470 278 1474 282
rect 3022 278 3026 282
rect 3478 278 3482 282
rect 4854 278 4858 282
rect 446 268 450 272
rect 462 268 466 272
rect 662 268 666 272
rect 694 268 698 272
rect 1078 268 1082 272
rect 1270 268 1274 272
rect 1350 268 1354 272
rect 1406 268 1410 272
rect 1502 268 1506 272
rect 1526 268 1530 272
rect 1590 268 1594 272
rect 1742 268 1746 272
rect 1926 268 1930 272
rect 2014 268 2018 272
rect 2702 268 2706 272
rect 2726 268 2730 272
rect 2774 268 2778 272
rect 3366 268 3370 272
rect 4174 268 4178 272
rect 4454 268 4458 272
rect 4470 268 4474 272
rect 4766 268 4770 272
rect 5118 268 5122 272
rect 134 258 138 262
rect 838 258 842 262
rect 1302 258 1306 262
rect 1622 258 1626 262
rect 1734 258 1738 262
rect 1878 258 1882 262
rect 2166 258 2170 262
rect 2214 258 2218 262
rect 2238 258 2242 262
rect 2566 258 2570 262
rect 2958 258 2962 262
rect 3310 258 3314 262
rect 4374 258 4378 262
rect 4446 258 4450 262
rect 4870 258 4874 262
rect 5134 258 5138 262
rect 550 248 554 252
rect 1910 248 1914 252
rect 3174 248 3178 252
rect 806 238 810 242
rect 1054 238 1058 242
rect 1486 238 1490 242
rect 3750 248 3754 252
rect 3998 248 4002 252
rect 4710 248 4714 252
rect 4758 248 4762 252
rect 2814 238 2818 242
rect 3462 238 3466 242
rect 3886 238 3890 242
rect 4878 238 4882 242
rect 670 228 674 232
rect 918 228 922 232
rect 1310 228 1314 232
rect 1990 228 1994 232
rect 2382 228 2386 232
rect 4622 228 4626 232
rect 646 218 650 222
rect 1582 218 1586 222
rect 1750 218 1754 222
rect 2862 218 2866 222
rect 3030 218 3034 222
rect 4238 218 4242 222
rect 5070 218 5074 222
rect 1502 208 1506 212
rect 2182 208 2186 212
rect 2694 208 2698 212
rect 3654 208 3658 212
rect 4606 208 4610 212
rect 538 203 542 207
rect 546 203 549 207
rect 549 203 550 207
rect 1562 203 1566 207
rect 1570 203 1573 207
rect 1573 203 1574 207
rect 2586 203 2590 207
rect 2594 203 2597 207
rect 2597 203 2598 207
rect 222 198 226 202
rect 1110 198 1114 202
rect 1662 198 1666 202
rect 2726 198 2730 202
rect 3610 203 3614 207
rect 3618 203 3621 207
rect 3621 203 3622 207
rect 4634 203 4638 207
rect 4642 203 4645 207
rect 4645 203 4646 207
rect 4102 198 4106 202
rect 4414 198 4418 202
rect 1582 188 1586 192
rect 1878 188 1882 192
rect 1918 188 1922 192
rect 3326 188 3330 192
rect 4494 188 4498 192
rect 4750 188 4754 192
rect 5102 188 5106 192
rect 1734 178 1738 182
rect 3398 178 3402 182
rect 3862 178 3866 182
rect 4182 178 4186 182
rect 966 168 970 172
rect 1454 168 1458 172
rect 1774 168 1778 172
rect 2158 168 2162 172
rect 2494 168 2498 172
rect 2742 168 2746 172
rect 2750 168 2754 172
rect 2846 168 2850 172
rect 4006 168 4010 172
rect 4446 168 4450 172
rect 4822 168 4826 172
rect 534 158 538 162
rect 1806 158 1810 162
rect 2854 158 2858 162
rect 2862 158 2866 162
rect 214 148 218 152
rect 342 148 346 152
rect 782 148 786 152
rect 1446 148 1450 152
rect 1494 148 1498 152
rect 230 138 234 142
rect 694 138 698 142
rect 798 138 802 142
rect 1254 138 1258 142
rect 1558 148 1562 152
rect 1742 148 1746 152
rect 1750 148 1754 152
rect 1862 148 1866 152
rect 1870 148 1874 152
rect 2022 148 2026 152
rect 2510 148 2514 152
rect 2702 148 2706 152
rect 3206 148 3210 152
rect 3310 148 3314 152
rect 3494 148 3498 152
rect 4438 148 4442 152
rect 4518 148 4522 152
rect 4758 148 4762 152
rect 4830 148 4834 152
rect 5174 148 5178 152
rect 1430 138 1434 142
rect 1462 138 1466 142
rect 1590 138 1594 142
rect 1758 138 1762 142
rect 1878 138 1882 142
rect 1934 138 1938 142
rect 2182 138 2186 142
rect 2286 138 2290 142
rect 2854 138 2858 142
rect 3414 138 3418 142
rect 3790 138 3794 142
rect 4206 138 4210 142
rect 4222 138 4226 142
rect 4382 138 4386 142
rect 4742 138 4746 142
rect 4798 138 4802 142
rect 4854 138 4858 142
rect 4966 138 4970 142
rect 758 128 762 132
rect 1718 128 1722 132
rect 1806 128 1810 132
rect 2582 128 2586 132
rect 2742 128 2746 132
rect 3566 128 3570 132
rect 3822 128 3826 132
rect 4470 128 4474 132
rect 4574 128 4578 132
rect 4758 128 4762 132
rect 798 118 802 122
rect 1918 118 1922 122
rect 2366 118 2370 122
rect 5078 118 5082 122
rect 766 108 770 112
rect 1470 108 1474 112
rect 2814 108 2818 112
rect 2822 108 2826 112
rect 4022 108 4026 112
rect 4606 108 4610 112
rect 4894 108 4898 112
rect 1050 103 1054 107
rect 1058 103 1061 107
rect 1061 103 1062 107
rect 2074 103 2078 107
rect 2082 103 2085 107
rect 2085 103 2086 107
rect 3098 103 3102 107
rect 3106 103 3109 107
rect 3109 103 3110 107
rect 4114 103 4118 107
rect 4122 103 4125 107
rect 4125 103 4126 107
rect 742 98 746 102
rect 758 98 762 102
rect 4198 98 4202 102
rect 4958 98 4962 102
rect 638 88 642 92
rect 694 88 698 92
rect 1678 88 1682 92
rect 1774 88 1778 92
rect 1990 88 1994 92
rect 2742 88 2746 92
rect 2998 88 3002 92
rect 5006 88 5010 92
rect 758 78 762 82
rect 918 78 922 82
rect 1870 78 1874 82
rect 2566 78 2570 82
rect 2686 78 2690 82
rect 3310 78 3314 82
rect 3662 78 3666 82
rect 4398 78 4402 82
rect 4942 78 4946 82
rect 4958 78 4962 82
rect 4998 78 5002 82
rect 982 68 986 72
rect 3654 68 3658 72
rect 3942 68 3946 72
rect 4214 68 4218 72
rect 5158 68 5162 72
rect 350 58 354 62
rect 798 58 802 62
rect 942 58 946 62
rect 1310 58 1314 62
rect 1462 58 1466 62
rect 1558 58 1562 62
rect 2278 58 2282 62
rect 2374 58 2378 62
rect 2758 58 2762 62
rect 3406 58 3410 62
rect 3822 58 3826 62
rect 4542 58 4546 62
rect 4582 58 4586 62
rect 4686 58 4690 62
rect 4750 58 4754 62
rect 4846 58 4850 62
rect 4990 58 4994 62
rect 1910 48 1914 52
rect 2646 48 2650 52
rect 3510 48 3514 52
rect 3998 48 4002 52
rect 4038 48 4042 52
rect 4086 48 4090 52
rect 4118 48 4122 52
rect 4550 48 4554 52
rect 4814 48 4818 52
rect 3222 8 3226 12
rect 538 3 542 7
rect 546 3 549 7
rect 549 3 550 7
rect 1562 3 1566 7
rect 1570 3 1573 7
rect 1573 3 1574 7
rect 2586 3 2590 7
rect 2594 3 2597 7
rect 2597 3 2598 7
rect 3610 3 3614 7
rect 3618 3 3621 7
rect 3621 3 3622 7
rect 4634 3 4638 7
rect 4642 3 4645 7
rect 4645 3 4646 7
<< metal4 >>
rect 1048 4903 1050 4907
rect 1054 4903 1057 4907
rect 1062 4903 1064 4907
rect 2072 4903 2074 4907
rect 2078 4903 2081 4907
rect 2086 4903 2088 4907
rect 3096 4903 3098 4907
rect 3102 4903 3105 4907
rect 3110 4903 3112 4907
rect 4112 4903 4114 4907
rect 4118 4903 4121 4907
rect 4126 4903 4128 4907
rect 582 4862 585 4868
rect 536 4803 538 4807
rect 542 4803 545 4807
rect 550 4803 552 4807
rect 94 3962 97 4368
rect 102 4062 105 4408
rect 110 4262 113 4478
rect 134 4222 137 4688
rect 150 4652 153 4658
rect 6 3512 9 3548
rect 94 3352 97 3958
rect 102 3762 105 4058
rect 142 4012 145 4318
rect 174 3952 177 4758
rect 250 4458 257 4461
rect 126 3262 129 3908
rect 134 3362 137 3948
rect 166 3662 169 3938
rect 118 3258 126 3261
rect 6 2742 9 3248
rect 18 3148 22 3151
rect 102 2872 105 3148
rect 118 3112 121 3258
rect 142 2562 145 3498
rect 174 3482 177 3948
rect 246 3482 249 4348
rect 254 4162 257 4458
rect 262 4342 265 4708
rect 286 4372 289 4578
rect 294 4362 297 4718
rect 342 4662 345 4678
rect 422 4658 430 4661
rect 422 4652 425 4658
rect 486 4552 489 4738
rect 574 4712 577 4858
rect 750 4832 753 4868
rect 674 4748 678 4751
rect 494 4662 497 4688
rect 318 4522 321 4538
rect 274 4348 278 4351
rect 262 4192 265 4248
rect 166 3478 174 3481
rect 158 3322 161 3468
rect 166 3332 169 3478
rect 222 3272 225 3468
rect 230 3452 233 3478
rect 262 3452 265 4188
rect 270 4138 278 4141
rect 270 3962 273 4138
rect 302 4112 305 4148
rect 274 3858 278 3861
rect 302 3642 305 4108
rect 318 4062 321 4138
rect 334 4062 337 4268
rect 238 3332 241 3418
rect 174 3061 177 3068
rect 174 3058 182 3061
rect 202 2948 206 2951
rect 210 2678 214 2681
rect 10 2548 14 2551
rect 6 2492 9 2518
rect 14 2442 17 2508
rect 118 2462 121 2488
rect 10 2348 14 2351
rect 10 2328 14 2331
rect 94 2322 97 2348
rect 94 2132 97 2148
rect 74 2088 78 2091
rect 134 2062 137 2508
rect 166 2082 169 2088
rect 126 1402 129 1838
rect 102 972 105 1268
rect 134 1152 137 1158
rect 130 868 134 871
rect 94 531 97 548
rect 90 528 97 531
rect 102 342 105 708
rect 126 542 129 868
rect 158 392 161 528
rect 166 332 169 1218
rect 190 822 193 2658
rect 214 2111 217 2278
rect 214 2108 222 2111
rect 218 2088 225 2091
rect 222 1542 225 2088
rect 238 1792 241 2908
rect 246 2902 249 3028
rect 262 2222 265 3448
rect 270 3282 273 3538
rect 270 2672 273 3278
rect 310 2762 313 4058
rect 318 3742 321 4058
rect 270 2622 273 2668
rect 222 1272 225 1468
rect 218 1158 222 1161
rect 222 1062 225 1068
rect 238 992 241 1248
rect 246 932 249 1128
rect 206 552 209 878
rect 214 662 217 778
rect 194 548 198 551
rect 182 442 185 458
rect 174 302 177 388
rect 210 348 217 351
rect 186 328 190 331
rect 134 262 137 268
rect 214 152 217 348
rect 222 202 225 688
rect 218 148 222 151
rect 230 142 233 748
rect 238 452 241 748
rect 262 702 265 928
rect 270 732 273 2258
rect 286 2122 289 2148
rect 302 2102 305 2268
rect 294 1952 297 1958
rect 278 1518 286 1521
rect 278 1322 281 1518
rect 262 562 265 698
rect 294 672 297 1418
rect 302 1282 305 1958
rect 318 1462 321 3738
rect 326 3222 329 3938
rect 334 3262 337 4048
rect 342 3562 345 4138
rect 326 3158 334 3161
rect 326 3082 329 3158
rect 342 3072 345 3328
rect 326 2622 329 2648
rect 350 2462 353 4338
rect 358 3982 361 4178
rect 366 4152 369 4178
rect 382 4062 385 4168
rect 422 4142 425 4148
rect 430 4142 433 4268
rect 390 4082 393 4128
rect 382 4022 385 4038
rect 358 3772 361 3818
rect 358 3722 361 3768
rect 382 3752 385 4018
rect 382 3742 385 3748
rect 358 3552 361 3558
rect 382 3502 385 3698
rect 390 3632 393 4078
rect 406 3691 409 3958
rect 414 3872 417 3878
rect 402 3688 409 3691
rect 398 3452 401 3548
rect 374 3142 377 3158
rect 382 3142 385 3318
rect 366 2941 369 2988
rect 362 2938 369 2941
rect 378 2758 382 2761
rect 362 2688 366 2691
rect 382 2282 385 2318
rect 382 2152 385 2168
rect 326 882 329 1528
rect 334 1292 337 2138
rect 378 2048 382 2051
rect 390 1892 393 3138
rect 398 3062 401 3258
rect 398 1862 401 2858
rect 406 2852 409 3628
rect 422 3562 425 4138
rect 406 2462 409 2788
rect 414 2782 417 3538
rect 422 3332 425 3348
rect 430 3322 433 3868
rect 430 3102 433 3208
rect 438 2672 441 3928
rect 446 3652 449 4228
rect 486 4102 489 4548
rect 494 4072 497 4658
rect 536 4603 538 4607
rect 542 4603 545 4607
rect 550 4603 552 4607
rect 558 4582 561 4608
rect 536 4403 538 4407
rect 542 4403 545 4407
rect 550 4403 552 4407
rect 550 4262 553 4318
rect 536 4203 538 4207
rect 542 4203 545 4207
rect 550 4203 552 4207
rect 462 3662 465 3688
rect 478 3672 481 3678
rect 446 3472 449 3478
rect 418 2548 422 2551
rect 374 1738 382 1741
rect 362 1668 366 1671
rect 374 1642 377 1738
rect 358 1552 361 1638
rect 342 962 345 1338
rect 358 1322 361 1548
rect 378 1428 382 1431
rect 398 1422 401 1858
rect 406 1542 409 1618
rect 422 1612 425 2478
rect 358 1282 361 1318
rect 350 1258 358 1261
rect 350 982 353 1258
rect 374 1212 377 1418
rect 386 1258 390 1261
rect 358 892 361 1118
rect 398 1112 401 1208
rect 366 822 369 948
rect 366 802 369 818
rect 302 741 305 768
rect 302 738 310 741
rect 398 682 401 1108
rect 406 972 409 1538
rect 414 1472 417 1528
rect 430 1472 433 2458
rect 446 2252 449 3268
rect 470 3192 473 3638
rect 478 3322 481 3528
rect 438 2162 441 2218
rect 438 2062 441 2158
rect 446 2112 449 2208
rect 446 1852 449 2108
rect 446 1681 449 1818
rect 442 1678 449 1681
rect 454 1632 457 2928
rect 470 2392 473 2468
rect 470 2342 473 2388
rect 478 2272 481 2518
rect 486 2392 489 4008
rect 494 3481 497 4068
rect 502 3662 505 4078
rect 518 4072 521 4178
rect 502 3502 505 3658
rect 510 3522 513 4038
rect 566 4032 569 4668
rect 582 4312 585 4518
rect 590 4242 593 4408
rect 630 4342 633 4448
rect 536 4003 538 4007
rect 542 4003 545 4007
rect 550 4003 552 4007
rect 526 3782 529 3808
rect 536 3803 538 3807
rect 542 3803 545 3807
rect 550 3803 552 3807
rect 574 3702 577 4068
rect 536 3603 538 3607
rect 542 3603 545 3607
rect 550 3603 552 3607
rect 494 3478 505 3481
rect 494 3372 497 3468
rect 502 2772 505 3478
rect 536 3403 538 3407
rect 542 3403 545 3407
rect 550 3403 552 3407
rect 550 3362 553 3368
rect 518 3332 521 3338
rect 518 3072 521 3318
rect 550 3232 553 3358
rect 536 3203 538 3207
rect 542 3203 545 3207
rect 550 3203 552 3207
rect 498 2568 502 2571
rect 502 2532 505 2568
rect 510 2342 513 2758
rect 518 2542 521 3068
rect 536 3003 538 3007
rect 542 3003 545 3007
rect 550 3003 552 3007
rect 518 2522 521 2538
rect 470 1961 473 2218
rect 502 2112 505 2328
rect 482 2048 486 2051
rect 466 1958 473 1961
rect 482 1948 489 1951
rect 486 1922 489 1948
rect 462 1858 470 1861
rect 462 1832 465 1858
rect 462 1562 465 1828
rect 478 1742 481 1848
rect 434 1448 438 1451
rect 418 1388 425 1391
rect 414 1042 417 1348
rect 422 1332 425 1388
rect 422 1062 425 1078
rect 354 468 358 471
rect 398 462 401 668
rect 406 472 409 838
rect 342 352 345 448
rect 346 348 350 351
rect 342 152 345 348
rect 406 342 409 468
rect 414 372 417 658
rect 422 622 425 888
rect 438 812 441 1428
rect 446 1312 449 1458
rect 446 1272 449 1308
rect 454 832 457 1218
rect 462 1132 465 1328
rect 470 1252 473 1268
rect 470 1152 473 1158
rect 478 1092 481 1738
rect 462 872 465 988
rect 462 742 465 868
rect 426 468 430 471
rect 446 292 449 678
rect 478 642 481 658
rect 454 462 457 568
rect 486 472 489 1448
rect 494 1012 497 1878
rect 518 1632 521 2368
rect 526 2352 529 2938
rect 558 2832 561 3358
rect 566 2952 569 3208
rect 574 3062 577 3198
rect 536 2803 538 2807
rect 542 2803 545 2807
rect 550 2803 552 2807
rect 536 2603 538 2607
rect 542 2603 545 2607
rect 550 2603 552 2607
rect 546 2478 550 2481
rect 536 2403 538 2407
rect 542 2403 545 2407
rect 550 2403 552 2407
rect 536 2203 538 2207
rect 542 2203 545 2207
rect 550 2203 552 2207
rect 566 2122 569 2948
rect 574 2862 577 2868
rect 582 2752 585 4058
rect 590 3982 593 4238
rect 590 3962 593 3968
rect 578 2688 582 2691
rect 582 2652 585 2658
rect 590 2622 593 3728
rect 598 3532 601 4128
rect 610 4068 617 4071
rect 614 3642 617 4068
rect 630 4032 633 4288
rect 638 4272 641 4598
rect 610 3548 614 3551
rect 598 2612 601 3518
rect 606 3282 609 3538
rect 574 2572 577 2578
rect 526 1542 529 2038
rect 536 2003 538 2007
rect 542 2003 545 2007
rect 550 2003 552 2007
rect 558 1912 561 1938
rect 536 1803 538 1807
rect 542 1803 545 1807
rect 550 1803 552 1807
rect 536 1603 538 1607
rect 542 1603 545 1607
rect 550 1603 552 1607
rect 558 1462 561 1908
rect 574 1872 577 2528
rect 582 2342 585 2538
rect 594 2458 598 2461
rect 606 2361 609 2558
rect 614 2412 617 3438
rect 622 3142 625 3278
rect 622 2542 625 3058
rect 630 2922 633 4028
rect 646 3732 649 4738
rect 682 4708 689 4711
rect 654 4472 657 4638
rect 686 4522 689 4708
rect 710 4572 713 4818
rect 766 4742 769 4858
rect 758 4722 761 4738
rect 646 2962 649 3328
rect 654 2952 657 4468
rect 710 4332 713 4458
rect 670 4071 673 4218
rect 666 4068 673 4071
rect 670 3742 673 3838
rect 670 3702 673 3738
rect 678 3552 681 3578
rect 686 3552 689 3748
rect 682 3448 686 3451
rect 670 3282 673 3328
rect 662 3252 665 3278
rect 678 3142 681 3438
rect 694 3362 697 3648
rect 686 3052 689 3138
rect 654 2762 657 2928
rect 662 2902 665 2998
rect 694 2952 697 3258
rect 646 2648 654 2651
rect 646 2642 649 2648
rect 622 2402 625 2538
rect 630 2502 633 2508
rect 630 2402 633 2428
rect 602 2358 609 2361
rect 590 2182 593 2258
rect 606 2162 609 2358
rect 622 2262 625 2388
rect 622 2072 625 2258
rect 630 2162 633 2198
rect 638 2162 641 2548
rect 662 2422 665 2898
rect 678 2752 681 2948
rect 686 2671 689 2678
rect 682 2668 689 2671
rect 646 2162 649 2348
rect 654 2262 657 2278
rect 614 1952 617 1958
rect 574 1742 577 1868
rect 578 1668 582 1671
rect 536 1403 538 1407
rect 542 1403 545 1407
rect 550 1403 552 1407
rect 502 1382 505 1388
rect 526 1382 529 1398
rect 558 1342 561 1458
rect 570 1348 574 1351
rect 590 1322 593 1678
rect 606 1552 609 1888
rect 614 1562 617 1648
rect 598 1352 601 1418
rect 622 1402 625 1608
rect 630 1342 633 1468
rect 638 1452 641 2128
rect 646 1662 649 1898
rect 654 1762 657 2158
rect 638 1362 641 1368
rect 594 1268 598 1271
rect 536 1203 538 1207
rect 542 1203 545 1207
rect 550 1203 552 1207
rect 558 1042 561 1148
rect 536 1003 538 1007
rect 542 1003 545 1007
rect 550 1003 552 1007
rect 558 902 561 1038
rect 510 772 513 858
rect 536 803 538 807
rect 542 803 545 807
rect 550 803 552 807
rect 582 672 585 1148
rect 590 862 593 1248
rect 618 1128 622 1131
rect 590 732 593 838
rect 536 603 538 607
rect 542 603 545 607
rect 550 603 552 607
rect 566 522 569 538
rect 590 502 593 558
rect 536 403 538 407
rect 542 403 545 407
rect 550 403 552 407
rect 574 322 577 338
rect 598 332 601 978
rect 606 872 609 938
rect 606 352 609 868
rect 614 552 617 818
rect 630 742 633 1208
rect 646 932 649 1658
rect 654 1392 657 1508
rect 662 1472 665 2038
rect 670 1712 673 2628
rect 678 2042 681 2638
rect 694 2632 697 2948
rect 702 2682 705 4228
rect 718 4182 721 4708
rect 758 4542 761 4718
rect 878 4652 881 4668
rect 738 4538 742 4541
rect 714 3938 718 3941
rect 718 3422 721 3648
rect 726 3562 729 4458
rect 734 3952 737 4038
rect 734 3622 737 3948
rect 766 3862 769 4568
rect 822 4512 825 4568
rect 858 4528 862 4531
rect 854 4342 857 4528
rect 854 4318 862 4321
rect 766 3702 769 3818
rect 726 3412 729 3558
rect 714 3148 718 3151
rect 710 3092 713 3118
rect 670 1652 673 1698
rect 670 1532 673 1628
rect 654 952 657 1128
rect 662 982 665 1408
rect 670 1272 673 1488
rect 678 1342 681 2038
rect 686 2032 689 2528
rect 694 2212 697 2618
rect 702 2482 705 2678
rect 694 2142 697 2148
rect 686 1402 689 1898
rect 694 1642 697 1848
rect 702 1752 705 2448
rect 710 2152 713 3008
rect 718 2182 721 2418
rect 702 1662 705 1718
rect 702 1261 705 1628
rect 710 1282 713 1748
rect 718 1522 721 1708
rect 726 1542 729 3358
rect 734 3142 737 3148
rect 734 1752 737 2948
rect 742 2772 745 3338
rect 750 3222 753 3448
rect 766 3242 769 3638
rect 774 3482 777 4288
rect 774 3182 777 3478
rect 770 3158 774 3161
rect 758 3092 761 3138
rect 774 3062 777 3068
rect 774 2952 777 2968
rect 742 2572 745 2748
rect 742 2082 745 2378
rect 750 2062 753 2938
rect 762 2868 766 2871
rect 774 2822 777 2918
rect 782 2822 785 4268
rect 810 4258 814 4261
rect 854 4242 857 4318
rect 794 4148 798 4151
rect 794 4068 798 4071
rect 870 4062 873 4628
rect 878 4042 881 4268
rect 806 3452 809 3818
rect 794 2938 798 2941
rect 758 2122 761 2668
rect 734 1582 737 1598
rect 702 1258 710 1261
rect 622 462 625 578
rect 634 538 638 541
rect 638 512 641 528
rect 618 458 622 461
rect 598 322 601 328
rect 446 272 449 288
rect 458 268 462 271
rect 550 242 553 248
rect 536 203 538 207
rect 542 203 545 207
rect 550 203 552 207
rect 534 152 537 158
rect 638 92 641 448
rect 646 222 649 508
rect 662 272 665 738
rect 678 442 681 728
rect 686 542 689 1208
rect 710 1072 713 1258
rect 670 232 673 338
rect 686 271 689 518
rect 694 472 697 988
rect 706 938 710 941
rect 702 722 705 748
rect 710 622 713 658
rect 718 542 721 1348
rect 734 1142 737 1568
rect 742 1472 745 1998
rect 750 1471 753 2058
rect 774 1952 777 2818
rect 782 2582 785 2598
rect 782 2562 785 2568
rect 790 2552 793 2848
rect 782 2132 785 2318
rect 758 1871 761 1928
rect 790 1902 793 2548
rect 798 2412 801 2728
rect 806 2552 809 3218
rect 814 3172 817 4028
rect 854 3938 862 3941
rect 814 3132 817 3138
rect 814 3102 817 3108
rect 822 3072 825 3858
rect 830 3552 833 3568
rect 830 3162 833 3378
rect 838 2892 841 3778
rect 846 3072 849 3388
rect 854 3232 857 3938
rect 878 3642 881 4028
rect 886 3752 889 4198
rect 926 4162 929 4298
rect 894 4132 897 4138
rect 902 3742 905 4048
rect 910 3902 913 4018
rect 862 3458 870 3461
rect 862 3452 865 3458
rect 826 2888 830 2891
rect 814 2662 817 2738
rect 822 2732 825 2778
rect 838 2682 841 2798
rect 834 2658 838 2661
rect 806 2492 809 2498
rect 806 2462 809 2468
rect 814 2342 817 2658
rect 814 2322 817 2328
rect 758 1868 766 1871
rect 758 1712 761 1748
rect 766 1672 769 1678
rect 766 1541 769 1658
rect 774 1552 777 1838
rect 782 1672 785 1678
rect 766 1538 777 1541
rect 766 1472 769 1478
rect 750 1468 758 1471
rect 742 1132 745 1408
rect 750 1292 753 1318
rect 726 852 729 938
rect 726 772 729 848
rect 742 722 745 1088
rect 750 752 753 1118
rect 750 292 753 748
rect 686 268 694 271
rect 694 142 697 268
rect 694 92 697 138
rect 750 101 753 278
rect 746 98 753 101
rect 758 132 761 618
rect 766 522 769 1128
rect 774 752 777 1538
rect 782 1262 785 1428
rect 782 1152 785 1258
rect 790 1072 793 1538
rect 798 1442 801 2308
rect 806 2112 809 2318
rect 814 2032 817 2198
rect 822 2002 825 2578
rect 846 2552 849 3068
rect 862 2921 865 3368
rect 870 3042 873 3448
rect 870 2942 873 2948
rect 854 2918 865 2921
rect 854 2752 857 2918
rect 846 2532 849 2548
rect 854 2482 857 2708
rect 830 2432 833 2448
rect 830 2132 833 2218
rect 838 2192 841 2458
rect 846 2432 849 2478
rect 806 1918 814 1921
rect 806 1442 809 1918
rect 806 1392 809 1398
rect 798 1328 806 1331
rect 798 1112 801 1328
rect 814 992 817 1698
rect 838 1692 841 2168
rect 846 2162 849 2388
rect 862 2262 865 2468
rect 870 2452 873 2848
rect 878 2341 881 3638
rect 874 2338 881 2341
rect 870 2232 873 2268
rect 858 2188 862 2191
rect 870 2122 873 2228
rect 878 2142 881 2148
rect 822 1442 825 1638
rect 822 1142 825 1438
rect 830 1361 833 1408
rect 846 1362 849 1578
rect 830 1358 838 1361
rect 830 1232 833 1318
rect 838 1232 841 1358
rect 846 1262 849 1358
rect 854 1352 857 1798
rect 862 1332 865 1928
rect 870 1782 873 2108
rect 878 1962 881 1968
rect 834 1148 838 1151
rect 870 1122 873 1778
rect 886 1552 889 3268
rect 894 3122 897 3568
rect 902 3452 905 3738
rect 894 2872 897 3098
rect 902 2882 905 3398
rect 910 3322 913 3878
rect 918 3252 921 4058
rect 926 4042 929 4068
rect 926 3562 929 4038
rect 894 2652 897 2678
rect 894 2392 897 2408
rect 894 2362 897 2388
rect 902 2372 905 2518
rect 894 1962 897 2228
rect 858 1078 862 1081
rect 862 1062 865 1068
rect 782 861 785 868
rect 782 858 790 861
rect 798 852 801 958
rect 814 942 817 978
rect 774 432 777 498
rect 782 472 785 728
rect 758 102 761 128
rect 766 112 769 408
rect 782 352 785 468
rect 790 151 793 668
rect 786 148 793 151
rect 798 142 801 408
rect 806 371 809 918
rect 814 462 817 868
rect 830 812 833 968
rect 822 752 825 758
rect 830 672 833 808
rect 870 642 873 1108
rect 878 722 881 1338
rect 886 1332 889 1348
rect 902 1202 905 2298
rect 910 2232 913 3218
rect 918 2992 921 3228
rect 934 3212 937 4438
rect 942 4062 945 4618
rect 950 3981 953 4568
rect 958 4271 961 4888
rect 1814 4862 1817 4868
rect 1242 4858 1246 4861
rect 1546 4858 1550 4861
rect 990 4572 993 4788
rect 1048 4703 1050 4707
rect 1054 4703 1057 4707
rect 1062 4703 1064 4707
rect 1150 4672 1153 4678
rect 1182 4622 1185 4748
rect 1206 4692 1209 4738
rect 1198 4662 1201 4688
rect 958 4268 966 4271
rect 966 4112 969 4118
rect 962 4068 966 4071
rect 942 3978 953 3981
rect 942 3952 945 3978
rect 942 3292 945 3658
rect 950 3212 953 3968
rect 958 3762 961 3898
rect 958 3422 961 3448
rect 966 3401 969 4038
rect 974 3872 977 4198
rect 982 3462 985 4538
rect 990 3462 993 4438
rect 998 4362 1001 4518
rect 1048 4503 1050 4507
rect 1054 4503 1057 4507
rect 1062 4503 1064 4507
rect 998 4338 1006 4341
rect 998 4332 1001 4338
rect 1006 4252 1009 4268
rect 998 4142 1001 4158
rect 1006 4152 1009 4238
rect 998 3672 1001 3678
rect 1006 3622 1009 4128
rect 1014 3982 1017 4258
rect 1022 4022 1025 4148
rect 1022 3992 1025 4018
rect 994 3458 998 3461
rect 966 3398 974 3401
rect 918 2622 921 2958
rect 918 2492 921 2518
rect 910 2142 913 2148
rect 910 1722 913 2008
rect 898 1148 902 1151
rect 894 1072 897 1138
rect 886 912 889 988
rect 894 912 897 1038
rect 886 842 889 848
rect 902 772 905 1118
rect 910 1032 913 1658
rect 918 1352 921 2418
rect 926 2162 929 3158
rect 934 3032 937 3038
rect 934 2852 937 2878
rect 934 2622 937 2628
rect 942 2382 945 3068
rect 950 3042 953 3148
rect 950 2892 953 3028
rect 958 2912 961 3028
rect 966 2932 969 3328
rect 982 3162 985 3288
rect 990 3272 993 3328
rect 1006 3252 1009 3618
rect 990 3152 993 3158
rect 978 3118 985 3121
rect 982 3112 985 3118
rect 974 2982 977 3048
rect 950 2732 953 2748
rect 958 2362 961 2468
rect 934 2332 937 2348
rect 934 2142 937 2328
rect 942 2252 945 2258
rect 958 2162 961 2228
rect 926 1662 929 1668
rect 934 1492 937 2048
rect 942 1942 945 1958
rect 942 1572 945 1918
rect 950 1692 953 2158
rect 958 2142 961 2148
rect 958 1922 961 2038
rect 966 2012 969 2468
rect 982 2292 985 2928
rect 978 2088 982 2091
rect 982 2022 985 2058
rect 990 2012 993 3138
rect 998 3122 1001 3188
rect 998 2712 1001 3078
rect 1006 2872 1009 3248
rect 1014 3142 1017 3968
rect 1022 3542 1025 3868
rect 1030 3762 1033 4378
rect 1048 4303 1050 4307
rect 1054 4303 1057 4307
rect 1062 4303 1064 4307
rect 1070 4272 1073 4488
rect 1086 4398 1094 4401
rect 1086 4362 1089 4398
rect 1038 4102 1041 4138
rect 1048 4103 1050 4107
rect 1054 4103 1057 4107
rect 1062 4103 1064 4107
rect 1038 3952 1041 3968
rect 1046 3951 1049 4068
rect 1046 3948 1054 3951
rect 1048 3903 1050 3907
rect 1054 3903 1057 3907
rect 1062 3903 1064 3907
rect 1070 3862 1073 4048
rect 1078 3982 1081 4228
rect 1078 3952 1081 3978
rect 1048 3703 1050 3707
rect 1054 3703 1057 3707
rect 1062 3703 1064 3707
rect 1034 3698 1038 3701
rect 1014 2972 1017 2978
rect 1014 2842 1017 2918
rect 1022 2882 1025 3518
rect 1030 3132 1033 3608
rect 1070 3602 1073 3858
rect 1078 3852 1081 3928
rect 1078 3682 1081 3778
rect 1038 3502 1041 3518
rect 1048 3503 1050 3507
rect 1054 3503 1057 3507
rect 1062 3503 1064 3507
rect 1038 3462 1041 3468
rect 1048 3303 1050 3307
rect 1054 3303 1057 3307
rect 1062 3303 1064 3307
rect 1048 3103 1050 3107
rect 1054 3103 1057 3107
rect 1062 3103 1064 3107
rect 1042 2948 1046 2951
rect 1048 2903 1050 2907
rect 1054 2903 1057 2907
rect 1062 2903 1064 2907
rect 1030 2892 1033 2898
rect 1006 2752 1009 2828
rect 998 2652 1001 2678
rect 998 2632 1001 2638
rect 998 2412 1001 2608
rect 1006 2351 1009 2748
rect 1014 2492 1017 2838
rect 1030 2692 1033 2698
rect 998 2348 1009 2351
rect 998 2062 1001 2348
rect 950 1682 953 1688
rect 950 1642 953 1668
rect 950 1542 953 1638
rect 942 1502 945 1518
rect 958 1472 961 1548
rect 918 1092 921 1348
rect 926 1172 929 1468
rect 966 1412 969 1958
rect 974 1922 977 1948
rect 1006 1862 1009 2208
rect 938 1358 942 1361
rect 938 1348 942 1351
rect 930 1058 937 1061
rect 918 812 921 828
rect 934 822 937 1058
rect 910 772 913 778
rect 910 672 913 768
rect 822 482 825 628
rect 870 552 873 588
rect 906 558 910 561
rect 862 542 865 548
rect 854 522 857 538
rect 886 522 889 558
rect 838 518 846 521
rect 838 462 841 518
rect 806 368 814 371
rect 806 242 809 368
rect 838 262 841 458
rect 866 338 870 341
rect 862 292 865 338
rect 918 232 921 788
rect 930 558 934 561
rect 942 561 945 1348
rect 950 802 953 1408
rect 958 1152 961 1158
rect 962 1058 966 1061
rect 974 882 977 1348
rect 982 1262 985 1708
rect 990 1552 993 1858
rect 1006 1842 1009 1858
rect 1014 1592 1017 2478
rect 990 1432 993 1538
rect 990 1102 993 1428
rect 998 1392 1001 1558
rect 1002 1268 1006 1271
rect 998 1132 1001 1138
rect 994 938 998 941
rect 962 858 966 861
rect 966 712 969 728
rect 974 712 977 718
rect 942 558 950 561
rect 926 482 929 548
rect 934 532 937 538
rect 926 472 929 478
rect 958 462 961 468
rect 798 122 801 138
rect 758 82 761 98
rect 918 82 921 228
rect 966 172 969 648
rect 974 372 977 708
rect 982 682 985 878
rect 990 761 993 828
rect 990 758 998 761
rect 998 612 1001 738
rect 1006 462 1009 1258
rect 1014 592 1017 1568
rect 1022 1552 1025 2588
rect 1030 2482 1033 2668
rect 1030 1952 1033 2118
rect 1038 2082 1041 2818
rect 1048 2703 1050 2707
rect 1054 2703 1057 2707
rect 1062 2703 1064 2707
rect 1070 2582 1073 3318
rect 1078 2912 1081 3658
rect 1086 3262 1089 4358
rect 1094 3872 1097 3918
rect 1102 3892 1105 3928
rect 1118 3842 1121 4328
rect 1150 4292 1153 4468
rect 1162 4458 1166 4461
rect 1166 4282 1169 4458
rect 1174 4271 1177 4278
rect 1170 4268 1177 4271
rect 1094 3332 1097 3728
rect 1086 2892 1089 3258
rect 1094 3192 1097 3198
rect 1048 2503 1050 2507
rect 1054 2503 1057 2507
rect 1062 2503 1064 2507
rect 1048 2303 1050 2307
rect 1054 2303 1057 2307
rect 1062 2303 1064 2307
rect 1070 2152 1073 2578
rect 1048 2103 1050 2107
rect 1054 2103 1057 2107
rect 1062 2103 1064 2107
rect 1078 2102 1081 2888
rect 1086 2682 1089 2868
rect 1094 2862 1097 2888
rect 1102 2861 1105 3698
rect 1110 3632 1113 3658
rect 1118 3532 1121 3838
rect 1126 3642 1129 4188
rect 1154 4068 1158 4071
rect 1142 3982 1145 3998
rect 1154 3968 1158 3971
rect 1150 3872 1153 3878
rect 1110 3092 1113 3408
rect 1118 3252 1121 3488
rect 1134 3232 1137 3748
rect 1142 3652 1145 3658
rect 1142 3412 1145 3578
rect 1150 3432 1153 3738
rect 1158 3672 1161 3868
rect 1166 3802 1169 4248
rect 1182 4142 1185 4618
rect 1214 4522 1217 4658
rect 1190 4472 1193 4518
rect 1178 3968 1182 3971
rect 1158 3422 1161 3668
rect 1166 3662 1169 3798
rect 1182 3742 1185 3938
rect 1166 3562 1169 3658
rect 1126 3151 1129 3168
rect 1134 3162 1137 3178
rect 1122 3148 1129 3151
rect 1142 3032 1145 3378
rect 1174 3262 1177 3728
rect 1182 3332 1185 3338
rect 1182 3272 1185 3298
rect 1190 3272 1193 4468
rect 1222 4402 1225 4748
rect 1230 4592 1233 4678
rect 1206 4092 1209 4258
rect 1214 4082 1217 4108
rect 1222 4062 1225 4388
rect 1230 4302 1233 4588
rect 1230 4122 1233 4138
rect 1230 4042 1233 4078
rect 1238 4062 1241 4448
rect 1198 3672 1201 3978
rect 1222 3972 1225 4028
rect 1210 3968 1214 3971
rect 1214 3932 1217 3958
rect 1150 3142 1153 3258
rect 1158 3172 1161 3178
rect 1158 3062 1161 3158
rect 1174 3142 1177 3158
rect 1122 2938 1126 2941
rect 1102 2858 1110 2861
rect 1110 2422 1113 2838
rect 1118 2512 1121 2788
rect 1046 1952 1049 2078
rect 1078 2051 1081 2098
rect 1078 2048 1089 2051
rect 1048 1903 1050 1907
rect 1054 1903 1057 1907
rect 1062 1903 1064 1907
rect 1030 1702 1033 1738
rect 1022 1182 1025 1518
rect 1030 1452 1033 1548
rect 1038 1472 1041 1828
rect 1048 1703 1050 1707
rect 1054 1703 1057 1707
rect 1062 1703 1064 1707
rect 1070 1652 1073 1968
rect 1078 1872 1081 2038
rect 1086 1952 1089 2048
rect 1094 2042 1097 2058
rect 1086 1892 1089 1938
rect 1046 1572 1049 1588
rect 1048 1503 1050 1507
rect 1054 1503 1057 1507
rect 1062 1503 1064 1507
rect 1038 1312 1041 1468
rect 1048 1303 1050 1307
rect 1054 1303 1057 1307
rect 1062 1303 1064 1307
rect 1026 1148 1030 1151
rect 1022 662 1025 1118
rect 1014 552 1017 588
rect 1030 562 1033 1028
rect 1014 402 1017 538
rect 1030 452 1033 538
rect 1038 482 1041 1298
rect 1046 1132 1049 1148
rect 1048 1103 1050 1107
rect 1054 1103 1057 1107
rect 1062 1103 1064 1107
rect 1070 1072 1073 1598
rect 1078 1582 1081 1818
rect 1094 1672 1097 2018
rect 1102 1992 1105 2078
rect 1110 2032 1113 2408
rect 1118 2282 1121 2468
rect 1126 2362 1129 2768
rect 1134 2572 1137 2978
rect 1142 2952 1145 2978
rect 1142 2752 1145 2948
rect 1150 2652 1153 2888
rect 1158 2582 1161 2598
rect 1150 2542 1153 2578
rect 1158 2552 1161 2558
rect 1134 2161 1137 2238
rect 1130 2158 1137 2161
rect 1122 2138 1126 2141
rect 1118 2052 1121 2058
rect 1110 2022 1113 2028
rect 1102 1922 1105 1958
rect 1126 1832 1129 2108
rect 1150 1981 1153 2538
rect 1158 2452 1161 2478
rect 1146 1978 1153 1981
rect 1158 1961 1161 2378
rect 1166 2362 1169 2658
rect 1174 2612 1177 2958
rect 1182 2922 1185 3248
rect 1190 3132 1193 3238
rect 1198 3172 1201 3408
rect 1206 3312 1209 3808
rect 1190 2932 1193 3018
rect 1182 2862 1185 2898
rect 1182 2672 1185 2858
rect 1174 2462 1177 2608
rect 1190 2582 1193 2928
rect 1198 2802 1201 3148
rect 1206 3062 1209 3108
rect 1198 2542 1201 2758
rect 1206 2602 1209 3048
rect 1214 2991 1217 3328
rect 1222 3192 1225 3668
rect 1230 3622 1233 4038
rect 1246 3982 1249 4548
rect 1278 4532 1281 4548
rect 1270 4032 1273 4408
rect 1214 2988 1222 2991
rect 1214 2862 1217 2868
rect 1222 2642 1225 2918
rect 1230 2892 1233 3598
rect 1238 3012 1241 3478
rect 1246 3002 1249 3558
rect 1254 3372 1257 4028
rect 1262 3512 1265 3758
rect 1270 3522 1273 4008
rect 1278 3962 1281 4528
rect 1286 3962 1289 4118
rect 1278 3892 1281 3958
rect 1270 3462 1273 3508
rect 1270 3332 1273 3348
rect 1254 3292 1257 3328
rect 1278 3252 1281 3638
rect 1182 2482 1185 2528
rect 1174 2392 1177 2398
rect 1170 2308 1177 2311
rect 1174 2172 1177 2308
rect 1190 2262 1193 2308
rect 1174 2062 1177 2108
rect 1190 2082 1193 2088
rect 1154 1958 1161 1961
rect 1138 1948 1142 1951
rect 1138 1938 1145 1941
rect 1114 1738 1118 1741
rect 1102 1722 1105 1728
rect 1094 1592 1097 1628
rect 1078 1142 1081 1568
rect 1086 1552 1089 1588
rect 1094 1362 1097 1588
rect 1102 1362 1105 1678
rect 1142 1572 1145 1938
rect 1102 1322 1105 1358
rect 1046 1058 1054 1061
rect 1046 1032 1049 1058
rect 1048 903 1050 907
rect 1054 903 1057 907
rect 1062 903 1064 907
rect 1066 758 1070 761
rect 1050 738 1054 741
rect 1048 703 1050 707
rect 1054 703 1057 707
rect 1062 703 1064 707
rect 1078 692 1081 1078
rect 1086 932 1089 1268
rect 1110 1262 1113 1418
rect 1126 1311 1129 1528
rect 1134 1412 1137 1458
rect 1118 1308 1129 1311
rect 1094 1062 1097 1068
rect 1102 1022 1105 1068
rect 1086 862 1089 918
rect 1086 712 1089 848
rect 1094 732 1097 748
rect 1070 552 1073 568
rect 1070 522 1073 538
rect 1048 503 1050 507
rect 1054 503 1057 507
rect 1062 503 1064 507
rect 1038 472 1041 478
rect 1078 372 1081 688
rect 1102 642 1105 878
rect 1110 742 1113 1238
rect 1118 742 1121 1308
rect 1126 1262 1129 1268
rect 1134 982 1137 1038
rect 1134 732 1137 978
rect 1142 552 1145 1558
rect 1150 1552 1153 1948
rect 1158 1932 1161 1938
rect 1158 1682 1161 1878
rect 1166 1822 1169 2038
rect 1182 2012 1185 2028
rect 1174 1872 1177 1878
rect 1190 1812 1193 2038
rect 1178 1748 1182 1751
rect 1150 1112 1153 1548
rect 1158 922 1161 1548
rect 1166 1512 1169 1618
rect 1174 1572 1177 1648
rect 1166 1442 1169 1508
rect 1166 1141 1169 1318
rect 1174 1162 1177 1468
rect 1182 1202 1185 1698
rect 1190 1462 1193 1778
rect 1198 1692 1201 2258
rect 1206 2032 1209 2548
rect 1214 2442 1217 2618
rect 1238 2552 1241 2928
rect 1270 2842 1273 2858
rect 1246 2662 1249 2668
rect 1230 2542 1233 2548
rect 1230 2528 1238 2531
rect 1230 2512 1233 2528
rect 1230 2472 1233 2488
rect 1230 2422 1233 2468
rect 1214 2282 1217 2418
rect 1222 2352 1225 2358
rect 1230 2352 1233 2358
rect 1214 2261 1217 2278
rect 1214 2258 1222 2261
rect 1214 1842 1217 1898
rect 1210 1748 1214 1751
rect 1198 1532 1201 1578
rect 1198 1462 1201 1468
rect 1166 1138 1174 1141
rect 1174 942 1177 1098
rect 1174 742 1177 938
rect 1182 802 1185 968
rect 1174 672 1177 738
rect 1134 472 1137 518
rect 1174 402 1177 668
rect 1190 572 1193 1438
rect 1198 1432 1201 1438
rect 1198 1342 1201 1368
rect 1198 1272 1201 1288
rect 1198 1252 1201 1258
rect 1198 912 1201 1208
rect 1206 892 1209 1678
rect 1214 1542 1217 1548
rect 1222 1482 1225 1908
rect 1230 1872 1233 1878
rect 1238 1802 1241 2438
rect 1246 2362 1249 2558
rect 1254 2462 1257 2628
rect 1262 2452 1265 2488
rect 1258 2438 1262 2441
rect 1254 2292 1257 2408
rect 1262 2352 1265 2368
rect 1254 2272 1257 2278
rect 1246 2202 1249 2268
rect 1230 1672 1233 1718
rect 1230 1432 1233 1448
rect 1218 1428 1222 1431
rect 1238 1402 1241 1708
rect 1246 1652 1249 1658
rect 1214 1262 1217 1388
rect 1230 1351 1233 1358
rect 1226 1348 1233 1351
rect 1238 1312 1241 1328
rect 1246 1322 1249 1648
rect 1254 1332 1257 1778
rect 1262 1632 1265 2308
rect 1270 2132 1273 2498
rect 1278 2442 1281 3108
rect 1286 2912 1289 3768
rect 1294 3342 1297 4108
rect 1302 3582 1305 4828
rect 1354 4748 1358 4751
rect 1310 4642 1313 4658
rect 1318 4642 1321 4698
rect 1310 4632 1313 4638
rect 1310 4142 1313 4478
rect 1326 4282 1329 4718
rect 1334 4672 1337 4678
rect 1386 4658 1390 4661
rect 1382 4552 1385 4598
rect 1382 4542 1385 4548
rect 1310 4042 1313 4128
rect 1334 3912 1337 4468
rect 1342 3962 1345 4078
rect 1310 3738 1318 3741
rect 1310 3712 1313 3738
rect 1310 3682 1313 3708
rect 1310 3601 1313 3608
rect 1310 3598 1318 3601
rect 1302 3462 1305 3538
rect 1310 3522 1313 3568
rect 1318 3552 1321 3558
rect 1294 3142 1297 3308
rect 1294 3062 1297 3138
rect 1294 2662 1297 3038
rect 1310 2962 1313 3488
rect 1318 3112 1321 3548
rect 1326 3482 1329 3538
rect 1334 3512 1337 3848
rect 1326 3222 1329 3448
rect 1334 3432 1337 3468
rect 1350 3451 1353 3778
rect 1358 3682 1361 4148
rect 1366 3742 1369 4118
rect 1374 4092 1377 4168
rect 1358 3471 1361 3678
rect 1358 3468 1366 3471
rect 1350 3448 1361 3451
rect 1350 3312 1353 3438
rect 1358 3432 1361 3448
rect 1374 3422 1377 3928
rect 1382 3572 1385 4538
rect 1422 4472 1425 4818
rect 1560 4803 1562 4807
rect 1566 4803 1569 4807
rect 1574 4803 1576 4807
rect 1506 4748 1510 4751
rect 1634 4748 1638 4751
rect 1622 4742 1625 4748
rect 1542 4652 1545 4708
rect 1446 4532 1449 4548
rect 1494 4542 1497 4548
rect 1446 4352 1449 4528
rect 1502 4461 1505 4618
rect 1502 4458 1510 4461
rect 1454 4422 1457 4458
rect 1462 4302 1465 4338
rect 1494 4322 1497 4458
rect 1406 4152 1409 4208
rect 1398 4092 1401 4148
rect 1390 3552 1393 3738
rect 1398 3712 1401 4088
rect 1414 4062 1417 4228
rect 1410 4058 1414 4061
rect 1318 2962 1321 2968
rect 1302 2942 1305 2948
rect 1314 2938 1318 2941
rect 1278 2372 1281 2378
rect 1286 2152 1289 2568
rect 1294 2342 1297 2658
rect 1302 2281 1305 2678
rect 1294 2278 1305 2281
rect 1286 2072 1289 2148
rect 1270 2032 1273 2068
rect 1270 1702 1273 2018
rect 1278 1972 1281 2038
rect 1294 2031 1297 2278
rect 1302 2072 1305 2268
rect 1294 2028 1305 2031
rect 1226 1308 1230 1311
rect 1194 528 1198 531
rect 1190 492 1193 528
rect 1214 472 1217 1148
rect 1222 682 1225 1288
rect 1262 1242 1265 1368
rect 1238 1142 1241 1148
rect 1230 512 1233 898
rect 1238 822 1241 858
rect 1238 792 1241 818
rect 1246 652 1249 1018
rect 1254 752 1257 878
rect 1086 332 1089 388
rect 1230 371 1233 398
rect 1226 368 1233 371
rect 1246 371 1249 648
rect 1242 368 1249 371
rect 1254 542 1257 748
rect 1270 552 1273 1648
rect 1278 912 1281 1738
rect 1286 1672 1289 1968
rect 1302 1962 1305 2028
rect 1302 1862 1305 1958
rect 1310 1952 1313 2888
rect 1318 2572 1321 2888
rect 1326 2872 1329 3128
rect 1334 2992 1337 3148
rect 1342 3021 1345 3268
rect 1362 3228 1369 3231
rect 1366 3112 1369 3228
rect 1374 3122 1377 3418
rect 1382 3262 1385 3478
rect 1390 3452 1393 3458
rect 1398 3442 1401 3698
rect 1406 3472 1409 3628
rect 1414 3522 1417 3868
rect 1430 3832 1433 4218
rect 1526 4162 1529 4588
rect 1534 4532 1537 4548
rect 1542 4272 1545 4648
rect 1560 4603 1562 4607
rect 1566 4603 1569 4607
rect 1574 4603 1576 4607
rect 1574 4522 1577 4528
rect 1558 4422 1561 4438
rect 1560 4403 1562 4407
rect 1566 4403 1569 4407
rect 1574 4403 1576 4407
rect 1582 4362 1585 4608
rect 1590 4462 1593 4648
rect 1606 4532 1609 4648
rect 1598 4452 1601 4468
rect 1494 4142 1497 4158
rect 1486 3942 1489 4078
rect 1446 3912 1449 3938
rect 1446 3872 1449 3908
rect 1442 3718 1446 3721
rect 1462 3671 1465 3928
rect 1478 3862 1481 3898
rect 1462 3668 1470 3671
rect 1422 3552 1425 3568
rect 1434 3518 1438 3521
rect 1450 3498 1454 3501
rect 1414 3482 1417 3498
rect 1358 3052 1361 3068
rect 1350 3032 1353 3048
rect 1342 3018 1353 3021
rect 1334 2951 1337 2988
rect 1334 2948 1342 2951
rect 1318 2532 1321 2538
rect 1326 2472 1329 2868
rect 1334 2832 1337 2948
rect 1350 2942 1353 3018
rect 1342 2772 1345 2838
rect 1350 2712 1353 2938
rect 1358 2832 1361 3028
rect 1374 2982 1377 3068
rect 1366 2672 1369 2678
rect 1318 2461 1321 2468
rect 1318 2458 1329 2461
rect 1318 2392 1321 2418
rect 1318 2382 1321 2388
rect 1318 2142 1321 2158
rect 1326 2112 1329 2458
rect 1350 2382 1353 2438
rect 1334 2222 1337 2278
rect 1342 2201 1345 2348
rect 1334 2198 1345 2201
rect 1350 2242 1353 2298
rect 1334 2112 1337 2198
rect 1298 1788 1302 1791
rect 1294 1212 1297 1778
rect 1302 1522 1305 1708
rect 1302 1052 1305 1488
rect 1310 1222 1313 1928
rect 1318 1792 1321 1838
rect 1326 1832 1329 2108
rect 1338 2088 1345 2091
rect 1342 2072 1345 2088
rect 1342 1952 1345 1988
rect 1350 1972 1353 2238
rect 1358 2192 1361 2458
rect 1366 2372 1369 2638
rect 1374 2512 1377 2898
rect 1382 2662 1385 3168
rect 1390 2982 1393 3398
rect 1398 3032 1401 3358
rect 1406 3332 1409 3358
rect 1414 3122 1417 3478
rect 1470 3472 1473 3668
rect 1422 3332 1425 3348
rect 1430 3312 1433 3468
rect 1414 3062 1417 3118
rect 1374 2432 1377 2498
rect 1390 2462 1393 2968
rect 1398 2682 1401 2978
rect 1422 2792 1425 2988
rect 1398 2552 1401 2668
rect 1406 2562 1409 2738
rect 1422 2732 1425 2758
rect 1430 2722 1433 2978
rect 1438 2952 1441 3128
rect 1446 3012 1449 3448
rect 1454 3222 1457 3458
rect 1462 3332 1465 3338
rect 1470 3322 1473 3378
rect 1454 3072 1457 3218
rect 1438 2942 1441 2948
rect 1462 2922 1465 3188
rect 1470 3142 1473 3248
rect 1478 3232 1481 3858
rect 1486 3652 1489 3788
rect 1486 3532 1489 3598
rect 1494 3542 1497 4138
rect 1510 4131 1513 4138
rect 1510 4128 1518 4131
rect 1494 3532 1497 3538
rect 1502 3452 1505 3978
rect 1510 3722 1513 4128
rect 1526 4042 1529 4058
rect 1534 4052 1537 4068
rect 1518 3462 1521 3968
rect 1486 3402 1489 3438
rect 1490 3358 1494 3361
rect 1502 3302 1505 3338
rect 1502 3292 1505 3298
rect 1510 3272 1513 3418
rect 1494 3202 1497 3248
rect 1494 3152 1497 3168
rect 1502 3162 1505 3228
rect 1486 3082 1489 3138
rect 1438 2802 1441 2808
rect 1414 2682 1417 2688
rect 1414 2592 1417 2648
rect 1422 2552 1425 2708
rect 1446 2682 1449 2908
rect 1454 2762 1457 2808
rect 1430 2602 1433 2658
rect 1462 2652 1465 2838
rect 1470 2552 1473 3058
rect 1478 2802 1481 3048
rect 1398 2512 1401 2548
rect 1358 1961 1361 2188
rect 1366 2152 1369 2368
rect 1354 1958 1361 1961
rect 1318 1592 1321 1788
rect 1326 1652 1329 1698
rect 1322 1558 1326 1561
rect 1286 782 1289 1038
rect 1318 982 1321 1518
rect 1326 1452 1329 1458
rect 1334 1342 1337 1948
rect 1342 1512 1345 1938
rect 1366 1782 1369 2138
rect 1374 1882 1377 2418
rect 1354 1768 1358 1771
rect 1342 1461 1345 1468
rect 1342 1458 1350 1461
rect 1326 1262 1329 1268
rect 1334 1192 1337 1308
rect 1342 1152 1345 1318
rect 1350 1312 1353 1358
rect 1358 1262 1361 1488
rect 1366 1432 1369 1658
rect 1374 1582 1377 1718
rect 1370 1358 1374 1361
rect 1342 722 1345 908
rect 1254 402 1257 538
rect 1278 472 1281 708
rect 1342 702 1345 718
rect 1110 338 1118 341
rect 1048 303 1050 307
rect 1054 303 1057 307
rect 1062 303 1064 307
rect 1078 272 1081 278
rect 1058 238 1062 241
rect 1110 202 1113 338
rect 1254 142 1257 398
rect 1270 312 1273 378
rect 1286 371 1289 678
rect 1286 368 1294 371
rect 1302 302 1305 528
rect 1330 368 1334 371
rect 1350 342 1353 938
rect 1270 272 1273 288
rect 1302 262 1305 298
rect 1310 232 1313 278
rect 1350 272 1353 338
rect 1358 282 1361 738
rect 1366 622 1369 1338
rect 1382 1302 1385 2328
rect 1390 2162 1393 2428
rect 1390 1552 1393 2148
rect 1398 2122 1401 2468
rect 1406 2322 1409 2328
rect 1406 2302 1409 2308
rect 1414 2162 1417 2408
rect 1398 1882 1401 2108
rect 1390 1502 1393 1508
rect 1390 1372 1393 1378
rect 1398 1352 1401 1868
rect 1406 1582 1409 2148
rect 1422 1932 1425 2548
rect 1446 2542 1449 2548
rect 1430 2412 1433 2538
rect 1430 2172 1433 2388
rect 1430 2052 1433 2158
rect 1414 1822 1417 1918
rect 1430 1802 1433 2048
rect 1406 1548 1414 1551
rect 1406 1362 1409 1548
rect 1422 1532 1425 1598
rect 1422 1472 1425 1488
rect 1382 1272 1385 1298
rect 1390 952 1393 1348
rect 1398 1272 1401 1348
rect 1406 1252 1409 1258
rect 1398 1238 1406 1241
rect 1398 1092 1401 1238
rect 1414 972 1417 1158
rect 1422 992 1425 1408
rect 1390 712 1393 898
rect 1430 861 1433 1748
rect 1446 1662 1449 2538
rect 1454 2442 1457 2448
rect 1462 2362 1465 2458
rect 1454 1752 1457 2078
rect 1462 1682 1465 2248
rect 1470 2142 1473 2548
rect 1470 2092 1473 2118
rect 1426 858 1433 861
rect 1414 812 1417 828
rect 1422 772 1425 778
rect 1430 772 1433 838
rect 1438 822 1441 1638
rect 1470 1542 1473 1868
rect 1478 1822 1481 2638
rect 1486 2632 1489 3018
rect 1494 2822 1497 2868
rect 1486 2552 1489 2568
rect 1494 2542 1497 2768
rect 1502 2732 1505 2998
rect 1518 2982 1521 3418
rect 1526 3271 1529 3858
rect 1534 3691 1537 3808
rect 1542 3722 1545 4038
rect 1550 3972 1553 4328
rect 1560 4203 1562 4207
rect 1566 4203 1569 4207
rect 1574 4203 1576 4207
rect 1560 4003 1562 4007
rect 1566 4003 1569 4007
rect 1574 4003 1576 4007
rect 1534 3688 1545 3691
rect 1534 3672 1537 3678
rect 1534 3282 1537 3468
rect 1526 3268 1537 3271
rect 1510 2932 1513 2958
rect 1510 2842 1513 2868
rect 1502 2652 1505 2678
rect 1510 2662 1513 2668
rect 1510 2552 1513 2648
rect 1502 2342 1505 2378
rect 1486 2312 1489 2338
rect 1486 2042 1489 2068
rect 1486 1992 1489 2038
rect 1494 2002 1497 2318
rect 1510 2282 1513 2348
rect 1502 2202 1505 2258
rect 1502 2072 1505 2078
rect 1502 1962 1505 1968
rect 1502 1938 1510 1941
rect 1478 1802 1481 1818
rect 1478 1742 1481 1748
rect 1478 1712 1481 1718
rect 1486 1662 1489 1818
rect 1494 1752 1497 1798
rect 1502 1742 1505 1938
rect 1518 1872 1521 2918
rect 1526 2902 1529 3138
rect 1534 3052 1537 3268
rect 1534 2992 1537 3048
rect 1534 2872 1537 2978
rect 1542 2912 1545 3688
rect 1550 3162 1553 3858
rect 1558 3852 1561 3938
rect 1570 3868 1574 3871
rect 1590 3862 1593 4418
rect 1598 3911 1601 4368
rect 1614 4242 1617 4538
rect 1622 4522 1625 4658
rect 1634 4538 1638 4541
rect 1622 4292 1625 4458
rect 1630 4201 1633 4508
rect 1630 4198 1638 4201
rect 1598 3908 1606 3911
rect 1560 3803 1562 3807
rect 1566 3803 1569 3807
rect 1574 3803 1576 3807
rect 1582 3692 1585 3808
rect 1590 3692 1593 3708
rect 1582 3652 1585 3678
rect 1598 3672 1601 3688
rect 1614 3672 1617 4058
rect 1622 4022 1625 4048
rect 1560 3603 1562 3607
rect 1566 3603 1569 3607
rect 1574 3603 1576 3607
rect 1582 3602 1585 3648
rect 1590 3622 1593 3648
rect 1560 3403 1562 3407
rect 1566 3403 1569 3407
rect 1574 3403 1576 3407
rect 1560 3203 1562 3207
rect 1566 3203 1569 3207
rect 1574 3203 1576 3207
rect 1582 3202 1585 3368
rect 1590 3272 1593 3528
rect 1598 3482 1601 3508
rect 1550 3152 1553 3158
rect 1606 3142 1609 3588
rect 1630 3582 1633 4048
rect 1638 3562 1641 4138
rect 1626 3548 1630 3551
rect 1630 3462 1633 3468
rect 1582 3012 1585 3048
rect 1560 3003 1562 3007
rect 1566 3003 1569 3007
rect 1574 3003 1576 3007
rect 1582 2892 1585 2998
rect 1542 2752 1545 2868
rect 1550 2812 1553 2828
rect 1560 2803 1562 2807
rect 1566 2803 1569 2807
rect 1574 2803 1576 2807
rect 1582 2802 1585 2878
rect 1570 2618 1574 2621
rect 1526 2562 1529 2588
rect 1542 2572 1545 2598
rect 1526 2312 1529 2538
rect 1534 2272 1537 2288
rect 1542 2221 1545 2488
rect 1534 2218 1545 2221
rect 1534 1972 1537 2218
rect 1530 1908 1534 1911
rect 1510 1792 1513 1828
rect 1494 1728 1502 1731
rect 1486 1552 1489 1658
rect 1494 1552 1497 1728
rect 1518 1642 1521 1848
rect 1526 1762 1529 1808
rect 1534 1532 1537 1818
rect 1542 1782 1545 2208
rect 1550 2062 1553 2608
rect 1560 2603 1562 2607
rect 1566 2603 1569 2607
rect 1574 2603 1576 2607
rect 1558 2442 1561 2488
rect 1582 2462 1585 2698
rect 1590 2612 1593 2848
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1574 2403 1576 2407
rect 1582 2301 1585 2448
rect 1590 2311 1593 2528
rect 1598 2371 1601 3098
rect 1606 2852 1609 3078
rect 1622 3072 1625 3458
rect 1630 3272 1633 3308
rect 1638 3282 1641 3558
rect 1614 3052 1617 3068
rect 1630 2952 1633 3268
rect 1622 2881 1625 2898
rect 1630 2892 1633 2948
rect 1622 2878 1630 2881
rect 1606 2842 1609 2848
rect 1630 2842 1633 2868
rect 1622 2742 1625 2758
rect 1606 2442 1609 2618
rect 1606 2392 1609 2408
rect 1598 2368 1606 2371
rect 1590 2308 1598 2311
rect 1582 2298 1593 2301
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1574 2203 1576 2207
rect 1582 2202 1585 2218
rect 1558 2122 1561 2128
rect 1582 2072 1585 2078
rect 1550 2012 1553 2038
rect 1566 2032 1569 2058
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1574 2003 1576 2007
rect 1542 1582 1545 1678
rect 1502 1492 1505 1528
rect 1482 1488 1486 1491
rect 1506 1488 1510 1491
rect 1446 1252 1449 1398
rect 1458 1278 1462 1281
rect 1446 1162 1449 1248
rect 1450 1068 1454 1071
rect 1462 962 1465 1218
rect 1398 462 1401 728
rect 1398 392 1401 458
rect 1406 272 1409 728
rect 1414 681 1417 768
rect 1414 678 1422 681
rect 1418 658 1425 661
rect 1422 432 1425 658
rect 1446 542 1449 698
rect 1422 362 1425 368
rect 1048 103 1050 107
rect 1054 103 1057 107
rect 1062 103 1064 107
rect 978 68 982 71
rect 350 62 353 68
rect 1310 62 1313 228
rect 1430 142 1433 408
rect 1438 352 1441 488
rect 1446 322 1449 538
rect 1454 432 1457 658
rect 1470 482 1473 1438
rect 1478 1152 1481 1488
rect 1494 1152 1497 1338
rect 1494 1082 1497 1148
rect 1502 952 1505 1358
rect 1518 1162 1521 1528
rect 1550 1492 1553 1978
rect 1590 1882 1593 2298
rect 1614 2292 1617 2458
rect 1618 2268 1622 2271
rect 1606 2242 1609 2258
rect 1630 2112 1633 2628
rect 1638 2321 1641 3178
rect 1646 2882 1649 3658
rect 1654 3422 1657 4028
rect 1662 3212 1665 3928
rect 1670 3752 1673 4808
rect 1678 4748 1686 4751
rect 1678 4732 1681 4748
rect 1702 4742 1705 4748
rect 1714 4528 1718 4531
rect 1678 3742 1681 4318
rect 1670 3732 1673 3738
rect 1686 3731 1689 4228
rect 1694 4062 1697 4318
rect 1726 4272 1729 4548
rect 1750 4292 1753 4808
rect 1766 4732 1769 4808
rect 1814 4752 1817 4858
rect 1766 4672 1769 4728
rect 1814 4562 1817 4748
rect 1710 4132 1713 4148
rect 1718 4142 1721 4148
rect 1702 3912 1705 4108
rect 1678 3728 1689 3731
rect 1670 3602 1673 3718
rect 1670 3262 1673 3598
rect 1678 3562 1681 3728
rect 1694 3722 1697 3748
rect 1686 3512 1689 3718
rect 1678 3452 1681 3468
rect 1654 2702 1657 3108
rect 1662 3032 1665 3088
rect 1670 3062 1673 3258
rect 1678 3162 1681 3378
rect 1686 3302 1689 3508
rect 1694 3462 1697 3678
rect 1702 3632 1705 3908
rect 1710 3772 1713 4128
rect 1718 3812 1721 4128
rect 1726 4082 1729 4268
rect 1734 4152 1737 4258
rect 1750 4182 1753 4208
rect 1726 4072 1729 4078
rect 1694 3292 1697 3458
rect 1702 3442 1705 3628
rect 1710 3562 1713 3738
rect 1718 3692 1721 3698
rect 1718 3462 1721 3678
rect 1710 3342 1713 3378
rect 1718 3342 1721 3358
rect 1706 3338 1710 3341
rect 1710 3208 1718 3211
rect 1670 2891 1673 2958
rect 1666 2888 1673 2891
rect 1662 2852 1665 2878
rect 1678 2872 1681 3088
rect 1650 2668 1654 2671
rect 1646 2422 1649 2588
rect 1662 2542 1665 2628
rect 1670 2562 1673 2858
rect 1678 2812 1681 2828
rect 1654 2482 1657 2518
rect 1654 2372 1657 2398
rect 1670 2392 1673 2548
rect 1638 2318 1649 2321
rect 1638 2182 1641 2308
rect 1634 2078 1638 2081
rect 1606 1992 1609 2008
rect 1606 1922 1609 1938
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1574 1803 1576 1807
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1574 1603 1576 1607
rect 1570 1558 1574 1561
rect 1558 1552 1561 1558
rect 1566 1532 1569 1548
rect 1550 1452 1553 1488
rect 1566 1452 1569 1528
rect 1526 1172 1529 1448
rect 1542 1322 1545 1348
rect 1550 1302 1553 1428
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1574 1403 1576 1407
rect 1558 1342 1561 1348
rect 1582 1282 1585 1878
rect 1590 1552 1593 1598
rect 1598 1552 1601 1558
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1574 1203 1576 1207
rect 1558 1122 1561 1148
rect 1482 948 1486 951
rect 1526 942 1529 1038
rect 1478 928 1486 931
rect 1478 792 1481 928
rect 1526 892 1529 898
rect 1542 812 1545 1058
rect 1558 1052 1561 1118
rect 1582 1012 1585 1278
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1574 1003 1576 1007
rect 1550 852 1553 958
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1574 803 1576 807
rect 1478 742 1481 788
rect 1590 762 1593 1318
rect 1598 1292 1601 1478
rect 1606 1362 1609 1868
rect 1614 1431 1617 2058
rect 1622 1442 1625 1918
rect 1630 1442 1633 2038
rect 1646 1941 1649 2318
rect 1654 2222 1657 2288
rect 1662 2162 1665 2308
rect 1678 2282 1681 2758
rect 1686 2552 1689 3128
rect 1710 3122 1713 3208
rect 1726 3162 1729 3988
rect 1742 3942 1745 3958
rect 1734 3682 1737 3718
rect 1734 3352 1737 3448
rect 1698 3078 1702 3081
rect 1698 3048 1702 3051
rect 1694 2952 1697 3028
rect 1694 2782 1697 2888
rect 1702 2792 1705 2938
rect 1702 2742 1705 2788
rect 1710 2722 1713 3118
rect 1718 2742 1721 2908
rect 1726 2782 1729 3138
rect 1734 3052 1737 3348
rect 1742 3122 1745 3878
rect 1750 3722 1753 4118
rect 1758 3772 1761 4498
rect 1766 4062 1769 4488
rect 1774 3962 1777 4508
rect 1886 4482 1889 4818
rect 1846 4468 1854 4471
rect 1750 3662 1753 3678
rect 1750 3622 1753 3658
rect 1750 3582 1753 3598
rect 1758 3592 1761 3688
rect 1766 3662 1769 3918
rect 1782 3862 1785 4278
rect 1806 4092 1809 4378
rect 1806 3962 1809 4018
rect 1814 3942 1817 4248
rect 1758 3552 1761 3558
rect 1758 3222 1761 3548
rect 1694 2562 1697 2638
rect 1718 2612 1721 2738
rect 1710 2582 1713 2598
rect 1726 2512 1729 2748
rect 1686 2422 1689 2508
rect 1734 2442 1737 3038
rect 1742 2492 1745 3108
rect 1750 2942 1753 3188
rect 1758 3042 1761 3218
rect 1758 2852 1761 2988
rect 1750 2752 1753 2848
rect 1750 2732 1753 2738
rect 1750 2632 1753 2678
rect 1750 2512 1753 2518
rect 1670 2272 1673 2278
rect 1662 2142 1665 2158
rect 1670 2108 1678 2111
rect 1638 1938 1649 1941
rect 1614 1428 1625 1431
rect 1598 1261 1601 1288
rect 1598 1258 1606 1261
rect 1614 1142 1617 1338
rect 1622 1202 1625 1428
rect 1638 1412 1641 1938
rect 1646 1722 1649 1928
rect 1638 1382 1641 1398
rect 1646 1392 1649 1468
rect 1598 982 1601 1028
rect 1614 982 1617 1058
rect 1598 852 1601 978
rect 1606 852 1609 978
rect 1638 882 1641 1258
rect 1646 1082 1649 1358
rect 1654 1102 1657 1858
rect 1662 1702 1665 2088
rect 1662 1262 1665 1638
rect 1670 1622 1673 2108
rect 1686 2062 1689 2408
rect 1694 2272 1697 2328
rect 1702 2242 1705 2438
rect 1714 2348 1718 2351
rect 1718 2152 1721 2208
rect 1694 2072 1697 2108
rect 1702 2102 1705 2108
rect 1682 2018 1686 2021
rect 1702 1602 1705 1998
rect 1710 1992 1713 2038
rect 1702 1552 1705 1578
rect 1694 1548 1702 1551
rect 1678 1492 1681 1498
rect 1686 1471 1689 1498
rect 1682 1468 1689 1471
rect 1654 1002 1657 1058
rect 1662 952 1665 968
rect 1678 932 1681 1138
rect 1606 802 1609 848
rect 1630 842 1633 858
rect 1642 848 1646 851
rect 1454 172 1457 428
rect 1450 148 1454 151
rect 1462 142 1465 388
rect 1470 282 1473 318
rect 1462 62 1465 138
rect 1470 112 1473 278
rect 1486 242 1489 558
rect 1494 492 1497 718
rect 1518 622 1521 638
rect 1518 471 1521 618
rect 1514 468 1521 471
rect 1518 442 1521 448
rect 1534 362 1537 728
rect 1622 712 1625 818
rect 1638 762 1641 848
rect 1686 822 1689 1468
rect 1630 698 1638 701
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1574 603 1576 607
rect 1542 551 1545 568
rect 1622 552 1625 698
rect 1630 652 1633 698
rect 1542 548 1550 551
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1574 403 1576 407
rect 1502 272 1505 348
rect 1534 292 1537 358
rect 1526 272 1529 278
rect 1502 212 1505 268
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1574 203 1576 207
rect 1582 192 1585 218
rect 1490 148 1494 151
rect 1558 62 1561 148
rect 1590 142 1593 268
rect 1622 262 1625 548
rect 1662 202 1665 778
rect 1674 748 1678 751
rect 1686 672 1689 788
rect 1694 752 1697 1548
rect 1710 1532 1713 1778
rect 1718 1532 1721 2128
rect 1726 2122 1729 2268
rect 1734 2262 1737 2388
rect 1742 2181 1745 2488
rect 1750 2432 1753 2468
rect 1750 2392 1753 2398
rect 1750 2322 1753 2348
rect 1734 2178 1745 2181
rect 1750 2242 1753 2268
rect 1726 1652 1729 2108
rect 1734 1902 1737 2178
rect 1742 2052 1745 2128
rect 1750 2122 1753 2238
rect 1758 2042 1761 2848
rect 1766 2452 1769 3658
rect 1774 3522 1777 3528
rect 1782 3422 1785 3778
rect 1790 3662 1793 3908
rect 1774 2862 1777 3248
rect 1782 3082 1785 3408
rect 1798 3172 1801 3898
rect 1814 3832 1817 3838
rect 1806 3312 1809 3748
rect 1814 3652 1817 3658
rect 1798 3112 1801 3168
rect 1782 2902 1785 3048
rect 1790 3042 1793 3108
rect 1806 2962 1809 3208
rect 1814 3012 1817 3498
rect 1822 3292 1825 4258
rect 1838 4252 1841 4418
rect 1846 4392 1849 4468
rect 1854 4372 1857 4458
rect 1894 4452 1897 4678
rect 1902 4372 1905 4718
rect 2030 4662 2033 4728
rect 2072 4703 2074 4707
rect 2078 4703 2081 4707
rect 2086 4703 2088 4707
rect 1830 3502 1833 4058
rect 1838 3952 1841 3998
rect 1854 3792 1857 4368
rect 1910 4312 1913 4528
rect 1918 4472 1921 4478
rect 1926 4382 1929 4518
rect 1958 4442 1961 4648
rect 1862 3962 1865 4158
rect 1862 3822 1865 3888
rect 1870 3882 1873 4198
rect 1910 4182 1913 4188
rect 1902 4062 1905 4068
rect 1894 4032 1897 4058
rect 1934 4052 1937 4068
rect 1886 3871 1889 4028
rect 1882 3868 1889 3871
rect 1842 3588 1849 3591
rect 1782 2802 1785 2898
rect 1806 2792 1809 2808
rect 1774 2742 1777 2768
rect 1774 2132 1777 2728
rect 1782 2492 1785 2778
rect 1798 2662 1801 2748
rect 1798 2542 1801 2608
rect 1806 2482 1809 2488
rect 1742 1982 1745 2038
rect 1734 1832 1737 1888
rect 1758 1842 1761 2038
rect 1766 1942 1769 2058
rect 1774 1942 1777 1948
rect 1766 1832 1769 1938
rect 1774 1862 1777 1878
rect 1734 1612 1737 1758
rect 1750 1742 1753 1778
rect 1742 1698 1750 1701
rect 1702 1152 1705 1478
rect 1710 1292 1713 1368
rect 1706 1148 1710 1151
rect 1718 1142 1721 1528
rect 1702 872 1705 1118
rect 1710 1072 1713 1108
rect 1674 658 1678 661
rect 1678 92 1681 598
rect 1686 552 1689 668
rect 1702 552 1705 858
rect 1710 692 1713 1068
rect 1726 922 1729 1598
rect 1734 1222 1737 1548
rect 1742 1432 1745 1698
rect 1750 1642 1753 1668
rect 1758 1452 1761 1758
rect 1774 1712 1777 1848
rect 1782 1762 1785 2428
rect 1790 2402 1793 2458
rect 1806 2402 1809 2448
rect 1790 2172 1793 2268
rect 1790 2152 1793 2158
rect 1798 2142 1801 2338
rect 1774 1592 1777 1668
rect 1766 1512 1769 1538
rect 1782 1522 1785 1558
rect 1742 1312 1745 1398
rect 1694 372 1697 458
rect 1694 361 1697 368
rect 1694 358 1702 361
rect 1718 292 1721 868
rect 1726 832 1729 858
rect 1726 548 1734 551
rect 1726 462 1729 548
rect 1726 322 1729 458
rect 1734 372 1737 488
rect 1750 382 1753 1428
rect 1766 1352 1769 1508
rect 1790 1471 1793 1708
rect 1798 1702 1801 2008
rect 1806 1892 1809 2298
rect 1814 2252 1817 2928
rect 1822 2682 1825 3278
rect 1830 2892 1833 3128
rect 1830 2752 1833 2878
rect 1838 2692 1841 3458
rect 1846 3092 1849 3588
rect 1854 3362 1857 3748
rect 1862 3532 1865 3798
rect 1894 3792 1897 3878
rect 1910 3762 1913 4028
rect 1930 3988 1937 3991
rect 1910 3702 1913 3758
rect 1862 3432 1865 3448
rect 1830 2552 1833 2578
rect 1838 2571 1841 2678
rect 1846 2592 1849 3088
rect 1854 2871 1857 3158
rect 1870 3071 1873 3278
rect 1878 3081 1881 3688
rect 1878 3078 1889 3081
rect 1870 3068 1881 3071
rect 1854 2868 1862 2871
rect 1854 2772 1857 2818
rect 1846 2582 1849 2588
rect 1838 2568 1849 2571
rect 1822 2532 1825 2548
rect 1838 2542 1841 2558
rect 1834 2478 1838 2481
rect 1822 2322 1825 2328
rect 1830 2311 1833 2448
rect 1846 2432 1849 2568
rect 1854 2552 1857 2678
rect 1862 2602 1865 2748
rect 1870 2662 1873 2988
rect 1878 2932 1881 3068
rect 1878 2732 1881 2828
rect 1870 2471 1873 2618
rect 1862 2468 1873 2471
rect 1838 2412 1841 2428
rect 1838 2332 1841 2348
rect 1822 2308 1833 2311
rect 1822 2222 1825 2308
rect 1830 2222 1833 2228
rect 1838 2222 1841 2318
rect 1846 2301 1849 2338
rect 1846 2298 1854 2301
rect 1814 2122 1817 2198
rect 1838 2182 1841 2208
rect 1822 1942 1825 2178
rect 1830 1952 1833 2048
rect 1838 1902 1841 1958
rect 1846 1872 1849 2078
rect 1806 1852 1809 1868
rect 1854 1862 1857 2028
rect 1838 1858 1846 1861
rect 1806 1622 1809 1848
rect 1814 1662 1817 1718
rect 1822 1622 1825 1658
rect 1790 1468 1798 1471
rect 1766 1232 1769 1348
rect 1758 702 1761 1108
rect 1766 852 1769 1228
rect 1774 1072 1777 1458
rect 1774 952 1777 978
rect 1774 692 1777 908
rect 1758 652 1761 658
rect 1758 382 1761 518
rect 1766 472 1769 668
rect 1782 482 1785 1448
rect 1798 1132 1801 1408
rect 1798 872 1801 1128
rect 1806 1042 1809 1108
rect 1806 512 1809 988
rect 1814 742 1817 1618
rect 1830 992 1833 1858
rect 1838 1852 1841 1858
rect 1838 1552 1841 1758
rect 1862 1702 1865 2468
rect 1878 2462 1881 2628
rect 1886 2522 1889 3078
rect 1894 2592 1897 3678
rect 1902 3662 1905 3668
rect 1926 3632 1929 3978
rect 1934 3712 1937 3988
rect 1958 3642 1961 4438
rect 1974 4382 1977 4538
rect 1974 4192 1977 4378
rect 1966 4022 1969 4138
rect 1902 3252 1905 3528
rect 1902 2872 1905 3198
rect 1910 3172 1913 3218
rect 1910 3062 1913 3158
rect 1918 3122 1921 3598
rect 1910 2912 1913 2918
rect 1902 2702 1905 2718
rect 1886 2482 1889 2498
rect 1894 2462 1897 2538
rect 1902 2462 1905 2698
rect 1870 2422 1873 2458
rect 1878 2372 1881 2438
rect 1878 2312 1881 2368
rect 1886 2292 1889 2458
rect 1894 2442 1897 2458
rect 1902 2412 1905 2438
rect 1910 2422 1913 2438
rect 1918 2392 1921 2768
rect 1926 2551 1929 3568
rect 1942 3222 1945 3638
rect 1950 3242 1953 3258
rect 1934 2772 1937 3158
rect 1942 3022 1945 3158
rect 1950 3142 1953 3148
rect 1950 3002 1953 3068
rect 1942 2872 1945 2968
rect 1950 2932 1953 2998
rect 1942 2732 1945 2748
rect 1934 2682 1937 2718
rect 1934 2572 1937 2588
rect 1926 2548 1934 2551
rect 1934 2482 1937 2518
rect 1926 2442 1929 2468
rect 1942 2462 1945 2728
rect 1950 2572 1953 2598
rect 1958 2562 1961 3638
rect 1966 3332 1969 4018
rect 1966 3082 1969 3238
rect 1974 3162 1977 4188
rect 1982 4082 1985 4528
rect 2030 4462 2033 4468
rect 1982 3662 1985 3768
rect 1990 3722 1993 4228
rect 1998 4102 2001 4378
rect 1982 3162 1985 3588
rect 1990 3452 1993 3458
rect 1998 3252 2001 3608
rect 2006 3472 2009 3778
rect 1974 3132 1977 3138
rect 1982 3062 1985 3118
rect 1974 3032 1977 3058
rect 1966 2802 1969 2918
rect 1974 2832 1977 3008
rect 1982 3002 1985 3058
rect 1966 2662 1969 2738
rect 1974 2682 1977 2818
rect 1950 2522 1953 2538
rect 1958 2512 1961 2528
rect 1910 2352 1913 2368
rect 1902 2311 1905 2328
rect 1918 2322 1921 2328
rect 1934 2322 1937 2368
rect 1902 2308 1913 2311
rect 1878 2192 1881 2288
rect 1910 2282 1913 2308
rect 1894 2262 1897 2278
rect 1886 2212 1889 2218
rect 1918 2202 1921 2278
rect 1910 2172 1913 2178
rect 1898 2168 1905 2171
rect 1870 1802 1873 2098
rect 1870 1782 1873 1798
rect 1870 1722 1873 1748
rect 1830 962 1833 968
rect 1822 872 1825 888
rect 1838 862 1841 1128
rect 1846 832 1849 1068
rect 1814 622 1817 738
rect 1822 482 1825 828
rect 1854 712 1857 1688
rect 1878 1662 1881 2118
rect 1886 1942 1889 2118
rect 1894 2092 1897 2148
rect 1894 1982 1897 2058
rect 1894 1902 1897 1938
rect 1886 1752 1889 1808
rect 1886 1712 1889 1738
rect 1894 1682 1897 1848
rect 1902 1682 1905 2168
rect 1926 2162 1929 2218
rect 1934 2182 1937 2188
rect 1926 2132 1929 2158
rect 1910 2082 1913 2118
rect 1934 2102 1937 2168
rect 1942 2142 1945 2448
rect 1950 2322 1953 2478
rect 1966 2452 1969 2518
rect 1966 2402 1969 2428
rect 1958 2272 1961 2288
rect 1966 2272 1969 2278
rect 1950 2202 1953 2208
rect 1958 2182 1961 2188
rect 1950 2112 1953 2138
rect 1958 2102 1961 2128
rect 1918 1862 1921 1888
rect 1878 1272 1881 1648
rect 1886 1592 1889 1658
rect 1886 1572 1889 1588
rect 1878 1092 1881 1268
rect 1894 1252 1897 1468
rect 1902 1382 1905 1678
rect 1910 1672 1913 1828
rect 1910 1522 1913 1578
rect 1918 1522 1921 1848
rect 1926 1582 1929 2088
rect 1902 1352 1905 1378
rect 1902 1072 1905 1138
rect 1878 1022 1881 1068
rect 1902 1042 1905 1068
rect 1778 478 1782 481
rect 1718 132 1721 288
rect 1734 262 1737 368
rect 1734 182 1737 258
rect 1742 152 1745 268
rect 1750 152 1753 218
rect 1762 138 1766 141
rect 1774 92 1777 168
rect 1806 132 1809 158
rect 1862 152 1865 658
rect 1910 412 1913 1068
rect 1926 452 1929 1558
rect 1934 1471 1937 1598
rect 1942 1512 1945 2098
rect 1966 2002 1969 2208
rect 1974 2132 1977 2598
rect 1950 1572 1953 1998
rect 1966 1892 1969 1928
rect 1954 1548 1958 1551
rect 1934 1468 1942 1471
rect 1934 782 1937 1468
rect 1958 1372 1961 1528
rect 1942 1292 1945 1298
rect 1942 832 1945 1278
rect 1950 862 1953 1268
rect 1966 1082 1969 1698
rect 1974 1602 1977 2068
rect 1982 1552 1985 2988
rect 1990 2772 1993 3168
rect 1998 2762 2001 3188
rect 2006 3092 2009 3468
rect 2014 3462 2017 3938
rect 2022 3922 2025 4038
rect 2030 3782 2033 4448
rect 2038 4262 2041 4588
rect 2072 4503 2074 4507
rect 2078 4503 2081 4507
rect 2086 4503 2088 4507
rect 2066 4448 2070 4451
rect 2072 4303 2074 4307
rect 2078 4303 2081 4307
rect 2086 4303 2088 4307
rect 2138 4278 2142 4281
rect 2134 4272 2137 4278
rect 2072 4103 2074 4107
rect 2078 4103 2081 4107
rect 2086 4103 2088 4107
rect 2038 3842 2041 3948
rect 2030 3752 2033 3758
rect 2030 3432 2033 3718
rect 2046 3672 2049 4078
rect 2054 3562 2057 4018
rect 2072 3903 2074 3907
rect 2078 3903 2081 3907
rect 2086 3903 2088 3907
rect 2062 3892 2065 3898
rect 2094 3712 2097 3728
rect 2072 3703 2074 3707
rect 2078 3703 2081 3707
rect 2086 3703 2088 3707
rect 2102 3692 2105 4208
rect 2134 4128 2142 4131
rect 2134 4052 2137 4128
rect 2134 4038 2142 4041
rect 2042 3548 2049 3551
rect 2014 2952 2017 3328
rect 2022 3142 2025 3358
rect 2010 2938 2014 2941
rect 2022 2912 2025 3128
rect 1990 2612 1993 2678
rect 1990 2442 1993 2538
rect 1998 2492 2001 2668
rect 2006 2482 2009 2888
rect 2014 2812 2017 2848
rect 2030 2602 2033 3428
rect 2038 3342 2041 3358
rect 2046 3352 2049 3548
rect 2054 3362 2057 3548
rect 2072 3503 2074 3507
rect 2078 3503 2081 3507
rect 2086 3503 2088 3507
rect 2082 3448 2086 3451
rect 2072 3303 2074 3307
rect 2078 3303 2081 3307
rect 2086 3303 2088 3307
rect 2046 3072 2049 3228
rect 2094 3182 2097 3508
rect 2110 3442 2113 3808
rect 2118 3472 2121 3938
rect 2126 3862 2129 3898
rect 2102 3302 2105 3438
rect 2118 3432 2121 3458
rect 2110 3272 2113 3378
rect 2126 3302 2129 3718
rect 2126 3242 2129 3248
rect 2054 3102 2057 3118
rect 2062 3112 2065 3148
rect 2072 3103 2074 3107
rect 2078 3103 2081 3107
rect 2086 3103 2088 3107
rect 2038 2872 2041 2938
rect 2046 2912 2049 2918
rect 2054 2892 2057 3098
rect 2046 2852 2049 2868
rect 2050 2848 2054 2851
rect 2014 2552 2017 2578
rect 2006 2442 2009 2458
rect 1990 2232 1993 2378
rect 2006 2352 2009 2368
rect 1998 2282 2001 2298
rect 1990 2222 1993 2228
rect 1990 2202 1993 2208
rect 1990 2162 1993 2198
rect 1990 1922 1993 1988
rect 1990 1802 1993 1838
rect 1974 1462 1977 1478
rect 1934 552 1937 718
rect 1926 272 1929 448
rect 1934 352 1937 548
rect 1950 302 1953 858
rect 1974 592 1977 1218
rect 1982 782 1985 1268
rect 1990 1172 1993 1798
rect 1998 1732 2001 2238
rect 2006 2072 2009 2318
rect 2014 2032 2017 2518
rect 2014 1982 2017 1988
rect 2006 1892 2009 1978
rect 2022 1952 2025 2578
rect 2030 2182 2033 2508
rect 2030 2032 2033 2108
rect 2038 2092 2041 2728
rect 2046 2672 2049 2798
rect 2054 2692 2057 2698
rect 2062 2622 2065 3088
rect 2072 2903 2074 2907
rect 2078 2903 2081 2907
rect 2086 2903 2088 2907
rect 2086 2762 2089 2788
rect 2094 2732 2097 3128
rect 2102 3112 2105 3178
rect 2134 3102 2137 4038
rect 2142 3322 2145 4018
rect 2150 3782 2153 4268
rect 2158 3972 2161 4728
rect 2214 4541 2217 4788
rect 2230 4662 2233 4738
rect 2214 4538 2225 4541
rect 2174 4342 2177 4348
rect 2166 4002 2169 4148
rect 2166 3932 2169 3958
rect 2102 2832 2105 3098
rect 2102 2802 2105 2828
rect 2118 2802 2121 2828
rect 2072 2703 2074 2707
rect 2078 2703 2081 2707
rect 2086 2703 2088 2707
rect 2082 2658 2086 2661
rect 2046 2592 2049 2618
rect 2046 2522 2049 2558
rect 2046 2432 2049 2498
rect 2054 2421 2057 2608
rect 2046 2418 2057 2421
rect 2062 2422 2065 2548
rect 2070 2542 2073 2628
rect 2086 2552 2089 2568
rect 2072 2503 2074 2507
rect 2078 2503 2081 2507
rect 2086 2503 2088 2507
rect 2046 2372 2049 2418
rect 2046 2202 2049 2358
rect 2054 2312 2057 2388
rect 2062 2262 2065 2418
rect 2086 2372 2089 2378
rect 2072 2303 2074 2307
rect 2078 2303 2081 2307
rect 2086 2303 2088 2307
rect 2062 2248 2070 2251
rect 2046 2082 2049 2168
rect 2054 2012 2057 2218
rect 2062 2212 2065 2248
rect 2094 2242 2097 2728
rect 2102 2712 2105 2748
rect 2102 2332 2105 2668
rect 2110 2542 2113 2778
rect 2102 2252 2105 2288
rect 2070 2192 2073 2218
rect 2078 2192 2081 2228
rect 2062 2162 2065 2188
rect 2102 2142 2105 2168
rect 2072 2103 2074 2107
rect 2078 2103 2081 2107
rect 2086 2103 2088 2107
rect 2078 2052 2081 2078
rect 2022 1842 2025 1908
rect 2038 1742 2041 1828
rect 1990 632 1993 1108
rect 1998 722 2001 1728
rect 2006 1012 2009 1348
rect 2022 1332 2025 1358
rect 2022 1272 2025 1328
rect 2014 1162 2017 1178
rect 2014 1101 2017 1138
rect 2014 1098 2025 1101
rect 2014 1052 2017 1058
rect 2014 1022 2017 1048
rect 2022 852 2025 1098
rect 2010 678 2014 681
rect 1998 652 2001 678
rect 2030 592 2033 1588
rect 2038 1212 2041 1458
rect 2046 1422 2049 1898
rect 2054 1552 2057 2008
rect 2062 1912 2065 1968
rect 2070 1932 2073 1978
rect 2094 1972 2097 2128
rect 2110 2082 2113 2538
rect 2118 2272 2121 2718
rect 2118 2242 2121 2248
rect 2118 2162 2121 2218
rect 2118 2082 2121 2158
rect 2102 2032 2105 2068
rect 2086 1951 2089 1968
rect 2082 1948 2089 1951
rect 2094 1912 2097 1938
rect 2072 1903 2074 1907
rect 2078 1903 2081 1907
rect 2086 1903 2088 1907
rect 2094 1891 2097 1898
rect 2086 1888 2097 1891
rect 2086 1872 2089 1888
rect 2062 1802 2065 1818
rect 2046 1362 2049 1418
rect 2038 672 2041 1208
rect 2046 1162 2049 1358
rect 2054 1142 2057 1408
rect 2062 1352 2065 1798
rect 2070 1752 2073 1828
rect 2078 1782 2081 1798
rect 2086 1752 2089 1838
rect 2072 1703 2074 1707
rect 2078 1703 2081 1707
rect 2086 1703 2088 1707
rect 2086 1682 2089 1688
rect 2094 1672 2097 1878
rect 2102 1692 2105 1718
rect 2098 1558 2102 1561
rect 2094 1512 2097 1528
rect 2072 1503 2074 1507
rect 2078 1503 2081 1507
rect 2086 1503 2088 1507
rect 2086 1422 2089 1468
rect 2086 1402 2089 1408
rect 2094 1342 2097 1438
rect 2072 1303 2074 1307
rect 2078 1303 2081 1307
rect 2086 1303 2088 1307
rect 2074 1268 2078 1271
rect 2086 1262 2089 1268
rect 2046 1132 2049 1138
rect 2062 1122 2065 1138
rect 2030 572 2033 588
rect 1958 312 1961 538
rect 2022 462 2025 558
rect 2046 482 2049 888
rect 2014 352 2017 388
rect 2014 272 2017 348
rect 1882 258 1886 261
rect 1870 82 1873 148
rect 1878 142 1881 188
rect 802 58 806 61
rect 938 58 942 61
rect 1910 52 1913 248
rect 1918 122 1921 188
rect 1930 138 1934 141
rect 1990 92 1993 228
rect 2022 152 2025 458
rect 2054 422 2057 978
rect 2062 942 2065 1118
rect 2072 1103 2074 1107
rect 2078 1103 2081 1107
rect 2086 1103 2088 1107
rect 2094 972 2097 1338
rect 2102 1222 2105 1438
rect 2110 1352 2113 2078
rect 2118 2012 2121 2038
rect 2118 1712 2121 1988
rect 2126 1852 2129 2888
rect 2142 2852 2145 3268
rect 2150 2932 2153 3778
rect 2158 3442 2161 3858
rect 2174 3732 2177 4338
rect 2182 4312 2185 4538
rect 2182 4252 2185 4258
rect 2182 3952 2185 4248
rect 2190 3932 2193 4338
rect 2182 3872 2185 3928
rect 2198 3862 2201 4168
rect 2206 4052 2209 4288
rect 2214 4102 2217 4528
rect 2222 4292 2225 4538
rect 2230 4522 2233 4658
rect 2262 4632 2265 4658
rect 2246 4502 2249 4518
rect 2254 4472 2257 4538
rect 2238 4462 2241 4468
rect 2262 4402 2265 4628
rect 2270 4472 2273 4508
rect 2270 4422 2273 4458
rect 2218 4098 2222 4101
rect 2134 2342 2137 2778
rect 2158 2762 2161 3218
rect 2166 3152 2169 3498
rect 2166 3002 2169 3148
rect 2182 3062 2185 3648
rect 2190 3242 2193 3278
rect 2166 2982 2169 2998
rect 2170 2938 2177 2941
rect 2174 2922 2177 2938
rect 2146 2738 2150 2741
rect 2146 2658 2150 2661
rect 2142 2392 2145 2618
rect 2150 2552 2153 2608
rect 2150 2522 2153 2528
rect 2142 2302 2145 2358
rect 2134 1872 2137 2298
rect 2150 2282 2153 2508
rect 2158 2302 2161 2738
rect 2166 2702 2169 2848
rect 2174 2462 2177 2898
rect 2182 2502 2185 3048
rect 2182 2432 2185 2478
rect 2174 2402 2177 2428
rect 2166 2372 2169 2398
rect 2150 2262 2153 2268
rect 2142 2131 2145 2258
rect 2150 2222 2153 2248
rect 2166 2202 2169 2238
rect 2150 2162 2153 2168
rect 2142 2128 2153 2131
rect 2142 2072 2145 2118
rect 2150 2072 2153 2128
rect 2134 1862 2137 1868
rect 2126 1682 2129 1808
rect 2142 1792 2145 1858
rect 2150 1752 2153 1928
rect 2134 1642 2137 1708
rect 2150 1682 2153 1748
rect 2118 1402 2121 1508
rect 2102 961 2105 1208
rect 2118 1101 2121 1128
rect 2114 1098 2121 1101
rect 2118 992 2121 1028
rect 2094 958 2105 961
rect 2086 952 2089 958
rect 2072 903 2074 907
rect 2078 903 2081 907
rect 2086 903 2088 907
rect 2086 842 2089 888
rect 2062 702 2065 838
rect 2072 703 2074 707
rect 2078 703 2081 707
rect 2086 703 2088 707
rect 2062 562 2065 578
rect 2072 503 2074 507
rect 2078 503 2081 507
rect 2086 503 2088 507
rect 2094 422 2097 958
rect 2106 888 2110 891
rect 2126 802 2129 1498
rect 2134 1402 2137 1428
rect 2142 1312 2145 1638
rect 2150 1502 2153 1648
rect 2158 1622 2161 2178
rect 2150 1392 2153 1498
rect 2158 1492 2161 1618
rect 2166 1602 2169 2198
rect 2174 2152 2177 2378
rect 2182 2162 2185 2388
rect 2182 2092 2185 2098
rect 2158 1471 2161 1488
rect 2158 1468 2166 1471
rect 2158 1332 2161 1428
rect 2166 1422 2169 1458
rect 2162 1258 2166 1261
rect 2134 1032 2137 1108
rect 2142 1032 2145 1248
rect 2150 1072 2153 1168
rect 2150 882 2153 918
rect 2134 862 2137 868
rect 2110 662 2113 698
rect 2106 648 2113 651
rect 2110 402 2113 648
rect 2118 541 2121 748
rect 2142 622 2145 648
rect 2118 538 2126 541
rect 2072 303 2074 307
rect 2078 303 2081 307
rect 2086 303 2088 307
rect 2158 172 2161 1048
rect 2174 692 2177 1848
rect 2182 1762 2185 2088
rect 2190 1742 2193 3238
rect 2198 2902 2201 3758
rect 2206 2822 2209 4008
rect 2214 3222 2217 3908
rect 2198 2752 2201 2768
rect 2206 2712 2209 2818
rect 2198 2502 2201 2598
rect 2214 2521 2217 3198
rect 2222 2992 2225 4058
rect 2230 3692 2233 3758
rect 2238 3652 2241 3808
rect 2230 3172 2233 3588
rect 2238 3422 2241 3448
rect 2222 2952 2225 2988
rect 2230 2952 2233 3038
rect 2222 2862 2225 2868
rect 2210 2518 2217 2521
rect 2198 2352 2201 2458
rect 2198 2162 2201 2298
rect 2206 2292 2209 2298
rect 2206 2212 2209 2228
rect 2206 2022 2209 2198
rect 2198 1932 2201 1948
rect 2198 1752 2201 1848
rect 2190 1722 2193 1728
rect 2182 1681 2185 1718
rect 2190 1692 2193 1698
rect 2182 1678 2190 1681
rect 2182 1432 2185 1478
rect 2190 1472 2193 1558
rect 2198 1552 2201 1748
rect 2206 1582 2209 1858
rect 2206 1552 2209 1558
rect 2198 1482 2201 1488
rect 2190 1451 2193 1458
rect 2190 1448 2198 1451
rect 2190 1132 2193 1438
rect 2202 1288 2206 1291
rect 2182 352 2185 1098
rect 2198 942 2201 1138
rect 2206 1062 2209 1248
rect 2214 1232 2217 2498
rect 2222 1742 2225 2728
rect 2230 2522 2233 2588
rect 2238 2542 2241 3418
rect 2246 3272 2249 4398
rect 2262 4362 2265 4398
rect 2286 4362 2289 4568
rect 2262 4102 2265 4358
rect 2262 3962 2265 4098
rect 2262 3692 2265 3878
rect 2278 3792 2281 4358
rect 2286 4152 2289 4258
rect 2294 4242 2297 4448
rect 2302 4392 2305 4468
rect 2310 4252 2313 4478
rect 2294 3912 2297 4238
rect 2302 4102 2305 4248
rect 2310 4102 2313 4248
rect 2318 4172 2321 4558
rect 2326 4172 2329 4178
rect 2254 3272 2257 3688
rect 2270 3222 2273 3748
rect 2278 3671 2281 3688
rect 2278 3668 2286 3671
rect 2294 3612 2297 3908
rect 2318 3842 2321 4148
rect 2334 4142 2337 4738
rect 2350 4692 2353 4868
rect 2370 4858 2374 4861
rect 2438 4822 2441 4868
rect 3190 4858 3198 4861
rect 2342 4322 2345 4328
rect 2350 4272 2353 4688
rect 2366 4432 2369 4458
rect 2378 4448 2382 4451
rect 2342 4062 2345 4258
rect 2366 4202 2369 4368
rect 2374 4262 2377 4288
rect 2350 4082 2353 4178
rect 2358 4062 2361 4068
rect 2330 3918 2334 3921
rect 2282 3348 2286 3351
rect 2286 3292 2289 3298
rect 2262 2992 2265 3088
rect 2270 3032 2273 3108
rect 2278 3032 2281 3288
rect 2294 3092 2297 3588
rect 2290 3048 2294 3051
rect 2246 2712 2249 2748
rect 2246 2682 2249 2708
rect 2262 2702 2265 2988
rect 2270 2732 2273 3028
rect 2246 2552 2249 2578
rect 2238 2442 2241 2468
rect 2230 2252 2233 2378
rect 2246 2372 2249 2468
rect 2238 2312 2241 2328
rect 2230 1892 2233 2178
rect 2238 1952 2241 2278
rect 2246 2062 2249 2358
rect 2254 2272 2257 2648
rect 2262 2402 2265 2578
rect 2270 2462 2273 2668
rect 2278 2632 2281 2658
rect 2254 2082 2257 2108
rect 2246 1982 2249 2058
rect 2246 1772 2249 1838
rect 2238 1752 2241 1768
rect 2254 1672 2257 2068
rect 2262 1992 2265 2348
rect 2270 2282 2273 2288
rect 2270 2272 2273 2278
rect 2270 2192 2273 2218
rect 2270 2112 2273 2148
rect 2278 2102 2281 2538
rect 2286 2402 2289 2938
rect 2294 2632 2297 2648
rect 2294 2452 2297 2578
rect 2302 2352 2305 3828
rect 2314 3808 2318 3811
rect 2326 3802 2329 3878
rect 2342 3872 2345 4058
rect 2350 3972 2353 4058
rect 2366 3992 2369 4158
rect 2326 3622 2329 3798
rect 2334 3611 2337 3818
rect 2326 3608 2337 3611
rect 2310 3252 2313 3518
rect 2310 2942 2313 3248
rect 2318 3172 2321 3268
rect 2318 3072 2321 3168
rect 2326 2942 2329 3608
rect 2334 3342 2337 3438
rect 2334 3072 2337 3208
rect 2342 3022 2345 3728
rect 2350 3612 2353 3968
rect 2358 3672 2361 3678
rect 2354 3538 2358 3541
rect 2318 2938 2326 2941
rect 2318 2902 2321 2938
rect 2310 2342 2313 2848
rect 2334 2662 2337 2858
rect 2350 2732 2353 3268
rect 2358 2992 2361 3138
rect 2358 2742 2361 2748
rect 2334 2592 2337 2608
rect 2318 2558 2326 2561
rect 2318 2552 2321 2558
rect 2350 2552 2353 2698
rect 2334 2491 2337 2548
rect 2342 2512 2345 2518
rect 2326 2488 2337 2491
rect 2318 2452 2321 2468
rect 2310 2332 2313 2338
rect 2286 2172 2289 2288
rect 2294 2172 2297 2328
rect 2318 2192 2321 2348
rect 2214 1222 2217 1228
rect 2222 1042 2225 1528
rect 2230 1082 2233 1578
rect 2238 1552 2241 1578
rect 2238 1072 2241 1538
rect 2262 1512 2265 1588
rect 2246 1448 2254 1451
rect 2246 1432 2249 1448
rect 2246 1412 2249 1428
rect 2270 1421 2273 2048
rect 2278 1982 2281 2008
rect 2286 1892 2289 1908
rect 2278 1572 2281 1738
rect 2286 1552 2289 1618
rect 2282 1528 2286 1531
rect 2270 1418 2281 1421
rect 2246 1152 2249 1398
rect 2270 1292 2273 1328
rect 2222 952 2225 1018
rect 2206 682 2209 908
rect 2214 852 2217 938
rect 2246 742 2249 1098
rect 2254 892 2257 1148
rect 2262 1061 2265 1208
rect 2262 1058 2270 1061
rect 2270 822 2273 848
rect 2246 542 2249 548
rect 2262 372 2265 648
rect 2270 492 2273 728
rect 2278 462 2281 1418
rect 2286 782 2289 1478
rect 2294 1272 2297 1648
rect 2302 1582 2305 2158
rect 2310 2102 2313 2108
rect 2310 2071 2313 2078
rect 2310 2068 2318 2071
rect 2310 1962 2313 1998
rect 2310 1582 2313 1948
rect 2326 1942 2329 2488
rect 2334 2392 2337 2458
rect 2334 2312 2337 2318
rect 2350 2252 2353 2528
rect 2334 2012 2337 2228
rect 2358 2222 2361 2658
rect 2306 1548 2310 1551
rect 2302 1392 2305 1418
rect 2310 1352 2313 1358
rect 2294 751 2297 1168
rect 2294 748 2302 751
rect 2302 562 2305 708
rect 2302 541 2305 558
rect 2298 538 2305 541
rect 2310 522 2313 898
rect 2318 702 2321 1898
rect 2330 1858 2334 1861
rect 2326 1482 2329 1628
rect 2326 1282 2329 1358
rect 2334 852 2337 1848
rect 2342 1602 2345 2168
rect 2350 2082 2353 2178
rect 2350 1862 2353 1888
rect 2358 1852 2361 2018
rect 2358 1822 2361 1848
rect 2366 1672 2369 3938
rect 2374 3842 2377 4188
rect 2374 3822 2377 3838
rect 2374 3632 2377 3808
rect 2382 3742 2385 4248
rect 2390 4192 2393 4358
rect 2390 4062 2393 4118
rect 2398 3962 2401 4498
rect 2422 4472 2425 4478
rect 2406 4352 2409 4458
rect 2430 4282 2433 4768
rect 2438 4272 2441 4818
rect 2584 4803 2586 4807
rect 2590 4803 2593 4807
rect 2598 4803 2600 4807
rect 2502 4532 2505 4538
rect 2478 4362 2481 4488
rect 2494 4432 2497 4528
rect 2422 4142 2425 4148
rect 2422 4072 2425 4078
rect 2422 3872 2425 3878
rect 2430 3862 2433 4158
rect 2446 4142 2449 4328
rect 2438 4062 2441 4068
rect 2422 3852 2425 3858
rect 2402 3848 2409 3851
rect 2406 3812 2409 3848
rect 2390 3772 2393 3788
rect 2374 3452 2377 3628
rect 2390 3502 2393 3668
rect 2414 3651 2417 3808
rect 2422 3662 2425 3848
rect 2430 3742 2433 3768
rect 2414 3648 2425 3651
rect 2390 3482 2393 3498
rect 2374 2702 2377 3448
rect 2382 3262 2385 3368
rect 2382 3192 2385 3258
rect 2374 2682 2377 2698
rect 2374 2412 2377 2668
rect 2382 2662 2385 2838
rect 2390 2632 2393 3458
rect 2398 3012 2401 3528
rect 2398 2892 2401 2928
rect 2406 2792 2409 3648
rect 2414 3122 2417 3548
rect 2422 3522 2425 3648
rect 2422 3172 2425 3518
rect 2430 3142 2433 3738
rect 2438 3552 2441 3738
rect 2438 3542 2441 3548
rect 2446 3192 2449 4138
rect 2454 4052 2457 4218
rect 2470 4062 2473 4148
rect 2462 3682 2465 3718
rect 2470 3422 2473 4058
rect 2494 3692 2497 3748
rect 2478 3672 2481 3678
rect 2478 3542 2481 3618
rect 2502 3572 2505 4318
rect 2478 3492 2481 3538
rect 2458 3358 2465 3361
rect 2462 3342 2465 3358
rect 2442 3168 2449 3171
rect 2398 2552 2401 2568
rect 2382 2412 2385 2508
rect 2406 2471 2409 2488
rect 2402 2468 2409 2471
rect 2374 2342 2377 2388
rect 2390 2362 2393 2458
rect 2398 2442 2401 2458
rect 2406 2402 2409 2438
rect 2414 2362 2417 2808
rect 2422 2522 2425 3058
rect 2438 3042 2441 3048
rect 2438 2972 2441 3028
rect 2422 2472 2425 2478
rect 2414 2262 2417 2358
rect 2414 2152 2417 2168
rect 2394 2088 2398 2091
rect 2374 1862 2377 1888
rect 2374 1652 2377 1718
rect 2390 1682 2393 1878
rect 2334 412 2337 778
rect 2342 522 2345 1498
rect 2350 812 2353 928
rect 2366 882 2369 1588
rect 2390 1542 2393 1628
rect 2398 1402 2401 1668
rect 2406 1422 2409 1988
rect 2414 1921 2417 1978
rect 2422 1932 2425 2268
rect 2430 1992 2433 2798
rect 2414 1918 2422 1921
rect 2430 1892 2433 1898
rect 2414 1722 2417 1748
rect 2422 1722 2425 1838
rect 2430 1782 2433 1848
rect 2430 1732 2433 1748
rect 2414 1632 2417 1718
rect 2438 1682 2441 2968
rect 2446 2302 2449 3168
rect 2454 2822 2457 3338
rect 2462 3262 2465 3298
rect 2454 2672 2457 2768
rect 2454 2352 2457 2618
rect 2462 2512 2465 2898
rect 2470 2872 2473 3118
rect 2486 3072 2489 3338
rect 2486 3062 2489 3068
rect 2486 2932 2489 2958
rect 2494 2952 2497 3398
rect 2502 3352 2505 3448
rect 2510 3262 2513 4208
rect 2518 4091 2521 4758
rect 2658 4738 2662 4741
rect 2526 4582 2529 4728
rect 2526 4532 2529 4548
rect 2534 4542 2537 4628
rect 2550 4622 2553 4688
rect 2526 4422 2529 4528
rect 2534 4382 2537 4538
rect 2534 4352 2537 4358
rect 2518 4088 2526 4091
rect 2518 3492 2521 4068
rect 2526 3672 2529 3908
rect 2542 3832 2545 4618
rect 2566 4542 2569 4638
rect 2584 4603 2586 4607
rect 2590 4603 2593 4607
rect 2598 4603 2600 4607
rect 2566 4512 2569 4538
rect 2678 4482 2681 4538
rect 2584 4403 2586 4407
rect 2590 4403 2593 4407
rect 2598 4403 2600 4407
rect 2550 4342 2553 4348
rect 2584 4203 2586 4207
rect 2590 4203 2593 4207
rect 2598 4203 2600 4207
rect 2606 4202 2609 4298
rect 2550 4012 2553 4058
rect 2534 3462 2537 3758
rect 2502 3082 2505 3138
rect 2510 3132 2513 3218
rect 2542 3122 2545 3808
rect 2550 3512 2553 4008
rect 2558 3502 2561 3858
rect 2566 3672 2569 3738
rect 2550 3332 2553 3348
rect 2558 3322 2561 3328
rect 2522 3108 2526 3111
rect 2518 3072 2521 3078
rect 2526 3072 2529 3078
rect 2502 3052 2505 3058
rect 2510 2902 2513 3048
rect 2470 2772 2473 2848
rect 2478 2812 2481 2848
rect 2510 2812 2513 2818
rect 2462 2452 2465 2458
rect 2446 2202 2449 2298
rect 2446 2142 2449 2158
rect 2446 1692 2449 1888
rect 2422 1442 2425 1648
rect 2446 1642 2449 1668
rect 2374 932 2377 998
rect 2382 932 2385 1348
rect 2390 1342 2393 1348
rect 2398 1312 2401 1398
rect 2422 1302 2425 1418
rect 2426 1258 2433 1261
rect 2362 738 2369 741
rect 2366 662 2369 738
rect 2374 672 2377 928
rect 2414 722 2417 1248
rect 2430 1032 2433 1258
rect 2438 762 2441 1488
rect 2418 718 2422 721
rect 2422 642 2425 648
rect 2398 522 2401 588
rect 2342 482 2345 518
rect 2350 392 2353 488
rect 2398 472 2401 518
rect 2422 472 2425 638
rect 2182 292 2185 348
rect 2166 262 2169 268
rect 2238 262 2241 268
rect 2210 258 2214 261
rect 2182 142 2185 208
rect 2286 142 2289 338
rect 2382 232 2385 448
rect 2438 302 2441 758
rect 2454 742 2457 2258
rect 2462 2172 2465 2238
rect 2462 1651 2465 2168
rect 2470 2162 2473 2768
rect 2490 2678 2494 2681
rect 2478 2442 2481 2458
rect 2494 2232 2497 2508
rect 2502 2372 2505 2698
rect 2510 2592 2513 2678
rect 2518 2602 2521 2778
rect 2510 2362 2513 2478
rect 2486 2212 2489 2218
rect 2486 1972 2489 2198
rect 2494 2012 2497 2058
rect 2502 1962 2505 2358
rect 2470 1942 2473 1948
rect 2494 1761 2497 1948
rect 2486 1758 2497 1761
rect 2486 1732 2489 1758
rect 2494 1742 2497 1748
rect 2462 1648 2470 1651
rect 2462 1502 2465 1548
rect 2462 892 2465 1458
rect 2470 892 2473 1648
rect 2486 1582 2489 1728
rect 2478 1232 2481 1378
rect 2478 912 2481 1008
rect 2486 952 2489 1348
rect 2502 822 2505 1808
rect 2510 1242 2513 2148
rect 2518 2032 2521 2498
rect 2526 2362 2529 3068
rect 2534 3042 2537 3088
rect 2550 3072 2553 3178
rect 2534 3012 2537 3038
rect 2534 2972 2537 3008
rect 2534 2942 2537 2948
rect 2534 2592 2537 2878
rect 2554 2868 2558 2871
rect 2542 2732 2545 2868
rect 2554 2748 2561 2751
rect 2558 2742 2561 2748
rect 2542 2642 2545 2648
rect 2558 2622 2561 2738
rect 2526 1802 2529 2168
rect 2534 2152 2537 2588
rect 2566 2572 2569 3668
rect 2574 3532 2577 4048
rect 2606 4022 2609 4068
rect 2584 4003 2586 4007
rect 2590 4003 2593 4007
rect 2598 4003 2600 4007
rect 2606 3972 2609 3998
rect 2598 3862 2601 3918
rect 2584 3803 2586 3807
rect 2590 3803 2593 3807
rect 2598 3803 2600 3807
rect 2614 3741 2617 4408
rect 2630 4262 2633 4298
rect 2622 3862 2625 3868
rect 2630 3782 2633 3938
rect 2614 3738 2622 3741
rect 2584 3603 2586 3607
rect 2590 3603 2593 3607
rect 2598 3603 2600 3607
rect 2606 3582 2609 3708
rect 2614 3592 2617 3648
rect 2614 3522 2617 3588
rect 2622 3491 2625 3698
rect 2618 3488 2625 3491
rect 2584 3403 2586 3407
rect 2590 3403 2593 3407
rect 2598 3403 2600 3407
rect 2574 3092 2577 3398
rect 2614 3262 2617 3468
rect 2584 3203 2586 3207
rect 2590 3203 2593 3207
rect 2598 3203 2600 3207
rect 2606 3172 2609 3198
rect 2542 2332 2545 2528
rect 2550 2412 2553 2458
rect 2534 1972 2537 2128
rect 2542 2022 2545 2278
rect 2542 2008 2550 2011
rect 2534 1912 2537 1918
rect 2542 1912 2545 2008
rect 2518 1302 2521 1558
rect 2526 1152 2529 1658
rect 2558 1392 2561 2228
rect 2566 1952 2569 2368
rect 2574 2242 2577 3068
rect 2614 3032 2617 3168
rect 2622 3122 2625 3438
rect 2630 3342 2633 3778
rect 2638 3752 2641 4088
rect 2646 3802 2649 4328
rect 2662 4258 2670 4261
rect 2662 4222 2665 4258
rect 2654 4012 2657 4048
rect 2662 4032 2665 4218
rect 2646 3742 2649 3758
rect 2646 3612 2649 3738
rect 2654 3482 2657 3998
rect 2662 3742 2665 3778
rect 2666 3648 2670 3651
rect 2584 3003 2586 3007
rect 2590 3003 2593 3007
rect 2598 3003 2600 3007
rect 2606 2952 2609 3008
rect 2606 2932 2609 2948
rect 2584 2803 2586 2807
rect 2590 2803 2593 2807
rect 2598 2803 2600 2807
rect 2606 2622 2609 2918
rect 2614 2702 2617 3028
rect 2630 2952 2633 3298
rect 2654 3282 2657 3428
rect 2670 3352 2673 3508
rect 2678 3482 2681 3918
rect 2686 3822 2689 4858
rect 3010 4738 3014 4741
rect 3096 4703 3098 4707
rect 3102 4703 3105 4707
rect 3110 4703 3112 4707
rect 2694 4512 2697 4658
rect 2718 4652 2721 4658
rect 2702 4472 2705 4578
rect 2714 4468 2718 4471
rect 2726 4372 2729 4488
rect 2734 4452 2737 4458
rect 2686 3642 2689 3758
rect 2678 3472 2681 3478
rect 2682 3348 2686 3351
rect 2638 3232 2641 3268
rect 2630 2942 2633 2948
rect 2622 2922 2625 2938
rect 2622 2802 2625 2908
rect 2630 2852 2633 2908
rect 2584 2603 2586 2607
rect 2590 2603 2593 2607
rect 2598 2603 2600 2607
rect 2606 2492 2609 2618
rect 2614 2462 2617 2608
rect 2584 2403 2586 2407
rect 2590 2403 2593 2407
rect 2598 2403 2600 2407
rect 2582 2342 2585 2368
rect 2584 2203 2586 2207
rect 2590 2203 2593 2207
rect 2598 2203 2600 2207
rect 2582 2092 2585 2188
rect 2584 2003 2586 2007
rect 2590 2003 2593 2007
rect 2598 2003 2600 2007
rect 2558 1371 2561 1378
rect 2554 1368 2561 1371
rect 2510 1032 2513 1058
rect 2518 852 2521 1088
rect 2526 942 2529 1138
rect 2534 862 2537 1338
rect 2546 1328 2550 1331
rect 2542 972 2545 1208
rect 2566 972 2569 1868
rect 2574 1672 2577 1998
rect 2584 1803 2586 1807
rect 2590 1803 2593 1807
rect 2598 1803 2600 1807
rect 2574 1402 2577 1658
rect 2584 1603 2586 1607
rect 2590 1603 2593 1607
rect 2598 1603 2600 1607
rect 2584 1403 2586 1407
rect 2590 1403 2593 1407
rect 2598 1403 2600 1407
rect 2574 1382 2577 1388
rect 2574 1272 2577 1338
rect 2582 1252 2585 1278
rect 2584 1203 2586 1207
rect 2590 1203 2593 1207
rect 2598 1203 2600 1207
rect 2606 1132 2609 2448
rect 2614 2432 2617 2448
rect 2622 2342 2625 2638
rect 2638 2542 2641 3208
rect 2646 2952 2649 2958
rect 2646 2892 2649 2928
rect 2654 2871 2657 3208
rect 2662 3142 2665 3268
rect 2694 3252 2697 4198
rect 2702 4102 2705 4368
rect 2710 4052 2713 4288
rect 2742 4272 2745 4688
rect 2750 4352 2753 4488
rect 2742 4258 2750 4261
rect 2726 3902 2729 4148
rect 2702 3762 2705 3848
rect 2662 2982 2665 2998
rect 2686 2971 2689 3048
rect 2682 2968 2689 2971
rect 2702 2972 2705 3758
rect 2662 2902 2665 2938
rect 2650 2868 2657 2871
rect 2666 2868 2670 2871
rect 2654 2722 2657 2868
rect 2678 2542 2681 2828
rect 2702 2712 2705 2728
rect 2702 2662 2705 2688
rect 2638 2502 2641 2528
rect 2630 2372 2633 2488
rect 2638 2471 2641 2498
rect 2646 2482 2649 2518
rect 2638 2468 2646 2471
rect 2654 2412 2657 2468
rect 2630 2232 2633 2348
rect 2670 2342 2673 2348
rect 2678 2332 2681 2538
rect 2614 1942 2617 2008
rect 2614 1472 2617 1888
rect 2622 1872 2625 2068
rect 2630 1932 2633 1968
rect 2622 1212 2625 1778
rect 2638 1361 2641 1778
rect 2646 1742 2649 1878
rect 2654 1792 2657 2218
rect 2670 2082 2673 2118
rect 2654 1752 2657 1788
rect 2638 1358 2646 1361
rect 2574 1002 2577 1098
rect 2590 1082 2593 1118
rect 2590 1062 2593 1078
rect 2584 1003 2586 1007
rect 2590 1003 2593 1007
rect 2598 1003 2600 1007
rect 2606 982 2609 1078
rect 2614 1012 2617 1188
rect 2622 1182 2625 1188
rect 2630 1172 2633 1358
rect 2642 1258 2646 1261
rect 2654 1172 2657 1358
rect 2654 1062 2657 1108
rect 2626 1058 2630 1061
rect 2662 982 2665 2048
rect 2558 962 2561 968
rect 2658 948 2662 951
rect 2630 862 2633 898
rect 2638 892 2641 918
rect 2646 852 2649 948
rect 2502 802 2505 818
rect 2606 812 2609 848
rect 2584 803 2586 807
rect 2590 803 2593 807
rect 2598 803 2600 807
rect 2614 752 2617 778
rect 2522 748 2526 751
rect 2622 632 2625 738
rect 2630 662 2633 678
rect 2654 672 2657 928
rect 2654 662 2657 668
rect 2584 603 2586 607
rect 2590 603 2593 607
rect 2598 603 2600 607
rect 2646 472 2649 478
rect 2654 472 2657 658
rect 2670 482 2673 1668
rect 2678 1372 2681 2078
rect 2686 1472 2689 2568
rect 2694 2532 2697 2648
rect 2702 2642 2705 2648
rect 2710 2612 2713 3598
rect 2718 3272 2721 3828
rect 2726 3642 2729 3858
rect 2734 3352 2737 3688
rect 2742 3292 2745 4258
rect 2750 3692 2753 4128
rect 2758 4072 2761 4628
rect 2798 4352 2801 4588
rect 2758 3922 2761 3968
rect 2766 3952 2769 4228
rect 2774 4082 2777 4348
rect 2798 4342 2801 4348
rect 2878 4342 2881 4428
rect 2886 4342 2889 4448
rect 2782 4102 2785 4328
rect 2830 4302 2833 4338
rect 2782 4001 2785 4098
rect 2774 3998 2785 4001
rect 2774 3871 2777 3998
rect 2774 3868 2782 3871
rect 2750 3472 2753 3668
rect 2758 3382 2761 3768
rect 2774 3392 2777 3858
rect 2782 3442 2785 3868
rect 2738 3248 2745 3251
rect 2718 3042 2721 3188
rect 2742 3102 2745 3248
rect 2718 2732 2721 3038
rect 2726 3022 2729 3048
rect 2734 2962 2737 3018
rect 2710 2552 2713 2598
rect 2702 2542 2705 2548
rect 2706 2468 2710 2471
rect 2694 2362 2697 2458
rect 2706 2368 2710 2371
rect 2694 2212 2697 2258
rect 2710 2062 2713 2128
rect 2694 1522 2697 1988
rect 2702 1862 2705 1948
rect 2702 1752 2705 1828
rect 2702 1742 2705 1748
rect 2678 1142 2681 1158
rect 2678 1072 2681 1138
rect 2678 952 2681 988
rect 2686 722 2689 1448
rect 2694 1062 2697 1488
rect 2702 1172 2705 1468
rect 2710 1222 2713 1928
rect 2702 1151 2705 1168
rect 2702 1148 2710 1151
rect 2694 732 2697 1058
rect 2702 832 2705 1138
rect 2718 1071 2721 2718
rect 2726 2012 2729 2578
rect 2734 2381 2737 2958
rect 2750 2832 2753 3198
rect 2758 2962 2761 3038
rect 2742 2552 2745 2808
rect 2758 2582 2761 2918
rect 2766 2682 2769 3378
rect 2774 3092 2777 3248
rect 2774 2902 2777 2968
rect 2782 2912 2785 3368
rect 2790 3302 2793 4098
rect 2798 3802 2801 4148
rect 2806 4112 2809 4188
rect 2822 4142 2825 4148
rect 2806 3912 2809 3988
rect 2790 3132 2793 3288
rect 2798 2862 2801 3248
rect 2806 2892 2809 3788
rect 2814 3472 2817 4138
rect 2830 4072 2833 4098
rect 2826 4058 2830 4061
rect 2838 4022 2841 4298
rect 2846 4292 2849 4318
rect 2846 4132 2849 4138
rect 2846 4002 2849 4018
rect 2842 3958 2846 3961
rect 2822 3922 2825 3928
rect 2858 3918 2862 3921
rect 2870 3842 2873 4188
rect 2910 4172 2913 4548
rect 2966 4332 2969 4538
rect 2974 4472 2977 4558
rect 2990 4552 2993 4658
rect 3022 4561 3025 4688
rect 3030 4652 3033 4658
rect 3018 4558 3025 4561
rect 2998 4542 3001 4548
rect 2990 4532 2993 4538
rect 2982 4451 2985 4528
rect 2978 4448 2985 4451
rect 2894 4062 2897 4118
rect 2882 3958 2886 3961
rect 2882 3928 2886 3931
rect 2902 3832 2905 3928
rect 2918 3832 2921 4258
rect 2926 4222 2929 4238
rect 2822 3342 2825 3388
rect 2818 3338 2822 3341
rect 2814 3222 2817 3258
rect 2814 3212 2817 3218
rect 2814 2922 2817 3208
rect 2822 2832 2825 3078
rect 2830 2842 2833 3098
rect 2838 3032 2841 3748
rect 2902 3742 2905 3758
rect 2850 3738 2857 3741
rect 2854 3552 2857 3738
rect 2838 2872 2841 2988
rect 2742 2502 2745 2508
rect 2742 2472 2745 2488
rect 2766 2462 2769 2678
rect 2734 2378 2745 2381
rect 2734 2042 2737 2368
rect 2742 2282 2745 2378
rect 2726 1551 2729 1838
rect 2734 1572 2737 1748
rect 2742 1622 2745 2218
rect 2750 1611 2753 2408
rect 2782 2312 2785 2648
rect 2790 2222 2793 2808
rect 2822 2791 2825 2828
rect 2818 2788 2825 2791
rect 2834 2788 2838 2791
rect 2814 2572 2817 2628
rect 2822 2522 2825 2578
rect 2798 2432 2801 2458
rect 2806 2172 2809 2508
rect 2814 2322 2817 2478
rect 2822 2462 2825 2478
rect 2822 2352 2825 2358
rect 2822 2332 2825 2348
rect 2814 2202 2817 2298
rect 2830 2141 2833 2788
rect 2854 2782 2857 3238
rect 2862 3162 2865 3528
rect 2882 3458 2886 3461
rect 2902 3342 2905 3348
rect 2890 3318 2894 3321
rect 2926 3302 2929 4168
rect 2950 4152 2953 4158
rect 2934 3772 2937 4068
rect 2958 4012 2961 4258
rect 2966 4212 2969 4278
rect 2942 3832 2945 3858
rect 2942 3672 2945 3828
rect 2950 3812 2953 3958
rect 2942 3482 2945 3668
rect 2862 3072 2865 3158
rect 2870 3122 2873 3248
rect 2838 2722 2841 2758
rect 2850 2718 2854 2721
rect 2842 2708 2846 2711
rect 2850 2668 2854 2671
rect 2862 2622 2865 3048
rect 2878 2912 2881 3128
rect 2886 2902 2889 2948
rect 2878 2741 2881 2828
rect 2874 2738 2881 2741
rect 2846 2552 2849 2568
rect 2846 2472 2849 2538
rect 2838 2432 2841 2448
rect 2822 2138 2833 2141
rect 2790 2062 2793 2068
rect 2822 2022 2825 2138
rect 2782 2008 2790 2011
rect 2782 1922 2785 2008
rect 2762 1678 2766 1681
rect 2742 1608 2753 1611
rect 2726 1548 2734 1551
rect 2742 1412 2745 1608
rect 2774 1602 2777 1708
rect 2782 1682 2785 1768
rect 2782 1672 2785 1678
rect 2754 1528 2758 1531
rect 2790 1502 2793 1918
rect 2734 1338 2742 1341
rect 2734 1102 2737 1338
rect 2718 1068 2726 1071
rect 2722 1058 2726 1061
rect 2734 1022 2737 1088
rect 2742 992 2745 1278
rect 2438 282 2441 298
rect 2494 172 2497 448
rect 2654 412 2657 468
rect 2584 403 2586 407
rect 2590 403 2593 407
rect 2598 403 2600 407
rect 2670 372 2673 478
rect 2682 348 2686 351
rect 2514 148 2518 151
rect 2370 118 2374 121
rect 2072 103 2074 107
rect 2078 103 2081 107
rect 2086 103 2088 107
rect 2566 82 2569 258
rect 2694 212 2697 728
rect 2750 632 2753 1488
rect 2758 1072 2761 1348
rect 2766 1162 2769 1198
rect 2758 682 2761 958
rect 2766 792 2769 838
rect 2702 272 2705 408
rect 2718 392 2721 478
rect 2718 362 2721 388
rect 2726 272 2729 578
rect 2774 402 2777 1498
rect 2798 1492 2801 1988
rect 2806 1892 2809 1908
rect 2806 1872 2809 1888
rect 2830 1652 2833 2048
rect 2838 1742 2841 2158
rect 2846 1702 2849 2228
rect 2854 2042 2857 2568
rect 2862 2022 2865 2528
rect 2870 1982 2873 2658
rect 2878 2622 2881 2668
rect 2878 2342 2881 2618
rect 2886 2482 2889 2558
rect 2894 2442 2897 3258
rect 2902 3082 2905 3228
rect 2918 3112 2921 3178
rect 2942 3152 2945 3358
rect 2934 3142 2937 3148
rect 2902 2782 2905 3068
rect 2902 2662 2905 2668
rect 2902 2281 2905 2518
rect 2910 2312 2913 3018
rect 2918 2572 2921 2888
rect 2942 2742 2945 3148
rect 2950 2992 2953 3808
rect 2958 3562 2961 3858
rect 2966 3792 2969 4148
rect 2982 3952 2985 4448
rect 2990 3972 2993 4528
rect 3002 4018 3006 4021
rect 3014 3942 3017 4508
rect 3030 4282 3033 4458
rect 3014 3908 3022 3911
rect 2998 3782 3001 3858
rect 2902 2278 2910 2281
rect 2858 1848 2862 1851
rect 2854 1762 2857 1798
rect 2870 1712 2873 1788
rect 2782 1042 2785 1488
rect 2782 952 2785 1038
rect 2798 802 2801 1438
rect 2806 1262 2809 1468
rect 2814 982 2817 1518
rect 2798 761 2801 768
rect 2798 758 2806 761
rect 2790 442 2793 748
rect 2802 548 2806 551
rect 2814 522 2817 878
rect 2822 832 2825 1348
rect 2830 1221 2833 1648
rect 2846 1552 2849 1578
rect 2862 1552 2865 1648
rect 2870 1622 2873 1708
rect 2854 1532 2857 1538
rect 2838 1382 2841 1388
rect 2830 1218 2841 1221
rect 2830 1022 2833 1208
rect 2838 962 2841 1218
rect 2584 203 2586 207
rect 2590 203 2593 207
rect 2598 203 2600 207
rect 2702 152 2705 268
rect 2726 132 2729 198
rect 2734 171 2737 328
rect 2778 268 2782 271
rect 2814 242 2817 518
rect 2830 452 2833 468
rect 2734 168 2742 171
rect 2586 128 2590 131
rect 2742 92 2745 128
rect 2750 122 2753 168
rect 2814 112 2817 238
rect 2838 142 2841 918
rect 2846 862 2849 1518
rect 2862 1512 2865 1548
rect 2870 1332 2873 1618
rect 2878 1552 2881 2268
rect 2894 1622 2897 2068
rect 2886 1372 2889 1558
rect 2894 1522 2897 1528
rect 2902 1522 2905 1918
rect 2910 1582 2913 2278
rect 2918 1882 2921 2328
rect 2926 2152 2929 2558
rect 2934 2502 2937 2508
rect 2934 2292 2937 2358
rect 2942 2312 2945 2738
rect 2950 2532 2953 2948
rect 2958 2612 2961 3528
rect 2966 3482 2969 3668
rect 2998 3662 3001 3778
rect 2974 3512 2977 3598
rect 3014 3542 3017 3908
rect 3030 3762 3033 4088
rect 3038 3952 3041 4658
rect 3190 4652 3193 4858
rect 3222 4632 3225 4858
rect 3608 4803 3610 4807
rect 3614 4803 3617 4807
rect 3622 4803 3624 4807
rect 3246 4682 3249 4798
rect 3382 4698 3390 4701
rect 3298 4638 3302 4641
rect 3038 3812 3041 3948
rect 3046 3872 3049 3948
rect 3034 3758 3041 3761
rect 3030 3612 3033 3708
rect 2966 3382 2969 3388
rect 2966 3182 2969 3258
rect 2974 3182 2977 3348
rect 2966 3142 2969 3148
rect 2974 3132 2977 3138
rect 2974 2941 2977 2948
rect 2982 2942 2985 3508
rect 2990 3102 2993 3248
rect 2998 3152 3001 3448
rect 2974 2938 2982 2941
rect 2978 2858 2985 2861
rect 2982 2842 2985 2858
rect 2958 2382 2961 2608
rect 2966 2302 2969 2348
rect 2950 2262 2953 2268
rect 2958 2212 2961 2288
rect 2966 2272 2969 2298
rect 2966 2212 2969 2228
rect 2862 1322 2865 1328
rect 2846 412 2849 618
rect 2854 552 2857 1298
rect 2870 902 2873 1318
rect 2850 408 2857 411
rect 2846 172 2849 398
rect 2854 162 2857 408
rect 2862 222 2865 368
rect 2870 312 2873 718
rect 2878 472 2881 1258
rect 2894 862 2897 868
rect 2894 332 2897 858
rect 2902 712 2905 998
rect 2910 762 2913 1548
rect 2918 1432 2921 1878
rect 2926 1632 2929 2128
rect 2934 1802 2937 2058
rect 2934 1462 2937 1798
rect 2942 1632 2945 1708
rect 2950 1662 2953 2128
rect 2958 1752 2961 1958
rect 2958 1532 2961 1738
rect 2966 1692 2969 2178
rect 2918 1382 2921 1408
rect 2902 672 2905 708
rect 2910 482 2913 698
rect 2918 692 2921 1378
rect 2930 1328 2934 1331
rect 2942 1252 2945 1528
rect 2950 1271 2953 1368
rect 2950 1268 2958 1271
rect 2930 1148 2934 1151
rect 2966 1052 2969 1658
rect 2974 952 2977 2688
rect 2982 2122 2985 2548
rect 2990 2332 2993 3098
rect 2998 2372 3001 3148
rect 3006 3082 3009 3418
rect 3022 3272 3025 3588
rect 3038 3582 3041 3758
rect 3046 3662 3049 3868
rect 3038 3432 3041 3578
rect 3030 3141 3033 3328
rect 3054 3302 3057 4548
rect 3078 4232 3081 4538
rect 3086 4512 3089 4628
rect 3096 4503 3098 4507
rect 3102 4503 3105 4507
rect 3110 4503 3112 4507
rect 3096 4303 3098 4307
rect 3102 4303 3105 4307
rect 3110 4303 3112 4307
rect 3126 4152 3129 4288
rect 3134 4212 3137 4458
rect 3198 4442 3201 4468
rect 3262 4462 3265 4548
rect 3382 4512 3385 4698
rect 3406 4482 3409 4648
rect 3486 4552 3489 4618
rect 3490 4548 3494 4551
rect 3150 4402 3153 4418
rect 3198 4412 3201 4438
rect 3150 4322 3153 4348
rect 3174 4342 3177 4348
rect 3150 4272 3153 4318
rect 3142 4242 3145 4258
rect 3096 4103 3098 4107
rect 3102 4103 3105 4107
rect 3110 4103 3112 4107
rect 3070 3872 3073 4048
rect 3070 3822 3073 3868
rect 3078 3862 3081 3908
rect 3096 3903 3098 3907
rect 3102 3903 3105 3907
rect 3110 3903 3112 3907
rect 3086 3702 3089 3748
rect 3096 3703 3098 3707
rect 3102 3703 3105 3707
rect 3110 3703 3112 3707
rect 3086 3551 3089 3688
rect 3118 3672 3121 3678
rect 3126 3592 3129 4128
rect 3134 3922 3137 4188
rect 3134 3592 3137 3918
rect 3150 3602 3153 4248
rect 3182 4072 3185 4258
rect 3198 4062 3201 4088
rect 3082 3548 3089 3551
rect 3096 3503 3098 3507
rect 3102 3503 3105 3507
rect 3110 3503 3112 3507
rect 3106 3478 3110 3481
rect 3070 3438 3078 3441
rect 3062 3262 3065 3328
rect 3062 3192 3065 3258
rect 3030 3138 3038 3141
rect 3030 3112 3033 3138
rect 3030 2982 3033 3108
rect 3046 3081 3049 3118
rect 3042 3078 3049 3081
rect 3022 2922 3025 2968
rect 3018 2848 3022 2851
rect 3046 2842 3049 3068
rect 3070 2912 3073 3438
rect 3078 3312 3081 3328
rect 3086 3302 3089 3358
rect 3096 3303 3098 3307
rect 3102 3303 3105 3307
rect 3110 3303 3112 3307
rect 3078 3052 3081 3088
rect 3086 2822 3089 3198
rect 3096 3103 3098 3107
rect 3102 3103 3105 3107
rect 3110 3103 3112 3107
rect 3110 2932 3113 2938
rect 3096 2903 3098 2907
rect 3102 2903 3105 2907
rect 3110 2903 3112 2907
rect 3118 2902 3121 3188
rect 3126 2952 3129 3558
rect 3134 3352 3137 3528
rect 3182 3462 3185 3568
rect 3206 3552 3209 4398
rect 3214 4292 3217 4398
rect 3214 4112 3217 4148
rect 3222 4092 3225 4278
rect 3238 4142 3241 4418
rect 3510 4412 3513 4698
rect 3678 4672 3681 4868
rect 4138 4838 4145 4841
rect 3874 4718 3881 4721
rect 3578 4668 3585 4671
rect 3554 4658 3558 4661
rect 3526 4522 3529 4538
rect 3538 4528 3542 4531
rect 3518 4472 3521 4488
rect 3214 3852 3217 3978
rect 3222 3722 3225 4078
rect 3230 4062 3233 4078
rect 3238 3852 3241 4078
rect 3214 3572 3217 3718
rect 3186 3458 3193 3461
rect 3150 3452 3153 3458
rect 3146 3318 3150 3321
rect 3142 3132 3145 3298
rect 3038 2762 3041 2768
rect 3006 2712 3009 2728
rect 3038 2662 3041 2758
rect 3054 2682 3057 2708
rect 3046 2678 3054 2681
rect 3006 2522 3009 2528
rect 3006 2492 3009 2498
rect 2994 2278 2998 2281
rect 2998 2171 3001 2178
rect 2994 2168 3001 2171
rect 2982 1972 2985 2118
rect 2998 2102 3001 2108
rect 2982 1942 2985 1948
rect 3006 1941 3009 2458
rect 3014 2222 3017 2568
rect 3022 2462 3025 2468
rect 3022 2172 3025 2228
rect 3014 2092 3017 2118
rect 2998 1938 3009 1941
rect 2982 1752 2985 1938
rect 2998 1772 3001 1938
rect 3006 1912 3009 1928
rect 2982 1592 2985 1748
rect 2982 1292 2985 1498
rect 2990 1082 2993 1768
rect 2998 1602 3001 1748
rect 3006 1582 3009 1598
rect 2998 1392 3001 1538
rect 3006 1352 3009 1538
rect 3014 1442 3017 1968
rect 3022 1682 3025 2168
rect 3030 1882 3033 2408
rect 3046 2272 3049 2678
rect 3062 2492 3065 2798
rect 3070 2702 3073 2718
rect 3058 2468 3065 2471
rect 3038 2142 3041 2158
rect 3046 2142 3049 2238
rect 3054 2152 3057 2338
rect 3062 2322 3065 2468
rect 3070 2312 3073 2688
rect 3078 2682 3081 2698
rect 3086 2652 3089 2818
rect 3102 2782 3105 2858
rect 3114 2848 3118 2851
rect 3126 2732 3129 2788
rect 3118 2712 3121 2728
rect 3096 2703 3098 2707
rect 3102 2703 3105 2707
rect 3110 2703 3112 2707
rect 3118 2682 3121 2698
rect 3130 2618 3134 2621
rect 3086 2532 3089 2608
rect 3038 2062 3041 2098
rect 3030 1752 3033 1808
rect 3030 1708 3038 1711
rect 3030 1652 3033 1708
rect 3022 1392 3025 1538
rect 3022 1182 3025 1318
rect 2970 928 2977 931
rect 2974 922 2977 928
rect 2950 872 2953 878
rect 2950 802 2953 868
rect 2926 652 2929 658
rect 2934 522 2937 668
rect 2950 362 2953 748
rect 2966 582 2969 818
rect 2970 578 2974 581
rect 2870 262 2873 298
rect 2958 262 2961 548
rect 2966 472 2969 558
rect 2990 522 2993 588
rect 2998 532 3001 1168
rect 3006 872 3009 1078
rect 3030 1022 3033 1558
rect 3038 1472 3041 1528
rect 3046 1471 3049 2138
rect 3054 2122 3057 2128
rect 3054 1552 3057 1768
rect 3062 1752 3065 2238
rect 3070 1752 3073 2308
rect 3078 2262 3081 2488
rect 3078 2142 3081 2258
rect 3078 1912 3081 2118
rect 3086 2022 3089 2528
rect 3096 2503 3098 2507
rect 3102 2503 3105 2507
rect 3110 2503 3112 2507
rect 3118 2432 3121 2508
rect 3134 2502 3137 2578
rect 3142 2522 3145 2708
rect 3126 2422 3129 2428
rect 3134 2412 3137 2468
rect 3110 2372 3113 2408
rect 3096 2303 3098 2307
rect 3102 2303 3105 2307
rect 3110 2303 3112 2307
rect 3118 2272 3121 2368
rect 3102 2232 3105 2258
rect 3110 2162 3113 2218
rect 3096 2103 3098 2107
rect 3102 2103 3105 2107
rect 3110 2103 3112 2107
rect 3118 2052 3121 2228
rect 3126 2112 3129 2208
rect 3134 2122 3137 2328
rect 3126 2082 3129 2098
rect 3096 1903 3098 1907
rect 3102 1903 3105 1907
rect 3110 1903 3112 1907
rect 3082 1898 3086 1901
rect 3070 1622 3073 1718
rect 3054 1502 3057 1548
rect 3062 1532 3065 1538
rect 3046 1468 3054 1471
rect 3070 1422 3073 1608
rect 3078 1462 3081 1888
rect 3118 1862 3121 2038
rect 3142 1911 3145 2478
rect 3150 2462 3153 2918
rect 3158 2412 3161 2838
rect 3150 2192 3153 2298
rect 3158 2212 3161 2388
rect 3150 1922 3153 2108
rect 3166 2042 3169 2828
rect 3174 2732 3177 2858
rect 3174 2352 3177 2648
rect 3182 2471 3185 3098
rect 3190 3072 3193 3458
rect 3198 3262 3201 3268
rect 3190 2982 3193 2998
rect 3182 2468 3190 2471
rect 3182 2402 3185 2408
rect 3190 2362 3193 2458
rect 3198 2402 3201 2928
rect 3206 2812 3209 3368
rect 3238 2932 3241 3848
rect 3246 3672 3249 4148
rect 3254 4062 3257 4158
rect 3254 3702 3257 3948
rect 3246 3332 3249 3668
rect 3254 3662 3257 3668
rect 3246 3052 3249 3208
rect 3254 2852 3257 3338
rect 3262 3282 3265 3868
rect 3206 2572 3209 2698
rect 3214 2572 3217 2728
rect 3230 2602 3233 2608
rect 3206 2402 3209 2528
rect 3214 2482 3217 2488
rect 3174 2252 3177 2348
rect 3174 2062 3177 2248
rect 3198 2112 3201 2358
rect 3206 2042 3209 2398
rect 3230 2372 3233 2538
rect 3230 2281 3233 2368
rect 3238 2302 3241 2468
rect 3246 2362 3249 2788
rect 3254 2552 3257 2848
rect 3262 2702 3265 3268
rect 3270 3212 3273 4138
rect 3278 3982 3281 4258
rect 3278 2942 3281 3978
rect 3294 3862 3297 4218
rect 3286 2972 3289 3768
rect 3318 3742 3321 4338
rect 3326 4332 3329 4338
rect 3326 4052 3329 4298
rect 3342 3942 3345 4008
rect 3366 3872 3369 4378
rect 3478 4338 3486 4341
rect 3422 4222 3425 4328
rect 3430 4252 3433 4258
rect 3398 4112 3401 4178
rect 3406 4142 3409 4178
rect 3390 3922 3393 3928
rect 3366 3862 3369 3868
rect 3334 3832 3337 3858
rect 3342 3852 3345 3858
rect 3294 3482 3297 3498
rect 3278 2782 3281 2878
rect 3302 2832 3305 3548
rect 3310 3522 3313 3548
rect 3326 3462 3329 3658
rect 3342 3562 3345 3628
rect 3326 3302 3329 3458
rect 3350 3332 3353 3418
rect 3310 3092 3313 3298
rect 3358 3242 3361 3438
rect 3322 3228 3326 3231
rect 3310 2792 3313 3088
rect 3326 3062 3329 3068
rect 3342 3042 3345 3068
rect 3318 2922 3321 2938
rect 3326 2922 3329 2978
rect 3358 2952 3361 3118
rect 3334 2842 3337 2848
rect 3262 2462 3265 2638
rect 3286 2542 3289 2728
rect 3310 2592 3313 2678
rect 3254 2362 3257 2448
rect 3230 2278 3238 2281
rect 3214 2192 3217 2218
rect 3174 1922 3177 2028
rect 3222 1972 3225 2278
rect 3202 1968 3206 1971
rect 3142 1908 3150 1911
rect 3086 1692 3089 1718
rect 3096 1703 3098 1707
rect 3102 1703 3105 1707
rect 3110 1703 3112 1707
rect 3086 1672 3089 1678
rect 3094 1612 3097 1678
rect 3118 1612 3121 1858
rect 3126 1692 3129 1908
rect 3138 1898 3145 1901
rect 3142 1852 3145 1898
rect 3134 1642 3137 1678
rect 3096 1503 3098 1507
rect 3102 1503 3105 1507
rect 3110 1503 3112 1507
rect 3118 1492 3121 1588
rect 3142 1562 3145 1738
rect 3150 1532 3153 1908
rect 3182 1872 3185 1928
rect 3158 1792 3161 1858
rect 3166 1652 3169 1858
rect 3190 1832 3193 1858
rect 3174 1692 3177 1818
rect 3174 1572 3177 1638
rect 3126 1422 3129 1448
rect 3038 1262 3041 1278
rect 3070 1052 3073 1078
rect 3078 1072 3081 1098
rect 3030 942 3033 1018
rect 2998 492 3001 528
rect 2986 338 2990 341
rect 2862 162 2865 218
rect 2854 142 2857 158
rect 2686 72 2689 78
rect 2374 62 2377 68
rect 2282 58 2286 61
rect 2754 58 2758 61
rect 2822 52 2825 108
rect 2998 92 3001 408
rect 3006 392 3009 668
rect 3014 592 3017 628
rect 3022 372 3025 728
rect 3022 282 3025 368
rect 3030 222 3033 898
rect 3062 672 3065 988
rect 3078 912 3081 1008
rect 3070 752 3073 778
rect 3070 742 3073 748
rect 3086 702 3089 1398
rect 3102 1352 3105 1418
rect 3110 1332 3113 1418
rect 3134 1332 3137 1498
rect 3142 1472 3145 1488
rect 3150 1421 3153 1528
rect 3150 1418 3158 1421
rect 3166 1352 3169 1568
rect 3182 1492 3185 1828
rect 3190 1732 3193 1748
rect 3186 1468 3190 1471
rect 3096 1303 3098 1307
rect 3102 1303 3105 1307
rect 3110 1303 3112 1307
rect 3110 1152 3113 1238
rect 3126 1122 3129 1138
rect 3096 1103 3098 1107
rect 3102 1103 3105 1107
rect 3110 1103 3112 1107
rect 3134 1082 3137 1298
rect 3150 1252 3153 1288
rect 3166 1282 3169 1308
rect 3158 1242 3161 1268
rect 3182 1262 3185 1278
rect 3150 1112 3153 1208
rect 3096 903 3098 907
rect 3102 903 3105 907
rect 3110 903 3112 907
rect 3098 718 3102 721
rect 3096 703 3098 707
rect 3102 703 3105 707
rect 3110 703 3112 707
rect 3062 662 3065 668
rect 3096 503 3098 507
rect 3102 503 3105 507
rect 3110 503 3112 507
rect 3118 392 3121 978
rect 3126 312 3129 958
rect 3142 932 3145 958
rect 3134 762 3137 768
rect 3150 712 3153 1108
rect 3158 762 3161 1228
rect 3174 1102 3177 1158
rect 3182 1082 3185 1168
rect 3134 432 3137 688
rect 3158 662 3161 668
rect 3166 662 3169 858
rect 3174 772 3177 848
rect 3182 792 3185 1048
rect 3182 552 3185 678
rect 3190 642 3193 1248
rect 3198 681 3201 1648
rect 3206 1462 3209 1678
rect 3214 1652 3217 1728
rect 3214 1532 3217 1538
rect 3206 1092 3209 1458
rect 3214 1342 3217 1488
rect 3214 1272 3217 1338
rect 3222 1312 3225 1498
rect 3230 1312 3233 1698
rect 3238 1532 3241 2118
rect 3246 2112 3249 2158
rect 3262 2052 3265 2058
rect 3262 1912 3265 2048
rect 3214 1192 3217 1228
rect 3206 912 3209 1088
rect 3206 732 3209 748
rect 3198 678 3209 681
rect 3198 662 3201 668
rect 3096 303 3098 307
rect 3102 303 3105 307
rect 3110 303 3112 307
rect 3174 252 3177 498
rect 3206 152 3209 678
rect 3214 672 3217 798
rect 3096 103 3098 107
rect 3102 103 3105 107
rect 3110 103 3112 107
rect 2650 48 2654 51
rect 3222 12 3225 1268
rect 3230 742 3233 1158
rect 3238 1002 3241 1498
rect 3246 1332 3249 1548
rect 3254 1422 3257 1868
rect 3262 1741 3265 1898
rect 3270 1752 3273 2158
rect 3262 1738 3273 1741
rect 3250 1318 3254 1321
rect 3246 1292 3249 1298
rect 3238 852 3241 888
rect 3246 762 3249 888
rect 3254 652 3257 1258
rect 3262 862 3265 1688
rect 3270 982 3273 1738
rect 3278 1722 3281 2318
rect 3286 2232 3289 2538
rect 3302 2452 3305 2458
rect 3302 2402 3305 2438
rect 3302 2351 3305 2388
rect 3310 2372 3313 2498
rect 3318 2472 3321 2638
rect 3298 2348 3305 2351
rect 3286 2162 3289 2198
rect 3302 2122 3305 2208
rect 3310 2202 3313 2348
rect 3318 2312 3321 2338
rect 3326 2272 3329 2818
rect 3334 2552 3337 2558
rect 3334 2282 3337 2518
rect 3342 2422 3345 2838
rect 3350 2752 3353 2868
rect 3358 2812 3361 2948
rect 3350 2682 3353 2748
rect 3350 2602 3353 2648
rect 3354 2558 3358 2561
rect 3366 2502 3369 3768
rect 3374 3762 3377 3908
rect 3382 3842 3385 3868
rect 3398 3832 3401 4008
rect 3414 3932 3417 4058
rect 3394 3698 3401 3701
rect 3390 3672 3393 3688
rect 3382 3512 3385 3518
rect 3382 3402 3385 3508
rect 3390 3192 3393 3448
rect 3398 3312 3401 3698
rect 3406 3622 3409 3748
rect 3406 3532 3409 3578
rect 3374 3152 3377 3158
rect 3398 2862 3401 3298
rect 3390 2802 3393 2858
rect 3382 2542 3385 2548
rect 3358 2488 3366 2491
rect 3350 2422 3353 2438
rect 3358 2362 3361 2488
rect 3286 2102 3289 2108
rect 3278 1652 3281 1658
rect 3278 1192 3281 1638
rect 3286 1392 3289 2018
rect 3294 1362 3297 2048
rect 3302 1942 3305 1948
rect 3286 1172 3289 1248
rect 3294 1212 3297 1318
rect 3302 1212 3305 1688
rect 3310 1302 3313 2198
rect 3318 2042 3321 2118
rect 3326 2052 3329 2268
rect 3342 2162 3345 2298
rect 3374 2272 3377 2518
rect 3382 2492 3385 2508
rect 3390 2462 3393 2748
rect 3406 2712 3409 2998
rect 3414 2842 3417 3928
rect 3422 3672 3425 4218
rect 3430 4112 3433 4148
rect 3434 3878 3438 3881
rect 3430 3471 3433 3618
rect 3438 3532 3441 3718
rect 3446 3672 3449 4068
rect 3446 3662 3449 3668
rect 3454 3662 3457 3968
rect 3462 3942 3465 4308
rect 3470 4092 3473 4288
rect 3478 4162 3481 4338
rect 3470 4002 3473 4038
rect 3478 3862 3481 4128
rect 3486 4042 3489 4058
rect 3450 3648 3457 3651
rect 3454 3642 3457 3648
rect 3426 3468 3433 3471
rect 3446 3212 3449 3438
rect 3454 3282 3457 3538
rect 3462 3262 3465 3688
rect 3478 3542 3481 3588
rect 3470 3262 3473 3488
rect 3478 3462 3481 3488
rect 3470 3248 3478 3251
rect 3406 2442 3409 2458
rect 3422 2442 3425 3178
rect 3470 3172 3473 3248
rect 3486 3241 3489 4008
rect 3494 3842 3497 4368
rect 3526 4292 3529 4508
rect 3534 4488 3542 4491
rect 3534 4482 3537 4488
rect 3502 4022 3505 4118
rect 3526 4092 3529 4178
rect 3494 3571 3497 3828
rect 3510 3592 3513 4068
rect 3518 3762 3521 3968
rect 3534 3962 3537 4258
rect 3542 3872 3545 4178
rect 3550 4102 3553 4508
rect 3558 4362 3561 4658
rect 3558 4152 3561 4278
rect 3566 4132 3569 4438
rect 3582 4112 3585 4668
rect 3608 4603 3610 4607
rect 3614 4603 3617 4607
rect 3622 4603 3624 4607
rect 3558 4072 3561 4108
rect 3522 3728 3526 3731
rect 3542 3662 3545 3728
rect 3494 3568 3502 3571
rect 3494 3352 3497 3458
rect 3518 3392 3521 3658
rect 3542 3602 3545 3638
rect 3518 3362 3521 3388
rect 3494 3332 3497 3338
rect 3478 3238 3489 3241
rect 3466 3138 3470 3141
rect 3430 3112 3433 3138
rect 3446 3132 3449 3138
rect 3430 2492 3433 2498
rect 3382 2362 3385 2438
rect 3414 2422 3417 2438
rect 3422 2422 3425 2428
rect 3438 2392 3441 3058
rect 3454 2562 3457 2728
rect 3462 2542 3465 3128
rect 3454 2531 3457 2538
rect 3454 2528 3462 2531
rect 3462 2462 3465 2508
rect 3470 2452 3473 3048
rect 3478 2772 3481 3238
rect 3518 3052 3521 3258
rect 3526 3062 3529 3068
rect 3478 2622 3481 2638
rect 3478 2432 3481 2528
rect 3446 2412 3449 2418
rect 3362 2238 3366 2241
rect 3350 2142 3353 2148
rect 3398 2062 3401 2348
rect 3414 2332 3417 2348
rect 3422 2322 3425 2348
rect 3414 2222 3417 2258
rect 3422 2232 3425 2318
rect 3438 2308 3446 2311
rect 3414 2072 3417 2088
rect 3422 2042 3425 2138
rect 3430 2062 3433 2068
rect 3342 2002 3345 2008
rect 3326 1852 3329 1958
rect 3350 1932 3353 1998
rect 3358 1962 3361 2008
rect 3358 1942 3361 1958
rect 3382 1941 3385 1948
rect 3382 1938 3390 1941
rect 3318 1492 3321 1618
rect 3322 1338 3326 1341
rect 3306 1188 3310 1191
rect 3294 1142 3297 1158
rect 3278 872 3281 938
rect 3294 912 3297 958
rect 3270 852 3273 858
rect 3278 842 3281 868
rect 3294 862 3297 908
rect 3262 752 3265 758
rect 3254 542 3257 638
rect 3254 342 3257 538
rect 3294 392 3297 748
rect 3302 492 3305 868
rect 3310 542 3313 1058
rect 3318 662 3321 1148
rect 3334 1072 3337 1608
rect 3342 1581 3345 1638
rect 3342 1578 3350 1581
rect 3342 1532 3345 1538
rect 3350 1532 3353 1538
rect 3350 1452 3353 1528
rect 3358 1292 3361 1358
rect 3342 1152 3345 1188
rect 3342 1042 3345 1068
rect 3358 922 3361 1198
rect 3366 1162 3369 1888
rect 3374 1842 3377 1938
rect 3414 1892 3417 1978
rect 3430 1962 3433 1998
rect 3422 1948 3430 1951
rect 3422 1942 3425 1948
rect 3430 1932 3433 1948
rect 3374 1662 3377 1838
rect 3382 1782 3385 1808
rect 3406 1762 3409 1848
rect 3406 1752 3409 1758
rect 3386 1718 3393 1721
rect 3382 1662 3385 1668
rect 3390 1382 3393 1718
rect 3414 1692 3417 1888
rect 3414 1582 3417 1618
rect 3374 1202 3377 1238
rect 3382 1172 3385 1368
rect 3366 1042 3369 1058
rect 3382 1042 3385 1148
rect 3374 872 3377 948
rect 3346 868 3350 871
rect 3378 868 3385 871
rect 3382 862 3385 868
rect 3342 858 3350 861
rect 3342 542 3345 858
rect 3362 738 3366 741
rect 3310 462 3313 538
rect 3294 292 3297 388
rect 3310 352 3313 458
rect 3310 262 3313 348
rect 3334 332 3337 368
rect 3326 192 3329 328
rect 3366 272 3369 338
rect 3398 182 3401 1278
rect 3406 482 3409 1418
rect 3422 1412 3425 1818
rect 3430 1412 3433 1648
rect 3438 1472 3441 2308
rect 3454 2122 3457 2328
rect 3470 2222 3473 2358
rect 3478 2302 3481 2308
rect 3462 2212 3465 2218
rect 3474 2198 3481 2201
rect 3478 2132 3481 2198
rect 3486 2112 3489 2418
rect 3494 2392 3497 2978
rect 3502 2792 3505 2988
rect 3510 2862 3513 3028
rect 3518 3012 3521 3038
rect 3526 2862 3529 3048
rect 3502 2392 3505 2748
rect 3494 2302 3497 2368
rect 3502 2082 3505 2338
rect 3510 2242 3513 2858
rect 3534 2752 3537 3468
rect 3542 3252 3545 3598
rect 3550 3312 3553 4058
rect 3566 3852 3569 3988
rect 3558 3432 3561 3798
rect 3550 2992 3553 3268
rect 3558 3252 3561 3278
rect 3550 2852 3553 2968
rect 3566 2842 3569 3848
rect 3574 3582 3577 4098
rect 3590 3762 3593 4538
rect 3608 4403 3610 4407
rect 3614 4403 3617 4407
rect 3622 4403 3624 4407
rect 3646 4392 3649 4658
rect 3678 4542 3681 4668
rect 3630 4248 3638 4251
rect 3598 4232 3601 4248
rect 3608 4203 3610 4207
rect 3614 4203 3617 4207
rect 3622 4203 3624 4207
rect 3598 4152 3601 4198
rect 3630 4192 3633 4248
rect 3582 3732 3585 3748
rect 3582 3532 3585 3728
rect 3590 3612 3593 3638
rect 3578 3418 3582 3421
rect 3590 3202 3593 3228
rect 3574 2932 3577 3128
rect 3558 2772 3561 2818
rect 3518 2532 3521 2718
rect 3534 2682 3537 2748
rect 3526 2522 3529 2568
rect 3526 2462 3529 2468
rect 3518 2322 3521 2338
rect 3510 2192 3513 2198
rect 3450 2068 3454 2071
rect 3462 2002 3465 2078
rect 3518 2072 3521 2308
rect 3526 2302 3529 2338
rect 3534 2152 3537 2578
rect 3470 2032 3473 2058
rect 3446 1822 3449 1848
rect 3446 1552 3449 1818
rect 3454 1762 3457 1998
rect 3462 1732 3465 1958
rect 3478 1882 3481 2038
rect 3486 1902 3489 2048
rect 3414 1282 3417 1378
rect 3438 1292 3441 1468
rect 3446 1302 3449 1438
rect 3454 1402 3457 1698
rect 3470 1592 3473 1848
rect 3454 1392 3457 1398
rect 3454 1252 3457 1288
rect 3462 1212 3465 1468
rect 3438 1051 3441 1068
rect 3438 1048 3446 1051
rect 3454 1041 3457 1198
rect 3462 1052 3465 1068
rect 3446 1038 3457 1041
rect 3418 958 3422 961
rect 3414 512 3417 938
rect 3422 532 3425 548
rect 3430 472 3433 888
rect 3438 842 3441 858
rect 3446 832 3449 1038
rect 3470 972 3473 1588
rect 3486 1462 3489 1868
rect 3494 1862 3497 1898
rect 3494 1732 3497 1848
rect 3502 1732 3505 1758
rect 3494 1672 3497 1728
rect 3510 1702 3513 2068
rect 3518 1712 3521 2068
rect 3526 1932 3529 2138
rect 3534 2092 3537 2138
rect 3534 1742 3537 1938
rect 3542 1812 3545 2648
rect 3550 2632 3553 2748
rect 3566 2662 3569 2828
rect 3550 2332 3553 2618
rect 3558 2352 3561 2568
rect 3566 2342 3569 2638
rect 3574 2632 3577 2878
rect 3582 2702 3585 2898
rect 3598 2842 3601 4138
rect 3608 4003 3610 4007
rect 3614 4003 3617 4007
rect 3622 4003 3624 4007
rect 3614 3871 3617 3988
rect 3610 3868 3617 3871
rect 3614 3822 3617 3868
rect 3630 3942 3633 4058
rect 3638 4042 3641 4158
rect 3608 3803 3610 3807
rect 3614 3803 3617 3807
rect 3622 3803 3624 3807
rect 3608 3603 3610 3607
rect 3614 3603 3617 3607
rect 3622 3603 3624 3607
rect 3608 3403 3610 3407
rect 3614 3403 3617 3407
rect 3622 3403 3624 3407
rect 3622 3332 3625 3348
rect 3608 3203 3610 3207
rect 3614 3203 3617 3207
rect 3622 3203 3624 3207
rect 3608 3003 3610 3007
rect 3614 3003 3617 3007
rect 3622 3003 3624 3007
rect 3606 2952 3609 2958
rect 3614 2862 3617 2968
rect 3630 2892 3633 3938
rect 3638 3762 3641 4038
rect 3670 4032 3673 4348
rect 3642 3688 3646 3691
rect 3654 3442 3657 3848
rect 3662 3742 3665 3968
rect 3670 3792 3673 4018
rect 3678 3892 3681 4538
rect 3710 4162 3713 4388
rect 3750 4382 3753 4618
rect 3798 4468 3806 4471
rect 3670 3742 3673 3788
rect 3662 3562 3665 3738
rect 3662 3452 3665 3468
rect 3638 2942 3641 3378
rect 3608 2803 3610 2807
rect 3614 2803 3617 2807
rect 3622 2803 3624 2807
rect 3614 2772 3617 2788
rect 3586 2658 3590 2661
rect 3562 2298 3569 2301
rect 3566 2292 3569 2298
rect 3574 2232 3577 2548
rect 3582 2492 3585 2528
rect 3590 2422 3593 2578
rect 3598 2352 3601 2758
rect 3630 2732 3633 2888
rect 3646 2822 3649 3278
rect 3654 2912 3657 3298
rect 3662 3272 3665 3408
rect 3678 3272 3681 3848
rect 3686 3652 3689 4008
rect 3694 3651 3697 3858
rect 3710 3802 3713 4158
rect 3718 3892 3721 4238
rect 3726 4062 3729 4148
rect 3742 4141 3745 4248
rect 3742 4138 3750 4141
rect 3742 4042 3745 4078
rect 3758 4072 3761 4368
rect 3770 4338 3774 4341
rect 3782 4272 3785 4348
rect 3790 4241 3793 4278
rect 3798 4261 3801 4468
rect 3798 4258 3806 4261
rect 3790 4238 3798 4241
rect 3790 4232 3793 4238
rect 3814 4202 3817 4568
rect 3862 4462 3865 4638
rect 3878 4592 3881 4718
rect 4046 4642 4049 4818
rect 3886 4442 3889 4518
rect 3822 4412 3825 4438
rect 3774 4198 3782 4201
rect 3750 3982 3753 4018
rect 3702 3682 3705 3748
rect 3694 3648 3702 3651
rect 3662 2942 3665 2948
rect 3608 2603 3610 2607
rect 3614 2603 3617 2607
rect 3622 2603 3624 2607
rect 3630 2602 3633 2618
rect 3606 2422 3609 2588
rect 3626 2548 3630 2551
rect 3614 2452 3617 2538
rect 3622 2462 3625 2478
rect 3614 2422 3617 2438
rect 3608 2403 3610 2407
rect 3614 2403 3617 2407
rect 3622 2403 3624 2407
rect 3614 2282 3617 2308
rect 3622 2241 3625 2368
rect 3630 2252 3633 2258
rect 3622 2238 3633 2241
rect 3574 2208 3582 2211
rect 3542 1752 3545 1808
rect 3550 1772 3553 2178
rect 3558 2162 3561 2188
rect 3566 2082 3569 2158
rect 3574 2012 3577 2208
rect 3582 2122 3585 2168
rect 3598 2152 3601 2228
rect 3608 2203 3610 2207
rect 3614 2203 3617 2207
rect 3622 2203 3624 2207
rect 3630 2202 3633 2238
rect 3630 2162 3633 2198
rect 3562 1948 3566 1951
rect 3574 1902 3577 1958
rect 3582 1872 3585 2058
rect 3598 2012 3601 2128
rect 3608 2003 3610 2007
rect 3614 2003 3617 2007
rect 3622 2003 3624 2007
rect 3598 1908 3606 1911
rect 3582 1762 3585 1808
rect 3608 1803 3610 1807
rect 3614 1803 3617 1807
rect 3622 1803 3624 1807
rect 3486 1072 3489 1078
rect 3438 542 3441 768
rect 3454 542 3457 828
rect 3470 562 3473 928
rect 3494 702 3497 1128
rect 3502 1072 3505 1658
rect 3518 1262 3521 1708
rect 3534 1532 3537 1738
rect 3562 1638 3566 1641
rect 3526 1242 3529 1248
rect 3510 1148 3518 1151
rect 3510 1012 3513 1148
rect 3518 1122 3521 1128
rect 3526 952 3529 1148
rect 3502 888 3510 891
rect 3502 642 3505 888
rect 3518 782 3521 798
rect 3522 648 3529 651
rect 3450 538 3454 541
rect 3438 442 3441 538
rect 3454 382 3457 508
rect 3470 402 3473 558
rect 3518 552 3521 628
rect 3526 522 3529 648
rect 3534 562 3537 1358
rect 3542 832 3545 1548
rect 3574 1502 3577 1758
rect 3598 1752 3601 1788
rect 3630 1652 3633 1878
rect 3598 1602 3601 1618
rect 3608 1603 3610 1607
rect 3614 1603 3617 1607
rect 3622 1603 3624 1607
rect 3622 1562 3625 1568
rect 3630 1562 3633 1598
rect 3558 1222 3561 1258
rect 3558 1042 3561 1118
rect 3542 812 3545 828
rect 3566 612 3569 1458
rect 3558 552 3561 558
rect 3462 242 3465 348
rect 3478 282 3481 508
rect 3490 148 3494 151
rect 3310 82 3313 148
rect 3410 138 3414 141
rect 3566 132 3569 588
rect 3574 562 3577 1448
rect 3582 572 3585 1538
rect 3590 1492 3593 1528
rect 3590 1101 3593 1488
rect 3608 1403 3610 1407
rect 3614 1403 3617 1407
rect 3622 1403 3624 1407
rect 3630 1372 3633 1458
rect 3618 1328 3622 1331
rect 3622 1262 3625 1268
rect 3630 1242 3633 1368
rect 3608 1203 3610 1207
rect 3614 1203 3617 1207
rect 3622 1203 3624 1207
rect 3638 1192 3641 2418
rect 3646 2102 3649 2728
rect 3654 2152 3657 2158
rect 3646 1822 3649 1828
rect 3654 1752 3657 2138
rect 3662 2072 3665 2688
rect 3670 2502 3673 3268
rect 3678 2892 3681 3208
rect 3686 3102 3689 3648
rect 3694 3202 3697 3528
rect 3694 3172 3697 3198
rect 3678 2852 3681 2878
rect 3678 2662 3681 2808
rect 3686 2722 3689 3078
rect 3702 2762 3705 3648
rect 3710 3362 3713 3798
rect 3718 3751 3721 3818
rect 3734 3752 3737 3778
rect 3718 3748 3726 3751
rect 3718 3682 3721 3688
rect 3734 3672 3737 3678
rect 3718 3252 3721 3578
rect 3750 3561 3753 3868
rect 3746 3558 3753 3561
rect 3742 3452 3745 3558
rect 3742 3351 3745 3448
rect 3738 3348 3745 3351
rect 3726 3282 3729 3348
rect 3710 2962 3713 2988
rect 3718 2962 3721 3218
rect 3726 3082 3729 3278
rect 3734 3272 3737 3348
rect 3742 3322 3745 3328
rect 3750 3142 3753 3528
rect 3758 3252 3761 4058
rect 3766 3962 3769 4128
rect 3774 3852 3777 4198
rect 3766 3632 3769 3638
rect 3766 3482 3769 3498
rect 3774 3292 3777 3848
rect 3782 3542 3785 4068
rect 3790 4052 3793 4058
rect 3790 3502 3793 4048
rect 3806 4032 3809 4058
rect 3738 3128 3745 3131
rect 3718 2842 3721 2948
rect 3726 2732 3729 3008
rect 3742 2732 3745 3128
rect 3762 2998 3769 3001
rect 3750 2902 3753 2948
rect 3766 2922 3769 2998
rect 3762 2848 3766 2851
rect 3750 2812 3753 2848
rect 3774 2832 3777 2958
rect 3782 2892 3785 3438
rect 3798 3382 3801 3728
rect 3814 3602 3817 3778
rect 3814 3512 3817 3528
rect 3810 3508 3814 3511
rect 3822 3482 3825 4178
rect 3846 3962 3849 4328
rect 3886 4302 3889 4438
rect 3870 4262 3873 4268
rect 3830 3928 3838 3931
rect 3830 3642 3833 3928
rect 3790 2902 3793 3208
rect 3830 3172 3833 3588
rect 3838 3342 3841 3598
rect 3838 3142 3841 3338
rect 3806 3082 3809 3118
rect 3822 3052 3825 3088
rect 3830 3082 3833 3088
rect 3838 3072 3841 3138
rect 3838 3042 3841 3068
rect 3766 2792 3769 2798
rect 3782 2742 3785 2788
rect 3726 2712 3729 2728
rect 3686 2672 3689 2678
rect 3670 2242 3673 2458
rect 3662 1952 3665 2068
rect 3678 2032 3681 2638
rect 3686 2562 3689 2668
rect 3694 2652 3697 2698
rect 3686 2302 3689 2558
rect 3694 2422 3697 2648
rect 3702 2482 3705 2488
rect 3670 1841 3673 1948
rect 3662 1838 3673 1841
rect 3678 1842 3681 1938
rect 3646 1582 3649 1748
rect 3638 1162 3641 1188
rect 3590 1098 3598 1101
rect 3608 1003 3610 1007
rect 3614 1003 3617 1007
rect 3622 1003 3624 1007
rect 3630 812 3633 978
rect 3608 803 3610 807
rect 3614 803 3617 807
rect 3622 803 3624 807
rect 3608 603 3610 607
rect 3614 603 3617 607
rect 3622 603 3624 607
rect 3646 572 3649 1518
rect 3654 1362 3657 1688
rect 3662 1352 3665 1838
rect 3678 1782 3681 1798
rect 3670 1352 3673 1578
rect 3678 1272 3681 1778
rect 3686 1762 3689 2298
rect 3694 2172 3697 2338
rect 3694 2152 3697 2158
rect 3694 1812 3697 1858
rect 3686 1532 3689 1668
rect 3678 1152 3681 1178
rect 3670 1091 3673 1098
rect 3666 1088 3673 1091
rect 3574 492 3577 548
rect 3582 532 3585 568
rect 3646 522 3649 568
rect 3608 403 3610 407
rect 3614 403 3617 407
rect 3622 403 3624 407
rect 3646 372 3649 398
rect 3654 212 3657 1078
rect 3662 312 3665 548
rect 3678 402 3681 1118
rect 3686 512 3689 1488
rect 3702 1232 3705 2448
rect 3718 2442 3721 2468
rect 3710 2222 3713 2248
rect 3710 1612 3713 2108
rect 3718 1672 3721 2248
rect 3726 1992 3729 2338
rect 3734 2232 3737 2238
rect 3742 2212 3745 2608
rect 3750 2502 3753 2558
rect 3766 2432 3769 2438
rect 3750 2262 3753 2368
rect 3758 2302 3761 2328
rect 3750 2192 3753 2258
rect 3758 2242 3761 2288
rect 3742 2152 3745 2178
rect 3758 2162 3761 2188
rect 3718 1452 3721 1538
rect 3734 1492 3737 2118
rect 3766 2022 3769 2358
rect 3774 2182 3777 2268
rect 3782 2262 3785 2618
rect 3790 2612 3793 2858
rect 3798 2742 3801 2928
rect 3806 2802 3809 2838
rect 3806 2732 3809 2748
rect 3806 2682 3809 2718
rect 3806 2472 3809 2528
rect 3790 2442 3793 2458
rect 3790 2382 3793 2418
rect 3806 2402 3809 2468
rect 3798 2388 3806 2391
rect 3798 2382 3801 2388
rect 3806 2362 3809 2368
rect 3814 2352 3817 2528
rect 3758 1962 3761 2008
rect 3758 1802 3761 1958
rect 3774 1812 3777 1978
rect 3782 1952 3785 2248
rect 3806 2222 3809 2238
rect 3782 1862 3785 1948
rect 3790 1932 3793 2018
rect 3758 1772 3761 1798
rect 3742 1692 3745 1768
rect 3750 1582 3753 1718
rect 3758 1602 3761 1708
rect 3766 1702 3769 1718
rect 3770 1648 3777 1651
rect 3774 1642 3777 1648
rect 3694 842 3697 1098
rect 3710 902 3713 1318
rect 3742 1271 3745 1388
rect 3738 1268 3745 1271
rect 3722 1248 3729 1251
rect 3726 1242 3729 1248
rect 3750 1152 3753 1228
rect 3746 1118 3753 1121
rect 3734 1058 3742 1061
rect 3734 872 3737 1058
rect 3750 1042 3753 1118
rect 3758 1062 3761 1348
rect 3766 1082 3769 1358
rect 3782 1171 3785 1858
rect 3790 1722 3793 1928
rect 3798 1782 3801 1878
rect 3794 1688 3798 1691
rect 3790 1568 3798 1571
rect 3790 1252 3793 1568
rect 3806 1361 3809 2218
rect 3822 2192 3825 2768
rect 3830 2752 3833 2918
rect 3838 2882 3841 3008
rect 3846 2902 3849 3688
rect 3854 2982 3857 3928
rect 3870 3762 3873 4248
rect 3878 4022 3881 4268
rect 3886 3772 3889 4238
rect 3894 3922 3897 4528
rect 3970 4498 3977 4501
rect 3902 4242 3905 4458
rect 3918 4272 3921 4458
rect 3942 4341 3945 4348
rect 3938 4338 3945 4341
rect 3934 4302 3937 4338
rect 3902 4122 3905 4238
rect 3918 3972 3921 4268
rect 3942 4252 3945 4268
rect 3934 3942 3937 4108
rect 3942 4082 3945 4248
rect 3950 4092 3953 4488
rect 3958 4332 3961 4348
rect 3946 4058 3950 4061
rect 3862 3391 3865 3738
rect 3870 3652 3873 3758
rect 3878 3652 3881 3658
rect 3894 3482 3897 3818
rect 3902 3752 3905 3758
rect 3890 3468 3894 3471
rect 3862 3388 3873 3391
rect 3854 2921 3857 2978
rect 3862 2932 3865 3378
rect 3870 2932 3873 3388
rect 3894 3232 3897 3238
rect 3902 3132 3905 3748
rect 3910 3512 3913 3548
rect 3918 3442 3921 3558
rect 3910 3322 3913 3328
rect 3854 2918 3865 2921
rect 3846 2852 3849 2858
rect 3854 2762 3857 2878
rect 3862 2762 3865 2918
rect 3830 2362 3833 2748
rect 3838 2562 3841 2718
rect 3846 2542 3849 2648
rect 3830 2342 3833 2348
rect 3822 1902 3825 2168
rect 3818 1878 3822 1881
rect 3814 1742 3817 1748
rect 3814 1552 3817 1708
rect 3822 1682 3825 1748
rect 3802 1358 3809 1361
rect 3814 1372 3817 1438
rect 3814 1312 3817 1368
rect 3830 1352 3833 1748
rect 3838 1662 3841 1928
rect 3846 1672 3849 2358
rect 3854 2252 3857 2758
rect 3862 2512 3865 2528
rect 3862 2452 3865 2458
rect 3870 2342 3873 2868
rect 3878 2772 3881 3118
rect 3918 3082 3921 3408
rect 3926 3332 3929 3688
rect 3934 3352 3937 3738
rect 3942 3642 3945 3848
rect 3926 3162 3929 3328
rect 3934 3151 3937 3348
rect 3926 3148 3937 3151
rect 3914 3068 3918 3071
rect 3886 2771 3889 2968
rect 3886 2768 3894 2771
rect 3894 2732 3897 2748
rect 3870 2242 3873 2248
rect 3854 2142 3857 2168
rect 3854 2042 3857 2138
rect 3862 2102 3865 2228
rect 3854 1952 3857 1958
rect 3862 1852 3865 1968
rect 3854 1692 3857 1698
rect 3774 1168 3785 1171
rect 3766 1012 3769 1048
rect 3774 802 3777 1168
rect 3782 1032 3785 1048
rect 3790 942 3793 1238
rect 3798 1152 3801 1158
rect 3806 1152 3809 1158
rect 3814 1022 3817 1268
rect 3830 1262 3833 1278
rect 3838 1252 3841 1548
rect 3822 1248 3830 1251
rect 3806 912 3809 928
rect 3782 802 3785 848
rect 3822 762 3825 1248
rect 3830 1152 3833 1158
rect 3830 842 3833 938
rect 3830 752 3833 788
rect 3722 748 3726 751
rect 3718 452 3721 738
rect 3726 612 3729 738
rect 3774 722 3777 748
rect 3838 742 3841 1238
rect 3846 1162 3849 1548
rect 3854 1482 3857 1678
rect 3862 1522 3865 1528
rect 3854 1172 3857 1478
rect 3870 1452 3873 2218
rect 3878 1952 3881 2728
rect 3886 2212 3889 2668
rect 3894 2241 3897 2708
rect 3902 2372 3905 2738
rect 3910 2562 3913 2848
rect 3926 2772 3929 3148
rect 3942 3102 3945 3638
rect 3950 3582 3953 4028
rect 3958 3902 3961 4058
rect 3926 2721 3929 2738
rect 3922 2718 3929 2721
rect 3910 2442 3913 2488
rect 3894 2238 3902 2241
rect 3894 2052 3897 2238
rect 3906 2078 3910 2081
rect 3878 1572 3881 1948
rect 3878 1332 3881 1458
rect 3870 1172 3873 1298
rect 3878 1242 3881 1248
rect 3886 1242 3889 2048
rect 3894 1872 3897 1938
rect 3902 1882 3905 1918
rect 3910 1632 3913 2038
rect 3898 1538 3902 1541
rect 3894 1342 3897 1528
rect 3902 1282 3905 1458
rect 3910 1172 3913 1498
rect 3918 1492 3921 2678
rect 3926 2642 3929 2668
rect 3934 2512 3937 2798
rect 3942 2752 3945 3068
rect 3926 1962 3929 2188
rect 3934 1822 3937 2488
rect 3942 2232 3945 2658
rect 3950 2532 3953 3448
rect 3958 3062 3961 3588
rect 3966 3372 3969 4358
rect 3974 4142 3977 4498
rect 3974 3692 3977 3998
rect 3974 3382 3977 3528
rect 3982 3452 3985 4408
rect 3994 4308 3998 4311
rect 4006 4232 4009 4548
rect 4022 4332 4025 4458
rect 3990 4142 3993 4178
rect 3990 4122 3993 4128
rect 3990 4072 3993 4088
rect 3990 3752 3993 4068
rect 3998 3982 4001 4138
rect 4006 4072 4009 4088
rect 3994 3658 3998 3661
rect 3966 3348 3974 3351
rect 3966 3342 3969 3348
rect 3966 3302 3969 3338
rect 3966 3272 3969 3278
rect 3966 3012 3969 3248
rect 3966 2912 3969 2948
rect 3974 2732 3977 3338
rect 3982 3278 3990 3281
rect 3982 3272 3985 3278
rect 3990 3172 3993 3258
rect 3998 3062 4001 3598
rect 4006 3042 4009 3988
rect 4014 3672 4017 4318
rect 4022 4252 4025 4258
rect 4022 3602 4025 4028
rect 4014 3152 4017 3458
rect 4014 3082 4017 3108
rect 3994 2988 3998 2991
rect 4006 2981 4009 2998
rect 3998 2978 4009 2981
rect 3950 2472 3953 2478
rect 3950 2452 3953 2458
rect 3950 2392 3953 2428
rect 3942 2092 3945 2138
rect 3942 2062 3945 2078
rect 3866 1058 3870 1061
rect 3846 811 3849 828
rect 3846 808 3854 811
rect 3682 368 3686 371
rect 3750 252 3753 288
rect 3608 203 3610 207
rect 3614 203 3617 207
rect 3622 203 3624 207
rect 3654 72 3657 208
rect 3790 142 3793 608
rect 3814 571 3817 708
rect 3810 568 3817 571
rect 3798 352 3801 418
rect 3838 332 3841 588
rect 3846 402 3849 588
rect 3846 371 3849 398
rect 3846 368 3854 371
rect 3862 182 3865 628
rect 3870 492 3873 848
rect 3878 352 3881 448
rect 3870 342 3873 348
rect 3886 242 3889 1128
rect 3902 362 3905 1148
rect 3918 962 3921 1438
rect 3918 942 3921 948
rect 3926 892 3929 1488
rect 3934 1442 3937 1758
rect 3942 1622 3945 2048
rect 3934 1072 3937 1418
rect 3950 1412 3953 2338
rect 3958 2132 3961 2568
rect 3970 2498 3974 2501
rect 3982 2472 3985 2958
rect 3974 2432 3977 2438
rect 3982 2432 3985 2458
rect 3990 2422 3993 2428
rect 3978 2248 3982 2251
rect 3982 2042 3985 2178
rect 3990 2152 3993 2178
rect 3998 2132 4001 2978
rect 4006 2462 4009 2728
rect 4014 2692 4017 3058
rect 4022 3022 4025 3158
rect 4014 2662 4017 2668
rect 4006 2032 4009 2208
rect 4014 1982 4017 2648
rect 4022 2152 4025 2998
rect 4030 2942 4033 4338
rect 4046 4302 4049 4638
rect 4038 4272 4041 4278
rect 4046 4262 4049 4268
rect 4038 4252 4041 4258
rect 4038 3952 4041 4068
rect 4054 4062 4057 4658
rect 4102 4582 4105 4738
rect 4112 4703 4114 4707
rect 4118 4703 4121 4707
rect 4126 4703 4128 4707
rect 4134 4632 4137 4778
rect 4142 4712 4145 4838
rect 4254 4772 4257 4858
rect 4170 4658 4177 4661
rect 4062 4272 4065 4538
rect 4082 4458 4086 4461
rect 4082 4348 4086 4351
rect 4046 4042 4049 4048
rect 4062 3872 4065 4268
rect 4070 3922 4073 4128
rect 4046 3732 4049 3738
rect 4038 3302 4041 3358
rect 4038 3282 4041 3288
rect 4038 3082 4041 3128
rect 4046 3121 4049 3588
rect 4054 3432 4057 3868
rect 4062 3142 4065 3578
rect 4046 3118 4057 3121
rect 4030 2342 4033 2928
rect 4038 2922 4041 2938
rect 4054 2912 4057 3118
rect 4070 3112 4073 3918
rect 4078 3342 4081 4148
rect 4094 4142 4097 4528
rect 4102 4312 4105 4558
rect 4112 4503 4114 4507
rect 4118 4503 4121 4507
rect 4126 4503 4128 4507
rect 4134 4312 4137 4438
rect 4142 4321 4145 4488
rect 4150 4392 4153 4428
rect 4142 4318 4150 4321
rect 4112 4303 4114 4307
rect 4118 4303 4121 4307
rect 4126 4303 4128 4307
rect 4038 2222 4041 2468
rect 4022 2022 4025 2148
rect 4030 2042 4033 2198
rect 4038 2162 4041 2198
rect 4022 1972 4025 1998
rect 4026 1948 4030 1951
rect 3958 1562 3961 1798
rect 3966 1702 3969 1718
rect 3950 1202 3953 1278
rect 3934 1042 3937 1068
rect 3942 972 3945 1128
rect 3926 882 3929 888
rect 3926 612 3929 858
rect 3934 752 3937 838
rect 3950 662 3953 868
rect 3958 752 3961 1518
rect 3966 1471 3969 1548
rect 3974 1482 3977 1858
rect 3982 1772 3985 1928
rect 4006 1762 4009 1878
rect 3990 1702 3993 1758
rect 3998 1702 4001 1708
rect 4002 1688 4006 1691
rect 3990 1682 3993 1688
rect 3966 1468 3977 1471
rect 3966 1212 3969 1398
rect 3974 862 3977 1468
rect 3990 1462 3993 1548
rect 3982 872 3985 1308
rect 3990 992 3993 1458
rect 3998 1212 4001 1288
rect 3990 952 3993 958
rect 3950 622 3953 658
rect 3950 592 3953 618
rect 3982 382 3985 868
rect 3998 592 4001 1178
rect 4006 952 4009 1588
rect 4014 1412 4017 1928
rect 4038 1922 4041 2128
rect 4014 962 4017 1348
rect 4022 1312 4025 1608
rect 4030 1592 4033 1908
rect 4038 1842 4041 1918
rect 4038 1592 4041 1598
rect 4046 1432 4049 2698
rect 4054 2632 4057 2718
rect 4062 2702 4065 2748
rect 4070 2552 4073 3038
rect 4078 2972 4081 3338
rect 4078 2732 4081 2928
rect 4086 2812 4089 4108
rect 4094 4082 4097 4138
rect 4112 4103 4114 4107
rect 4118 4103 4121 4107
rect 4126 4103 4128 4107
rect 4094 4042 4097 4048
rect 4094 3342 4097 3708
rect 4102 3642 4105 3968
rect 4112 3903 4114 3907
rect 4118 3903 4121 3907
rect 4126 3903 4128 3907
rect 4134 3862 4137 4298
rect 4158 4282 4161 4508
rect 4174 4162 4177 4658
rect 4206 4372 4209 4648
rect 4214 4212 4217 4678
rect 4214 4192 4217 4208
rect 4174 4042 4177 4048
rect 4146 3958 4150 3961
rect 4174 3952 4177 4038
rect 4222 3982 4225 4378
rect 4230 4252 4233 4318
rect 4246 4292 4249 4588
rect 4230 4062 4233 4068
rect 4198 3918 4206 3921
rect 4182 3892 4185 3918
rect 4112 3703 4114 3707
rect 4118 3703 4121 3707
rect 4126 3703 4128 3707
rect 4102 3132 4105 3628
rect 4118 3532 4121 3538
rect 4112 3503 4114 3507
rect 4118 3503 4121 3507
rect 4126 3503 4128 3507
rect 4112 3303 4114 3307
rect 4118 3303 4121 3307
rect 4126 3303 4128 3307
rect 4134 3262 4137 3548
rect 4166 3442 4169 3878
rect 4182 3632 4185 3888
rect 4198 3862 4201 3918
rect 4190 3692 4193 3708
rect 4174 3412 4177 3428
rect 4054 2122 4057 2528
rect 4070 2332 4073 2398
rect 4058 2068 4062 2071
rect 4054 1562 4057 2068
rect 4062 1872 4065 1928
rect 4070 1792 4073 2328
rect 4078 2152 4081 2588
rect 4086 2492 4089 2748
rect 4094 2462 4097 3018
rect 4102 2712 4105 3108
rect 4112 3103 4114 3107
rect 4118 3103 4121 3107
rect 4126 3103 4128 3107
rect 4134 3052 4137 3258
rect 4142 3222 4145 3348
rect 4150 3322 4153 3328
rect 4142 3052 4145 3058
rect 4126 2932 4129 2938
rect 4112 2903 4114 2907
rect 4118 2903 4121 2907
rect 4126 2903 4128 2907
rect 4134 2772 4137 2938
rect 4112 2703 4114 2707
rect 4118 2703 4121 2707
rect 4126 2703 4128 2707
rect 4126 2522 4129 2548
rect 4102 2502 4105 2508
rect 4112 2503 4114 2507
rect 4118 2503 4121 2507
rect 4126 2503 4128 2507
rect 4112 2303 4114 2307
rect 4118 2303 4121 2307
rect 4126 2303 4128 2307
rect 4086 2022 4089 2218
rect 4094 2011 4097 2118
rect 4090 2008 4097 2011
rect 4078 1792 4081 1958
rect 4086 1952 4089 1958
rect 4094 1902 4097 1978
rect 4062 1572 4065 1768
rect 4078 1762 4081 1768
rect 4078 1692 4081 1718
rect 4078 1632 4081 1638
rect 4070 1562 4073 1628
rect 4078 1552 4081 1578
rect 4046 1352 4049 1368
rect 4054 1332 4057 1358
rect 4014 752 4017 958
rect 3998 542 4001 588
rect 3962 348 3966 351
rect 3666 78 3670 81
rect 3822 62 3825 128
rect 3946 68 3950 71
rect 3410 58 3414 61
rect 3510 52 3513 58
rect 3998 52 4001 248
rect 4006 172 4009 748
rect 4014 462 4017 688
rect 4022 622 4025 818
rect 4030 692 4033 1078
rect 4022 112 4025 618
rect 4030 552 4033 558
rect 4030 362 4033 458
rect 4038 142 4041 928
rect 4046 672 4049 1258
rect 4054 1162 4057 1168
rect 4054 1052 4057 1118
rect 4062 852 4065 1508
rect 4070 1182 4073 1318
rect 4078 1112 4081 1348
rect 4086 1222 4089 1898
rect 4094 1832 4097 1898
rect 4094 1072 4097 1828
rect 4102 1592 4105 2258
rect 4118 2252 4121 2268
rect 4112 2103 4114 2107
rect 4118 2103 4121 2107
rect 4126 2103 4128 2107
rect 4134 2082 4137 2348
rect 4110 2002 4113 2038
rect 4118 2032 4121 2038
rect 4134 2022 4137 2058
rect 4112 1903 4114 1907
rect 4118 1903 4121 1907
rect 4126 1903 4128 1907
rect 4118 1722 4121 1868
rect 4112 1703 4114 1707
rect 4118 1703 4121 1707
rect 4126 1703 4128 1707
rect 4102 1512 4105 1578
rect 4112 1503 4114 1507
rect 4118 1503 4121 1507
rect 4126 1503 4128 1507
rect 4126 1482 4129 1488
rect 4134 1392 4137 1998
rect 4142 1422 4145 2858
rect 4150 2652 4153 3268
rect 4158 3122 4161 3318
rect 4150 2152 4153 2558
rect 4158 2552 4161 3038
rect 4166 3022 4169 3358
rect 4174 3132 4177 3408
rect 4190 3332 4193 3688
rect 4198 3462 4201 3798
rect 4206 3472 4209 3638
rect 4214 3592 4217 3978
rect 4226 3958 4230 3961
rect 4222 3852 4225 3948
rect 4230 3872 4233 3928
rect 4206 3302 4209 3468
rect 4166 2892 4169 3018
rect 4182 2962 4185 3288
rect 4190 3192 4193 3278
rect 4182 2932 4185 2938
rect 4170 2858 4174 2861
rect 4182 2852 4185 2888
rect 4190 2862 4193 2878
rect 4174 2758 4182 2761
rect 4158 2542 4161 2548
rect 4158 2292 4161 2508
rect 4174 2472 4177 2758
rect 4182 2642 4185 2728
rect 4190 2512 4193 2848
rect 4198 2812 4201 3068
rect 4206 3022 4209 3148
rect 4206 2992 4209 3018
rect 4206 2682 4209 2938
rect 4214 2532 4217 3528
rect 4222 3272 4225 3408
rect 4222 2822 4225 3238
rect 4230 2882 4233 3868
rect 4238 3352 4241 4268
rect 4246 4142 4249 4278
rect 4246 3882 4249 4058
rect 4254 3932 4257 4768
rect 4262 4262 4265 4268
rect 4270 4092 4273 4408
rect 4278 4342 4281 4538
rect 4294 4342 4297 4738
rect 4350 4672 4353 4748
rect 4366 4692 4369 4808
rect 4310 4352 4313 4528
rect 4350 4522 4353 4668
rect 4446 4662 4449 4798
rect 4326 4442 4329 4458
rect 4398 4422 4401 4538
rect 4262 4062 4265 4088
rect 4270 3922 4273 4068
rect 4258 3878 4262 3881
rect 4262 3832 4265 3838
rect 4238 3222 4241 3258
rect 4246 3192 4249 3338
rect 4182 2372 4185 2408
rect 4178 2348 4182 2351
rect 4150 2032 4153 2148
rect 4166 2138 4174 2141
rect 4166 2102 4169 2138
rect 4150 1692 4153 1958
rect 4166 1942 4169 2018
rect 4174 1872 4177 2048
rect 4182 1972 4185 2258
rect 4190 2032 4193 2448
rect 4198 2072 4201 2348
rect 4206 2292 4209 2458
rect 4222 2422 4225 2588
rect 4230 2232 4233 2738
rect 4238 2382 4241 3088
rect 4246 2322 4249 2338
rect 4206 2192 4209 2208
rect 4222 2152 4225 2228
rect 4162 1848 4166 1851
rect 4174 1848 4182 1851
rect 4174 1822 4177 1848
rect 4158 1532 4161 1648
rect 4138 1368 4145 1371
rect 4112 1303 4114 1307
rect 4118 1303 4121 1307
rect 4126 1303 4128 1307
rect 4102 912 4105 1148
rect 4114 1128 4118 1131
rect 4112 1103 4114 1107
rect 4118 1103 4121 1107
rect 4126 1103 4128 1107
rect 4142 1002 4145 1368
rect 4150 932 4153 1518
rect 4166 1512 4169 1528
rect 4158 1172 4161 1498
rect 4112 903 4114 907
rect 4118 903 4121 907
rect 4126 903 4128 907
rect 4062 682 4065 688
rect 4050 658 4054 661
rect 4054 542 4057 548
rect 4070 362 4073 648
rect 4086 472 4089 748
rect 4112 703 4114 707
rect 4118 703 4121 707
rect 4126 703 4128 707
rect 4094 562 4097 598
rect 4102 202 4105 548
rect 4130 518 4134 521
rect 4112 503 4114 507
rect 4118 503 4121 507
rect 4126 503 4128 507
rect 4138 348 4142 351
rect 4112 303 4114 307
rect 4118 303 4121 307
rect 4126 303 4128 307
rect 4174 272 4177 1158
rect 4182 972 4185 1498
rect 4190 1352 4193 1938
rect 4202 1848 4206 1851
rect 4214 1692 4217 2128
rect 4230 1972 4233 2228
rect 4238 2032 4241 2308
rect 4254 2232 4257 3638
rect 4262 3312 4265 3698
rect 4270 3662 4273 3868
rect 4278 3702 4281 4338
rect 4286 4052 4289 4138
rect 4286 3862 4289 3998
rect 4294 3992 4297 4338
rect 4310 4072 4313 4258
rect 4298 3968 4302 3971
rect 4262 3162 4265 3298
rect 4262 3112 4265 3158
rect 4262 3062 4265 3068
rect 4262 2472 4265 2918
rect 4270 2482 4273 3148
rect 4278 3032 4281 3698
rect 4310 3592 4313 4068
rect 4318 3872 4321 4068
rect 4318 3752 4321 3848
rect 4318 3742 4321 3748
rect 4294 3352 4297 3588
rect 4310 3542 4313 3568
rect 4286 3012 4289 3048
rect 4278 2612 4281 2758
rect 4286 2662 4289 2688
rect 4238 1882 4241 1978
rect 4222 1762 4225 1798
rect 4222 1712 4225 1738
rect 4226 1688 4230 1691
rect 4182 552 4185 968
rect 4190 722 4193 1048
rect 4198 1012 4201 1648
rect 4198 912 4201 938
rect 4198 472 4201 908
rect 4206 882 4209 1588
rect 4246 1472 4249 2168
rect 4262 1952 4265 2328
rect 4258 1758 4262 1761
rect 4254 1452 4257 1468
rect 4230 1142 4233 1368
rect 4206 472 4209 538
rect 4182 182 4185 468
rect 4202 348 4206 351
rect 4112 103 4114 107
rect 4118 103 4121 107
rect 4126 103 4128 107
rect 4198 102 4201 338
rect 4238 222 4241 1258
rect 4246 892 4249 1408
rect 4254 1192 4257 1248
rect 4250 838 4254 841
rect 4270 822 4273 2478
rect 4278 1892 4281 2558
rect 4302 2332 4305 3508
rect 4310 2952 4313 3218
rect 4318 3122 4321 3618
rect 4286 2252 4289 2258
rect 4294 2072 4297 2198
rect 4278 1692 4281 1888
rect 4278 1341 4281 1548
rect 4286 1352 4289 1868
rect 4294 1792 4297 1888
rect 4294 1672 4297 1758
rect 4302 1752 4305 1998
rect 4278 1338 4286 1341
rect 4302 1322 4305 1708
rect 4310 1302 4313 2318
rect 4318 2172 4321 3118
rect 4326 2692 4329 3948
rect 4334 3462 4337 4348
rect 4342 3472 4345 4068
rect 4350 3782 4353 4318
rect 4358 4062 4361 4388
rect 4358 3842 4361 3918
rect 4374 3902 4377 4168
rect 4394 3958 4398 3961
rect 4358 3652 4361 3658
rect 4334 2942 4337 3388
rect 4342 3062 4345 3068
rect 4334 2912 4337 2938
rect 4342 2932 4345 3038
rect 4334 2812 4337 2828
rect 4326 2322 4329 2638
rect 4318 1492 4321 1968
rect 4326 1882 4329 1988
rect 4334 1942 4337 2538
rect 4342 2522 4345 2928
rect 4350 2852 4353 3068
rect 4350 2812 4353 2818
rect 4342 2452 4345 2488
rect 4350 2372 4353 2768
rect 4358 2542 4361 3478
rect 4366 3472 4369 3698
rect 4366 2682 4369 3438
rect 4374 2832 4377 3868
rect 4382 3262 4385 3458
rect 4390 3352 4393 3948
rect 4398 3862 4401 3938
rect 4398 3472 4401 3828
rect 4406 3632 4409 4518
rect 4422 4372 4425 4628
rect 4478 4548 4486 4551
rect 4430 4532 4433 4548
rect 4478 4542 4481 4548
rect 4494 4522 4497 4548
rect 4510 4542 4513 4718
rect 4550 4632 4553 4698
rect 4554 4578 4558 4581
rect 4522 4538 4526 4541
rect 4430 4372 4433 4458
rect 4430 4262 4433 4368
rect 4414 3702 4417 3838
rect 4422 3812 4425 4058
rect 4430 4042 4433 4228
rect 4438 3951 4441 4468
rect 4446 4352 4449 4368
rect 4454 4192 4457 4488
rect 4502 4312 4505 4438
rect 4538 4408 4542 4411
rect 4446 4032 4449 4118
rect 4438 3948 4446 3951
rect 4458 3948 4465 3951
rect 4442 3858 4446 3861
rect 4454 3662 4457 3888
rect 4462 3822 4465 3948
rect 4454 3648 4462 3651
rect 4454 3612 4457 3648
rect 4390 3232 4393 3348
rect 4366 2592 4369 2678
rect 4358 2472 4361 2478
rect 4350 2292 4353 2348
rect 4358 2312 4361 2318
rect 4346 2148 4350 2151
rect 4342 2102 4345 2138
rect 4342 1892 4345 2098
rect 4334 1652 4337 1678
rect 4322 1468 4329 1471
rect 4326 972 4329 1468
rect 4334 1322 4337 1648
rect 4342 1602 4345 1888
rect 4350 1652 4353 1888
rect 4346 1588 4353 1591
rect 4350 1582 4353 1588
rect 4358 1482 4361 2258
rect 4366 2172 4369 2528
rect 4382 2452 4385 3008
rect 4398 2942 4401 3458
rect 4406 3262 4409 3548
rect 4430 3532 4433 3568
rect 4470 3522 4473 3858
rect 4478 3622 4481 4138
rect 4490 3808 4494 3811
rect 4502 3672 4505 3978
rect 4510 3752 4513 4378
rect 4558 4342 4561 4528
rect 4582 4442 4585 4638
rect 4590 4352 4593 4648
rect 4598 4642 4601 4658
rect 4606 4462 4609 4618
rect 4558 4332 4561 4338
rect 4606 4262 4609 4268
rect 4530 4148 4534 4151
rect 4542 4142 4545 4158
rect 4550 4132 4553 4138
rect 4502 3542 4505 3668
rect 4510 3562 4513 3718
rect 4458 3468 4465 3471
rect 4426 3298 4430 3301
rect 4438 3222 4441 3288
rect 4398 2742 4401 2928
rect 4390 2562 4393 2568
rect 4374 2132 4377 2348
rect 4382 2322 4385 2438
rect 4382 2132 4385 2318
rect 4390 2302 4393 2308
rect 4366 1662 4369 2118
rect 4374 1832 4377 1948
rect 4382 1931 4385 2118
rect 4390 2052 4393 2228
rect 4398 2202 4401 2718
rect 4382 1928 4390 1931
rect 4382 1872 4385 1918
rect 4374 1782 4377 1818
rect 4378 1748 4382 1751
rect 4374 1602 4377 1658
rect 4362 1468 4366 1471
rect 4374 1262 4377 1598
rect 4390 1572 4393 1908
rect 4398 1552 4401 2198
rect 4406 2062 4409 2858
rect 4414 2472 4417 2728
rect 4414 2252 4417 2338
rect 4414 2062 4417 2228
rect 4406 1882 4409 2008
rect 4406 1672 4409 1708
rect 4390 1342 4393 1358
rect 4346 1258 4350 1261
rect 4342 1162 4345 1168
rect 4326 832 4329 968
rect 4270 731 4273 738
rect 4270 728 4278 731
rect 4286 262 4289 708
rect 4294 542 4297 808
rect 4302 792 4305 808
rect 4310 752 4313 758
rect 4326 472 4329 758
rect 4350 732 4353 1238
rect 4358 1162 4361 1178
rect 4358 932 4361 1018
rect 4366 862 4369 1258
rect 4374 1138 4382 1141
rect 4358 858 4366 861
rect 4358 502 4361 858
rect 4314 468 4318 471
rect 4358 362 4361 498
rect 4366 442 4369 748
rect 4374 722 4377 1138
rect 4390 962 4393 1148
rect 4414 972 4417 1958
rect 4422 1682 4425 2828
rect 4430 2502 4433 2828
rect 4438 2742 4441 3218
rect 4462 3012 4465 3468
rect 4470 3242 4473 3518
rect 4510 3362 4513 3548
rect 4518 3512 4521 4008
rect 4526 3332 4529 3858
rect 4550 3852 4553 3948
rect 4558 3902 4561 4248
rect 4598 4172 4601 4198
rect 4522 3328 4526 3331
rect 4534 3272 4537 3528
rect 4542 3282 4545 3838
rect 4502 3148 4510 3151
rect 4462 2982 4465 2988
rect 4454 2942 4457 2978
rect 4470 2972 4473 3098
rect 4490 3058 4497 3061
rect 4462 2922 4465 2958
rect 4454 2852 4457 2878
rect 4462 2772 4465 2898
rect 4450 2718 4454 2721
rect 4430 2492 4433 2498
rect 4430 1962 4433 2468
rect 4438 2462 4441 2468
rect 4446 2292 4449 2608
rect 4454 1962 4457 2488
rect 4462 2262 4465 2728
rect 4470 2352 4473 2538
rect 4478 2402 4481 3018
rect 4486 2442 4489 3038
rect 4494 2992 4497 3058
rect 4494 2532 4497 2568
rect 4470 2342 4473 2348
rect 4466 2258 4473 2261
rect 4470 2222 4473 2258
rect 4486 2172 4489 2178
rect 4494 2102 4497 2528
rect 4474 2078 4478 2081
rect 4438 1832 4441 1888
rect 4454 1862 4457 1958
rect 4462 1902 4465 2048
rect 4434 1748 4438 1751
rect 4422 1312 4425 1678
rect 4446 1662 4449 1698
rect 4422 1132 4425 1138
rect 4430 1032 4433 1478
rect 4438 1242 4441 1658
rect 4390 762 4393 958
rect 4430 772 4433 1028
rect 4446 662 4449 1418
rect 4454 882 4457 1838
rect 4462 1212 4465 1888
rect 4478 1872 4481 2008
rect 4486 1851 4489 2028
rect 4494 1972 4497 2098
rect 4482 1848 4489 1851
rect 4470 1752 4473 1788
rect 4470 1662 4473 1668
rect 4470 912 4473 1598
rect 4478 892 4481 1158
rect 4486 1142 4489 1218
rect 4486 892 4489 938
rect 4410 548 4414 551
rect 4386 468 4390 471
rect 4370 258 4374 261
rect 4382 142 4385 398
rect 4210 138 4214 141
rect 4226 138 4230 141
rect 4406 81 4409 418
rect 4414 202 4417 448
rect 4422 392 4425 538
rect 4446 262 4449 538
rect 4454 272 4457 608
rect 4470 492 4473 838
rect 4478 532 4481 538
rect 4486 492 4489 828
rect 4494 552 4497 1958
rect 4502 1652 4505 3148
rect 4518 2862 4521 3118
rect 4526 2872 4529 3048
rect 4526 2842 4529 2848
rect 4526 2542 4529 2548
rect 4534 2502 4537 3148
rect 4550 2891 4553 3528
rect 4558 3442 4561 3868
rect 4566 3452 4569 4118
rect 4574 3862 4577 3878
rect 4574 3742 4577 3748
rect 4558 3262 4561 3348
rect 4550 2888 4561 2891
rect 4546 2858 4550 2861
rect 4510 1862 4513 2068
rect 4502 1162 4505 1488
rect 4518 1342 4521 2458
rect 4526 2132 4529 2498
rect 4550 2452 4553 2488
rect 4538 2358 4542 2361
rect 4518 1201 4521 1338
rect 4510 1198 4521 1201
rect 4526 1202 4529 2068
rect 4534 2002 4537 2288
rect 4550 2172 4553 2448
rect 4558 2262 4561 2888
rect 4566 2782 4569 3368
rect 4574 3352 4577 3498
rect 4574 3332 4577 3338
rect 4574 2921 4577 3248
rect 4582 3042 4585 3928
rect 4590 3372 4593 4078
rect 4606 3872 4609 4258
rect 4590 3352 4593 3358
rect 4590 3282 4593 3308
rect 4590 2962 4593 2968
rect 4598 2962 4601 3748
rect 4606 3472 4609 3738
rect 4574 2918 4582 2921
rect 4574 2732 4577 2918
rect 4566 2502 4569 2668
rect 4598 2562 4601 2868
rect 4566 2232 4569 2478
rect 4574 2432 4577 2538
rect 4542 1852 4545 1998
rect 4542 1672 4545 1818
rect 4550 1812 4553 2128
rect 4550 1672 4553 1808
rect 4550 1642 4553 1668
rect 4510 942 4513 1198
rect 4502 782 4505 908
rect 4518 802 4521 1188
rect 4526 1168 4534 1171
rect 4526 1162 4529 1168
rect 4542 1152 4545 1158
rect 4526 1062 4529 1118
rect 4550 1072 4553 1348
rect 4518 762 4521 798
rect 4514 748 4518 751
rect 4482 348 4486 351
rect 4470 272 4473 338
rect 4446 172 4449 258
rect 4402 78 4409 81
rect 4206 71 4209 78
rect 4438 72 4441 148
rect 4470 132 4473 268
rect 4494 192 4497 518
rect 4518 362 4521 548
rect 4526 452 4529 1058
rect 4558 862 4561 1848
rect 4566 1422 4569 2128
rect 4574 2052 4577 2428
rect 4598 2282 4601 2548
rect 4598 2222 4601 2278
rect 4574 1922 4577 1998
rect 4582 1802 4585 2158
rect 4574 1792 4577 1798
rect 4590 1762 4593 1938
rect 4578 1728 4582 1731
rect 4582 1661 4585 1678
rect 4578 1658 4585 1661
rect 4578 1268 4582 1271
rect 4534 452 4537 718
rect 4558 352 4561 728
rect 4566 372 4569 1158
rect 4574 992 4577 1258
rect 4530 348 4534 351
rect 4518 142 4521 148
rect 4566 131 4569 138
rect 4566 128 4574 131
rect 4206 68 4214 71
rect 4086 52 4089 68
rect 4542 62 4545 68
rect 4582 62 4585 1198
rect 4590 702 4593 1748
rect 4606 1602 4609 3468
rect 4614 3362 4617 4858
rect 4632 4803 4634 4807
rect 4638 4803 4641 4807
rect 4646 4803 4648 4807
rect 4622 4612 4625 4668
rect 4632 4603 4634 4607
rect 4638 4603 4641 4607
rect 4646 4603 4648 4607
rect 4710 4512 4713 4748
rect 4750 4542 4753 4548
rect 4632 4403 4634 4407
rect 4638 4403 4641 4407
rect 4646 4403 4648 4407
rect 4622 4192 4625 4218
rect 4632 4203 4634 4207
rect 4638 4203 4641 4207
rect 4646 4203 4648 4207
rect 4650 4158 4654 4161
rect 4626 4148 4630 4151
rect 4654 4092 4657 4098
rect 4632 4003 4634 4007
rect 4638 4003 4641 4007
rect 4646 4003 4648 4007
rect 4654 3952 4657 3998
rect 4662 3992 4665 4468
rect 4694 4358 4702 4361
rect 4694 4342 4697 4358
rect 4710 4302 4713 4508
rect 4674 4258 4681 4261
rect 4678 4222 4681 4258
rect 4694 4162 4697 4168
rect 4710 4142 4713 4298
rect 4734 4082 4737 4138
rect 4738 4078 4742 4081
rect 4678 4052 4681 4058
rect 4678 3932 4681 4048
rect 4694 3932 4697 3938
rect 4632 3803 4634 3807
rect 4638 3803 4641 3807
rect 4646 3803 4648 3807
rect 4622 3482 4625 3648
rect 4662 3632 4665 3718
rect 4632 3603 4634 3607
rect 4638 3603 4641 3607
rect 4646 3603 4648 3607
rect 4632 3403 4634 3407
rect 4638 3403 4641 3407
rect 4646 3403 4648 3407
rect 4654 3372 4657 3628
rect 4614 3052 4617 3318
rect 4632 3203 4634 3207
rect 4638 3203 4641 3207
rect 4646 3203 4648 3207
rect 4614 1932 4617 2958
rect 4622 2882 4625 3008
rect 4632 3003 4634 3007
rect 4638 3003 4641 3007
rect 4646 3003 4648 3007
rect 4630 2942 4633 2948
rect 4622 2862 4625 2868
rect 4622 2572 4625 2838
rect 4632 2803 4634 2807
rect 4638 2803 4641 2807
rect 4646 2803 4648 2807
rect 4646 2672 4649 2788
rect 4654 2612 4657 3358
rect 4670 3302 4673 3718
rect 4678 3452 4681 3928
rect 4686 3602 4689 3738
rect 4702 3702 4705 3978
rect 4706 3658 4710 3661
rect 4710 3552 4713 3638
rect 4714 3468 4718 3471
rect 4662 3142 4665 3188
rect 4662 2792 4665 3138
rect 4670 3062 4673 3298
rect 4682 3138 4686 3141
rect 4686 2958 4694 2961
rect 4686 2902 4689 2958
rect 4702 2892 4705 3308
rect 4632 2603 4634 2607
rect 4638 2603 4641 2607
rect 4646 2603 4648 2607
rect 4654 2412 4657 2518
rect 4632 2403 4634 2407
rect 4638 2403 4641 2407
rect 4646 2403 4648 2407
rect 4642 2318 4649 2321
rect 4646 2312 4649 2318
rect 4642 2278 4646 2281
rect 4632 2203 4634 2207
rect 4638 2203 4641 2207
rect 4646 2203 4648 2207
rect 4654 2141 4657 2388
rect 4650 2138 4657 2141
rect 4632 2003 4634 2007
rect 4638 2003 4641 2007
rect 4646 2003 4648 2007
rect 4646 1952 4649 1968
rect 4614 1712 4617 1928
rect 4654 1882 4657 2138
rect 4662 2072 4665 2298
rect 4632 1803 4634 1807
rect 4638 1803 4641 1807
rect 4646 1803 4648 1807
rect 4630 1672 4633 1678
rect 4598 1232 4601 1278
rect 4598 552 4601 648
rect 4606 212 4609 1588
rect 4614 872 4617 1668
rect 4654 1612 4657 1628
rect 4632 1603 4634 1607
rect 4638 1603 4641 1607
rect 4646 1603 4648 1607
rect 4632 1403 4634 1407
rect 4638 1403 4641 1407
rect 4646 1403 4648 1407
rect 4632 1203 4634 1207
rect 4638 1203 4641 1207
rect 4646 1203 4648 1207
rect 4642 1148 4646 1151
rect 4632 1003 4634 1007
rect 4638 1003 4641 1007
rect 4646 1003 4648 1007
rect 4614 682 4617 868
rect 4622 622 4625 828
rect 4632 803 4634 807
rect 4638 803 4641 807
rect 4646 803 4648 807
rect 4654 792 4657 1488
rect 4662 1272 4665 2018
rect 4670 1922 4673 2668
rect 4678 2152 4681 2748
rect 4686 2652 4689 2678
rect 4670 1672 4673 1908
rect 4686 1692 4689 2558
rect 4694 2312 4697 2618
rect 4702 2452 4705 2718
rect 4702 2322 4705 2338
rect 4694 2258 4702 2261
rect 4670 1662 4673 1668
rect 4678 1302 4681 1648
rect 4678 1262 4681 1268
rect 4630 672 4633 768
rect 4662 742 4665 1138
rect 4678 1092 4681 1258
rect 4670 952 4673 958
rect 4678 942 4681 1008
rect 4632 603 4634 607
rect 4638 603 4641 607
rect 4646 603 4648 607
rect 4654 542 4657 618
rect 4622 232 4625 538
rect 4632 403 4634 407
rect 4638 403 4641 407
rect 4646 403 4648 407
rect 4686 382 4689 1638
rect 4694 1412 4697 2258
rect 4702 2242 4705 2248
rect 4702 1952 4705 1958
rect 4710 1912 4713 2848
rect 4718 1872 4721 3448
rect 4726 3382 4729 3458
rect 4734 3161 4737 3788
rect 4742 3492 4745 3728
rect 4750 3572 4753 4538
rect 4758 4452 4761 4458
rect 4766 3942 4769 4648
rect 4762 3938 4766 3941
rect 4758 3742 4761 3748
rect 4742 3302 4745 3488
rect 4758 3361 4761 3538
rect 4758 3358 4766 3361
rect 4730 3158 4737 3161
rect 4726 2192 4729 3148
rect 4734 2462 4737 2858
rect 4742 2742 4745 3208
rect 4750 3032 4753 3328
rect 4758 3132 4761 3138
rect 4750 2862 4753 2868
rect 4758 2772 4761 3128
rect 4758 2662 4761 2748
rect 4742 2492 4745 2578
rect 4766 2562 4769 3278
rect 4774 3102 4777 4788
rect 4782 3702 4785 4838
rect 4798 3652 4801 3678
rect 4786 3358 4790 3361
rect 4782 3222 4785 3258
rect 4774 2692 4777 3078
rect 4782 2972 4785 3218
rect 4790 2852 4793 3338
rect 4806 3242 4809 4868
rect 4866 4858 4870 4861
rect 4814 4452 4817 4458
rect 4814 4242 4817 4448
rect 4814 3892 4817 3958
rect 4822 3722 4825 4858
rect 4858 4648 4862 4651
rect 4870 4532 4873 4698
rect 4834 4408 4841 4411
rect 4838 4322 4841 4408
rect 4870 4312 4873 4358
rect 4870 4042 4873 4308
rect 4758 2548 4766 2551
rect 4746 2468 4750 2471
rect 4750 2252 4753 2268
rect 4742 2162 4745 2178
rect 4726 1882 4729 2148
rect 4742 1952 4745 2068
rect 4702 1292 4705 1818
rect 4710 1592 4713 1868
rect 4734 1682 4737 1938
rect 4750 1851 4753 1958
rect 4746 1848 4753 1851
rect 4718 1632 4721 1668
rect 4710 1232 4713 1438
rect 4726 1432 4729 1638
rect 4742 1521 4745 1788
rect 4734 1518 4745 1521
rect 4694 1152 4697 1158
rect 4694 1002 4697 1018
rect 4694 942 4697 948
rect 4702 881 4705 1178
rect 4710 1062 4713 1228
rect 4710 952 4713 958
rect 4698 878 4705 881
rect 4694 302 4697 848
rect 4710 252 4713 938
rect 4718 912 4721 1248
rect 4726 882 4729 1428
rect 4734 482 4737 1518
rect 4742 1482 4745 1488
rect 4750 1432 4753 1848
rect 4742 542 4745 1018
rect 4750 702 4753 1238
rect 4758 1062 4761 2548
rect 4790 2532 4793 2548
rect 4778 2528 4785 2531
rect 4766 2122 4769 2348
rect 4766 1842 4769 2108
rect 4766 1482 4769 1838
rect 4774 1282 4777 2188
rect 4782 2062 4785 2528
rect 4790 2152 4793 2158
rect 4782 1672 4785 1698
rect 4782 1302 4785 1408
rect 4758 1052 4761 1058
rect 4766 862 4769 1278
rect 4774 952 4777 1258
rect 4782 942 4785 948
rect 4766 712 4769 858
rect 4790 832 4793 2128
rect 4798 2072 4801 2158
rect 4806 1951 4809 3158
rect 4814 2082 4817 2908
rect 4830 2752 4833 3278
rect 4822 2322 4825 2728
rect 4838 2482 4841 2948
rect 4846 2902 4849 3668
rect 4854 3292 4857 3658
rect 4862 3232 4865 3278
rect 4870 3002 4873 3348
rect 4878 2672 4881 4868
rect 4930 4858 4934 4861
rect 4886 4562 4889 4578
rect 4886 2952 4889 3538
rect 4894 3342 4897 4848
rect 4918 4472 4921 4758
rect 4918 4382 4921 4468
rect 4902 3942 4905 4268
rect 4918 3972 4921 4378
rect 4902 3582 4905 3938
rect 4918 3882 4921 3968
rect 4918 3352 4921 3848
rect 4934 3442 4937 4818
rect 4942 4152 4945 4528
rect 4894 3092 4897 3168
rect 4834 2278 4838 2281
rect 4806 1948 4814 1951
rect 4822 1892 4825 2148
rect 4806 1742 4809 1848
rect 4806 1592 4809 1738
rect 4750 662 4753 668
rect 4742 422 4745 538
rect 4632 203 4634 207
rect 4638 203 4641 207
rect 4646 203 4648 207
rect 4742 142 4745 418
rect 4750 192 4753 518
rect 4758 252 4761 338
rect 4766 272 4769 578
rect 4758 152 4761 248
rect 4758 132 4761 148
rect 4798 142 4801 1568
rect 4806 792 4809 1238
rect 4814 1062 4817 1858
rect 4806 462 4809 748
rect 4814 322 4817 1048
rect 4822 172 4825 1878
rect 4830 1562 4833 2198
rect 4838 942 4841 2208
rect 4846 1872 4849 2568
rect 4862 2472 4865 2598
rect 4866 2468 4873 2471
rect 4854 2172 4857 2468
rect 4854 2158 4862 2161
rect 4854 2142 4857 2158
rect 4846 1792 4849 1858
rect 4854 1702 4857 1878
rect 4862 1852 4865 1978
rect 4870 1892 4873 2468
rect 4886 2421 4889 2948
rect 4902 2892 4905 2898
rect 4898 2758 4902 2761
rect 4878 2418 4889 2421
rect 4878 1932 4881 2418
rect 4886 2282 4889 2388
rect 4870 1722 4873 1868
rect 4854 1532 4857 1688
rect 4862 1682 4865 1688
rect 4854 1472 4857 1528
rect 4870 1502 4873 1718
rect 4846 992 4849 1368
rect 4830 152 4833 658
rect 4602 108 4606 111
rect 4846 62 4849 988
rect 4854 862 4857 1408
rect 4862 1142 4865 1378
rect 4854 692 4857 858
rect 4862 542 4865 1138
rect 4854 282 4857 368
rect 4854 142 4857 278
rect 4866 258 4870 261
rect 4878 242 4881 1918
rect 4886 1332 4889 2258
rect 4886 712 4889 958
rect 4894 112 4897 2458
rect 4902 2352 4905 2728
rect 4902 2152 4905 2158
rect 4910 2132 4913 3138
rect 4902 2092 4905 2098
rect 4910 1762 4913 1848
rect 4918 1832 4921 3308
rect 4926 2352 4929 3238
rect 4934 3162 4937 3278
rect 4950 3182 4953 4828
rect 4982 4022 4985 4818
rect 4978 3358 4982 3361
rect 4966 3352 4969 3358
rect 4998 3351 5001 3378
rect 4998 3348 5006 3351
rect 4942 3132 4945 3138
rect 4942 2971 4945 3078
rect 4942 2968 4950 2971
rect 4918 1772 4921 1828
rect 4918 1732 4921 1738
rect 4902 1471 4905 1568
rect 4902 1468 4910 1471
rect 4926 1382 4929 2268
rect 4934 2152 4937 2618
rect 4942 2432 4945 2968
rect 4942 2362 4945 2428
rect 4942 2322 4945 2358
rect 4934 1482 4937 2098
rect 4942 1492 4945 2068
rect 4902 952 4905 968
rect 4918 372 4921 698
rect 4926 592 4929 1118
rect 4942 82 4945 888
rect 4950 732 4953 2118
rect 4958 102 4961 2738
rect 4966 1852 4969 3338
rect 4974 3092 4977 3298
rect 4974 2832 4977 3088
rect 4982 2972 4985 3188
rect 4974 2542 4977 2828
rect 4974 1772 4977 2478
rect 4982 1732 4985 2678
rect 4982 1362 4985 1728
rect 4966 142 4969 728
rect 4982 662 4985 1348
rect 4954 78 4958 81
rect 4990 62 4993 3148
rect 4998 2692 5001 2948
rect 5014 2822 5017 4808
rect 5022 2922 5025 4788
rect 5034 4478 5038 4481
rect 5022 2898 5030 2901
rect 5022 2782 5025 2898
rect 5014 2742 5017 2758
rect 4998 2082 5001 2518
rect 5006 2092 5009 2578
rect 5014 2112 5017 2658
rect 5022 2452 5025 2778
rect 5030 2402 5033 2888
rect 5046 2642 5049 4858
rect 5054 4662 5057 4668
rect 5054 4152 5057 4458
rect 5062 4371 5065 4868
rect 5106 4858 5110 4861
rect 5070 4382 5073 4858
rect 5062 4368 5073 4371
rect 5062 4102 5065 4268
rect 5054 3832 5057 3848
rect 5054 3562 5057 3828
rect 5058 3348 5062 3351
rect 5070 3042 5073 4368
rect 5078 3342 5081 3858
rect 5086 3682 5089 4218
rect 4998 82 5001 2058
rect 5006 942 5009 2068
rect 5014 1872 5017 1878
rect 5022 1722 5025 1998
rect 5014 1542 5017 1558
rect 5014 1242 5017 1248
rect 5006 582 5009 938
rect 5022 792 5025 1698
rect 5030 1262 5033 2318
rect 5038 2062 5041 2508
rect 5046 1572 5049 2368
rect 5038 732 5041 1528
rect 5046 1361 5049 1558
rect 5054 1502 5057 2348
rect 5062 2312 5065 2888
rect 5078 2792 5081 3328
rect 5086 3112 5089 3338
rect 5086 3082 5089 3108
rect 5062 2082 5065 2298
rect 5070 2132 5073 2668
rect 5070 2072 5073 2128
rect 5062 1932 5065 2068
rect 5062 1672 5065 1928
rect 5070 1652 5073 2048
rect 5078 1742 5081 2618
rect 5086 2032 5089 3038
rect 5094 2432 5097 4808
rect 5102 2932 5105 4838
rect 5110 2762 5113 3668
rect 5118 2962 5121 4668
rect 5158 3541 5161 4538
rect 5166 4002 5169 4558
rect 5154 3538 5161 3541
rect 5110 2642 5113 2648
rect 5094 2382 5097 2428
rect 5094 2362 5097 2368
rect 5102 2351 5105 2538
rect 5110 2472 5113 2628
rect 5118 2572 5121 2938
rect 5126 2572 5129 3358
rect 5134 3062 5137 3348
rect 5158 3332 5161 3538
rect 5166 3362 5169 3428
rect 5118 2542 5121 2568
rect 5126 2552 5129 2558
rect 5126 2442 5129 2538
rect 5134 2472 5137 3058
rect 5142 2971 5145 3168
rect 5154 3048 5158 3051
rect 5142 2968 5153 2971
rect 5094 2348 5105 2351
rect 5094 2072 5097 2348
rect 5106 2338 5110 2341
rect 5086 1511 5089 1968
rect 5078 1508 5089 1511
rect 5046 1358 5054 1361
rect 5054 1272 5057 1358
rect 5058 1268 5065 1271
rect 5038 652 5041 728
rect 5054 542 5057 1228
rect 5062 982 5065 1268
rect 5062 742 5065 928
rect 5066 738 5073 741
rect 5070 222 5073 738
rect 5078 122 5081 1508
rect 5086 1492 5089 1498
rect 5094 1262 5097 2068
rect 5102 1532 5105 2008
rect 5110 1452 5113 2068
rect 5118 272 5121 1868
rect 5126 932 5129 2338
rect 5134 2282 5137 2428
rect 5142 2292 5145 2658
rect 5134 262 5137 2038
rect 5142 1912 5145 2278
rect 5150 2272 5153 2968
rect 5158 2552 5161 2968
rect 5174 2961 5177 3368
rect 5166 2958 5177 2961
rect 5166 2662 5169 2958
rect 5166 2642 5169 2648
rect 5158 2422 5161 2528
rect 5150 1932 5153 2258
rect 5106 188 5110 191
rect 5010 88 5014 91
rect 5142 62 5145 1878
rect 5150 1622 5153 1928
rect 5158 72 5161 2258
rect 5166 2052 5169 2638
rect 5174 2452 5177 2948
rect 5182 2672 5185 4498
rect 5190 3252 5193 3478
rect 5190 2762 5193 2768
rect 5186 2648 5190 2651
rect 5182 2431 5185 2488
rect 5174 2428 5185 2431
rect 5174 2102 5177 2428
rect 5166 2032 5169 2038
rect 5174 1982 5177 2078
rect 5166 1562 5169 1958
rect 5166 932 5169 938
rect 5174 152 5177 1938
rect 5182 1762 5185 2418
rect 5190 2062 5193 2068
rect 5182 852 5185 858
rect 5186 288 5190 291
rect 4690 58 4694 61
rect 4754 58 4758 61
rect 4042 48 4046 51
rect 4122 48 4126 51
rect 4554 48 4558 51
rect 4818 48 4822 51
rect 536 3 538 7
rect 542 3 545 7
rect 550 3 552 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1574 3 1576 7
rect 2584 3 2586 7
rect 2590 3 2593 7
rect 2598 3 2600 7
rect 3608 3 3610 7
rect 3614 3 3617 7
rect 3622 3 3624 7
rect 4632 3 4634 7
rect 4638 3 4641 7
rect 4646 3 4648 7
<< m5contact >>
rect 1050 4903 1054 4907
rect 1057 4903 1058 4907
rect 1058 4903 1061 4907
rect 2074 4903 2078 4907
rect 2081 4903 2082 4907
rect 2082 4903 2085 4907
rect 3098 4903 3102 4907
rect 3105 4903 3106 4907
rect 3106 4903 3109 4907
rect 4114 4903 4118 4907
rect 4121 4903 4122 4907
rect 4122 4903 4125 4907
rect 582 4858 586 4862
rect 538 4803 542 4807
rect 545 4803 546 4807
rect 546 4803 549 4807
rect 150 4648 154 4652
rect 134 3358 138 3362
rect 22 3148 26 3152
rect 422 4648 426 4652
rect 766 4858 770 4862
rect 670 4748 674 4752
rect 494 4688 498 4692
rect 318 4518 322 4522
rect 278 4348 282 4352
rect 262 4248 266 4252
rect 246 3478 250 3482
rect 166 3328 170 3332
rect 302 4108 306 4112
rect 270 3958 274 3962
rect 278 3858 282 3862
rect 318 4058 322 4062
rect 174 3068 178 3072
rect 198 2948 202 2952
rect 214 2678 218 2682
rect 14 2548 18 2552
rect 6 2518 10 2522
rect 118 2488 122 2492
rect 14 2438 18 2442
rect 14 2348 18 2352
rect 14 2328 18 2332
rect 94 2318 98 2322
rect 94 2128 98 2132
rect 78 2088 82 2092
rect 166 2088 170 2092
rect 134 1158 138 1162
rect 134 868 138 872
rect 270 3278 274 3282
rect 310 2758 314 2762
rect 270 2258 274 2262
rect 262 2218 266 2222
rect 238 1788 242 1792
rect 222 1468 226 1472
rect 214 1158 218 1162
rect 222 1058 226 1062
rect 198 548 202 552
rect 190 328 194 332
rect 134 268 138 272
rect 222 148 226 152
rect 294 1948 298 1952
rect 294 1418 298 1422
rect 342 3558 346 3562
rect 334 3258 338 3262
rect 326 2618 330 2622
rect 366 4178 370 4182
rect 422 4138 426 4142
rect 390 4078 394 4082
rect 382 4018 386 4022
rect 382 3738 386 3742
rect 358 3558 362 3562
rect 414 3868 418 3872
rect 374 3158 378 3162
rect 374 2758 378 2762
rect 366 2688 370 2692
rect 350 2458 354 2462
rect 382 2278 386 2282
rect 382 2148 386 2152
rect 334 2138 338 2142
rect 382 2048 386 2052
rect 390 1888 394 1892
rect 406 2848 410 2852
rect 430 3318 434 3322
rect 414 2778 418 2782
rect 538 4603 542 4607
rect 545 4603 546 4607
rect 546 4603 549 4607
rect 538 4403 542 4407
rect 545 4403 546 4407
rect 546 4403 549 4407
rect 550 4318 554 4322
rect 538 4203 542 4207
rect 545 4203 546 4207
rect 546 4203 549 4207
rect 478 3678 482 3682
rect 446 3478 450 3482
rect 438 2668 442 2672
rect 414 2548 418 2552
rect 366 1668 370 1672
rect 382 1428 386 1432
rect 406 1618 410 1622
rect 398 1418 402 1422
rect 358 1318 362 1322
rect 382 1258 386 1262
rect 350 978 354 982
rect 302 768 306 772
rect 414 1528 418 1532
rect 470 3188 474 3192
rect 630 4448 634 4452
rect 630 4288 634 4292
rect 566 4028 570 4032
rect 538 4003 542 4007
rect 545 4003 546 4007
rect 546 4003 549 4007
rect 538 3803 542 3807
rect 545 3803 546 3807
rect 546 3803 549 3807
rect 538 3603 542 3607
rect 545 3603 546 3607
rect 546 3603 549 3607
rect 502 3498 506 3502
rect 538 3403 542 3407
rect 545 3403 546 3407
rect 546 3403 549 3407
rect 550 3358 554 3362
rect 518 3328 522 3332
rect 518 3318 522 3322
rect 538 3203 542 3207
rect 545 3203 546 3207
rect 546 3203 549 3207
rect 510 2758 514 2762
rect 494 2568 498 2572
rect 486 2388 490 2392
rect 538 3003 542 3007
rect 545 3003 546 3007
rect 546 3003 549 3007
rect 518 2368 522 2372
rect 478 2268 482 2272
rect 470 2218 474 2222
rect 478 2048 482 2052
rect 462 1828 466 1832
rect 454 1628 458 1632
rect 430 1448 434 1452
rect 422 1078 426 1082
rect 350 468 354 472
rect 350 348 354 352
rect 446 1308 450 1312
rect 470 1248 474 1252
rect 470 1158 474 1162
rect 486 1448 490 1452
rect 462 868 466 872
rect 422 468 426 472
rect 574 3198 578 3202
rect 558 2828 562 2832
rect 538 2803 542 2807
rect 545 2803 546 2807
rect 546 2803 549 2807
rect 538 2603 542 2607
rect 545 2603 546 2607
rect 546 2603 549 2607
rect 542 2478 546 2482
rect 538 2403 542 2407
rect 545 2403 546 2407
rect 546 2403 549 2407
rect 538 2203 542 2207
rect 545 2203 546 2207
rect 546 2203 549 2207
rect 574 2868 578 2872
rect 590 3968 594 3972
rect 574 2688 578 2692
rect 582 2658 586 2662
rect 614 3548 618 3552
rect 598 2608 602 2612
rect 574 2578 578 2582
rect 574 2528 578 2532
rect 538 2003 542 2007
rect 545 2003 546 2007
rect 546 2003 549 2007
rect 538 1803 542 1807
rect 545 1803 546 1807
rect 546 1803 549 1807
rect 538 1603 542 1607
rect 545 1603 546 1607
rect 546 1603 549 1607
rect 590 2458 594 2462
rect 654 4468 658 4472
rect 646 3328 650 3332
rect 710 4328 714 4332
rect 670 3838 674 3842
rect 670 3698 674 3702
rect 678 3578 682 3582
rect 686 3548 690 3552
rect 678 3448 682 3452
rect 662 3278 666 3282
rect 670 3278 674 3282
rect 694 3358 698 3362
rect 678 3138 682 3142
rect 662 2998 666 3002
rect 694 2948 698 2952
rect 646 2638 650 2642
rect 614 2408 618 2412
rect 630 2498 634 2502
rect 590 2178 594 2182
rect 622 2388 626 2392
rect 630 2198 634 2202
rect 678 2748 682 2752
rect 686 2678 690 2682
rect 662 2418 666 2422
rect 654 2278 658 2282
rect 638 2158 642 2162
rect 654 2158 658 2162
rect 622 2068 626 2072
rect 614 1958 618 1962
rect 606 1888 610 1892
rect 590 1678 594 1682
rect 574 1668 578 1672
rect 538 1403 542 1407
rect 545 1403 546 1407
rect 546 1403 549 1407
rect 502 1388 506 1392
rect 574 1348 578 1352
rect 598 1418 602 1422
rect 622 1398 626 1402
rect 646 1898 650 1902
rect 662 2038 666 2042
rect 638 1358 642 1362
rect 630 1338 634 1342
rect 598 1268 602 1272
rect 590 1248 594 1252
rect 538 1203 542 1207
rect 545 1203 546 1207
rect 546 1203 549 1207
rect 538 1003 542 1007
rect 545 1003 546 1007
rect 546 1003 549 1007
rect 510 858 514 862
rect 538 803 542 807
rect 545 803 546 807
rect 546 803 549 807
rect 622 1128 626 1132
rect 598 978 602 982
rect 590 838 594 842
rect 538 603 542 607
rect 545 603 546 607
rect 546 603 549 607
rect 590 558 594 562
rect 566 518 570 522
rect 538 403 542 407
rect 545 403 546 407
rect 546 403 549 407
rect 742 4538 746 4542
rect 718 3938 722 3942
rect 862 4528 866 4532
rect 766 3818 770 3822
rect 718 3418 722 3422
rect 726 3408 730 3412
rect 726 3358 730 3362
rect 710 3148 714 3152
rect 710 3118 714 3122
rect 710 3008 714 3012
rect 694 2628 698 2632
rect 678 2038 682 2042
rect 670 1708 674 1712
rect 670 1648 674 1652
rect 702 2478 706 2482
rect 694 2138 698 2142
rect 686 2028 690 2032
rect 702 1718 706 1722
rect 718 1708 722 1712
rect 734 3148 738 3152
rect 766 3238 770 3242
rect 750 3218 754 3222
rect 774 3178 778 3182
rect 774 3158 778 3162
rect 758 3088 762 3092
rect 774 3058 778 3062
rect 774 2968 778 2972
rect 742 2748 746 2752
rect 758 2868 762 2872
rect 814 4258 818 4262
rect 854 4238 858 4242
rect 790 4148 794 4152
rect 798 4068 802 4072
rect 878 4028 882 4032
rect 798 2938 802 2942
rect 790 2848 794 2852
rect 782 2818 786 2822
rect 758 2668 762 2672
rect 742 1998 746 2002
rect 726 1538 730 1542
rect 718 1348 722 1352
rect 638 538 642 542
rect 638 528 642 532
rect 622 458 626 462
rect 598 328 602 332
rect 446 288 450 292
rect 454 268 458 272
rect 550 238 554 242
rect 538 203 542 207
rect 545 203 546 207
rect 546 203 549 207
rect 534 148 538 152
rect 694 988 698 992
rect 686 518 690 522
rect 710 938 714 942
rect 702 718 706 722
rect 710 618 714 622
rect 782 2578 786 2582
rect 782 2558 786 2562
rect 814 3128 818 3132
rect 814 3108 818 3112
rect 830 3568 834 3572
rect 894 4128 898 4132
rect 902 4048 906 4052
rect 910 3898 914 3902
rect 862 3448 866 3452
rect 854 3228 858 3232
rect 846 3068 850 3072
rect 830 2888 834 2892
rect 822 2778 826 2782
rect 838 2678 842 2682
rect 838 2658 842 2662
rect 806 2498 810 2502
rect 806 2468 810 2472
rect 822 2578 826 2582
rect 814 2328 818 2332
rect 790 1898 794 1902
rect 758 1748 762 1752
rect 766 1668 770 1672
rect 782 1678 786 1682
rect 766 1478 770 1482
rect 750 1318 754 1322
rect 750 1118 754 1122
rect 726 848 730 852
rect 726 768 730 772
rect 742 718 746 722
rect 758 618 762 622
rect 782 1258 786 1262
rect 870 2938 874 2942
rect 846 2528 850 2532
rect 830 2428 834 2432
rect 838 2168 842 2172
rect 806 1438 810 1442
rect 806 1388 810 1392
rect 790 1068 794 1072
rect 870 2448 874 2452
rect 886 3268 890 3272
rect 854 2188 858 2192
rect 878 2148 882 2152
rect 870 2108 874 2112
rect 862 1928 866 1932
rect 854 1798 858 1802
rect 822 1638 826 1642
rect 846 1578 850 1582
rect 822 1438 826 1442
rect 830 1408 834 1412
rect 878 1958 882 1962
rect 838 1228 842 1232
rect 838 1148 842 1152
rect 926 4038 930 4042
rect 918 3228 922 3232
rect 910 3218 914 3222
rect 894 2678 898 2682
rect 894 2408 898 2412
rect 894 2388 898 2392
rect 894 2228 898 2232
rect 886 1548 890 1552
rect 870 1118 874 1122
rect 854 1078 858 1082
rect 862 1058 866 1062
rect 814 988 818 992
rect 814 978 818 982
rect 798 958 802 962
rect 782 868 786 872
rect 782 348 786 352
rect 822 748 826 752
rect 886 1328 890 1332
rect 1246 4858 1250 4862
rect 1542 4858 1546 4862
rect 1222 4748 1226 4752
rect 1050 4703 1054 4707
rect 1057 4703 1058 4707
rect 1058 4703 1061 4707
rect 1150 4678 1154 4682
rect 1206 4688 1210 4692
rect 1198 4658 1202 4662
rect 966 4108 970 4112
rect 966 4068 970 4072
rect 942 3288 946 3292
rect 958 3418 962 3422
rect 1050 4503 1054 4507
rect 1057 4503 1058 4507
rect 1058 4503 1061 4507
rect 998 4328 1002 4332
rect 1006 4238 1010 4242
rect 998 3668 1002 3672
rect 1022 3988 1026 3992
rect 1006 3618 1010 3622
rect 998 3458 1002 3462
rect 990 3328 994 3332
rect 950 3208 954 3212
rect 918 2958 922 2962
rect 918 2488 922 2492
rect 918 2418 922 2422
rect 910 2148 914 2152
rect 910 2008 914 2012
rect 902 1148 906 1152
rect 894 1138 898 1142
rect 886 988 890 992
rect 886 838 890 842
rect 934 3028 938 3032
rect 934 2848 938 2852
rect 934 2618 938 2622
rect 950 3028 954 3032
rect 982 3288 986 3292
rect 998 3188 1002 3192
rect 990 3158 994 3162
rect 990 3138 994 3142
rect 982 3108 986 3112
rect 974 3048 978 3052
rect 966 2928 970 2932
rect 950 2728 954 2732
rect 942 2378 946 2382
rect 926 2158 930 2162
rect 942 2248 946 2252
rect 950 2158 954 2162
rect 958 2158 962 2162
rect 926 1668 930 1672
rect 942 1938 946 1942
rect 958 2138 962 2142
rect 982 2088 986 2092
rect 982 2018 986 2022
rect 998 3078 1002 3082
rect 1050 4303 1054 4307
rect 1057 4303 1058 4307
rect 1058 4303 1061 4307
rect 1086 4358 1090 4362
rect 1050 4103 1054 4107
rect 1057 4103 1058 4107
rect 1058 4103 1061 4107
rect 1050 3903 1054 3907
rect 1057 3903 1058 3907
rect 1058 3903 1061 3907
rect 1078 3978 1082 3982
rect 1050 3703 1054 3707
rect 1057 3703 1058 3707
rect 1058 3703 1061 3707
rect 1030 3698 1034 3702
rect 1022 3538 1026 3542
rect 1014 2978 1018 2982
rect 1006 2868 1010 2872
rect 1070 3598 1074 3602
rect 1050 3503 1054 3507
rect 1057 3503 1058 3507
rect 1058 3503 1061 3507
rect 1038 3468 1042 3472
rect 1050 3303 1054 3307
rect 1057 3303 1058 3307
rect 1058 3303 1061 3307
rect 1050 3103 1054 3107
rect 1057 3103 1058 3107
rect 1058 3103 1061 3107
rect 1038 2948 1042 2952
rect 1050 2903 1054 2907
rect 1057 2903 1058 2907
rect 1058 2903 1061 2907
rect 1030 2898 1034 2902
rect 1022 2878 1026 2882
rect 1014 2838 1018 2842
rect 1006 2828 1010 2832
rect 998 2678 1002 2682
rect 998 2648 1002 2652
rect 998 2638 1002 2642
rect 1038 2818 1042 2822
rect 1030 2688 1034 2692
rect 1014 2488 1018 2492
rect 1014 2478 1018 2482
rect 1006 2208 1010 2212
rect 950 1678 954 1682
rect 950 1668 954 1672
rect 958 1548 962 1552
rect 942 1518 946 1522
rect 974 1918 978 1922
rect 990 1858 994 1862
rect 950 1408 954 1412
rect 966 1408 970 1412
rect 934 1358 938 1362
rect 934 1348 938 1352
rect 918 1088 922 1092
rect 918 808 922 812
rect 910 768 914 772
rect 870 588 874 592
rect 902 558 906 562
rect 862 548 866 552
rect 854 518 858 522
rect 838 458 842 462
rect 870 338 874 342
rect 862 288 866 292
rect 926 558 930 562
rect 958 1158 962 1162
rect 966 1058 970 1062
rect 1006 1838 1010 1842
rect 990 1538 994 1542
rect 998 1268 1002 1272
rect 998 1128 1002 1132
rect 990 938 994 942
rect 982 878 986 882
rect 966 858 970 862
rect 966 728 970 732
rect 974 718 978 722
rect 926 548 930 552
rect 934 528 938 532
rect 958 468 962 472
rect 990 828 994 832
rect 1030 2478 1034 2482
rect 1030 2118 1034 2122
rect 1050 2703 1054 2707
rect 1057 2703 1058 2707
rect 1058 2703 1061 2707
rect 1102 3928 1106 3932
rect 1094 3918 1098 3922
rect 1166 4458 1170 4462
rect 1150 4288 1154 4292
rect 1174 4278 1178 4282
rect 1094 3328 1098 3332
rect 1094 3188 1098 3192
rect 1086 2888 1090 2892
rect 1050 2503 1054 2507
rect 1057 2503 1058 2507
rect 1058 2503 1061 2507
rect 1050 2303 1054 2307
rect 1057 2303 1058 2307
rect 1058 2303 1061 2307
rect 1070 2148 1074 2152
rect 1050 2103 1054 2107
rect 1057 2103 1058 2107
rect 1058 2103 1061 2107
rect 1110 3628 1114 3632
rect 1158 4068 1162 4072
rect 1158 3968 1162 3972
rect 1150 3878 1154 3882
rect 1126 3638 1130 3642
rect 1118 3488 1122 3492
rect 1142 3648 1146 3652
rect 1190 4518 1194 4522
rect 1182 3968 1186 3972
rect 1150 3428 1154 3432
rect 1182 3738 1186 3742
rect 1142 3408 1146 3412
rect 1134 3228 1138 3232
rect 1126 3168 1130 3172
rect 1134 3158 1138 3162
rect 1182 3328 1186 3332
rect 1182 3298 1186 3302
rect 1214 4078 1218 4082
rect 1230 4118 1234 4122
rect 1230 4078 1234 4082
rect 1214 3968 1218 3972
rect 1222 3968 1226 3972
rect 1214 3958 1218 3962
rect 1198 3668 1202 3672
rect 1158 3168 1162 3172
rect 1158 3158 1162 3162
rect 1150 3138 1154 3142
rect 1174 3138 1178 3142
rect 1142 2978 1146 2982
rect 1126 2938 1130 2942
rect 1118 2468 1122 2472
rect 1110 2418 1114 2422
rect 1046 2078 1050 2082
rect 1094 2058 1098 2062
rect 1070 1968 1074 1972
rect 1050 1903 1054 1907
rect 1057 1903 1058 1907
rect 1058 1903 1061 1907
rect 1030 1738 1034 1742
rect 1050 1703 1054 1707
rect 1057 1703 1058 1707
rect 1058 1703 1061 1707
rect 1086 1888 1090 1892
rect 1078 1868 1082 1872
rect 1050 1503 1054 1507
rect 1057 1503 1058 1507
rect 1058 1503 1061 1507
rect 1038 1308 1042 1312
rect 1050 1303 1054 1307
rect 1057 1303 1058 1307
rect 1058 1303 1061 1307
rect 1022 1178 1026 1182
rect 1030 1148 1034 1152
rect 1022 1118 1026 1122
rect 1030 1028 1034 1032
rect 1046 1128 1050 1132
rect 1050 1103 1054 1107
rect 1057 1103 1058 1107
rect 1058 1103 1061 1107
rect 1150 2888 1154 2892
rect 1158 2598 1162 2602
rect 1150 2578 1154 2582
rect 1158 2558 1162 2562
rect 1134 2238 1138 2242
rect 1118 2138 1122 2142
rect 1118 2048 1122 2052
rect 1110 2028 1114 2032
rect 1102 1988 1106 1992
rect 1142 1978 1146 1982
rect 1158 2378 1162 2382
rect 1206 3308 1210 3312
rect 1198 3168 1202 3172
rect 1190 3018 1194 3022
rect 1182 2918 1186 2922
rect 1182 2898 1186 2902
rect 1182 2668 1186 2672
rect 1278 4528 1282 4532
rect 1254 4028 1258 4032
rect 1270 4028 1274 4032
rect 1230 3598 1234 3602
rect 1222 2988 1226 2992
rect 1214 2858 1218 2862
rect 1286 3958 1290 3962
rect 1278 3888 1282 3892
rect 1262 3508 1266 3512
rect 1270 3458 1274 3462
rect 1270 3348 1274 3352
rect 1254 3328 1258 3332
rect 1246 2998 1250 3002
rect 1238 2928 1242 2932
rect 1222 2638 1226 2642
rect 1206 2598 1210 2602
rect 1206 2548 1210 2552
rect 1174 2458 1178 2462
rect 1174 2398 1178 2402
rect 1190 2308 1194 2312
rect 1174 2168 1178 2172
rect 1190 2078 1194 2082
rect 1134 1948 1138 1952
rect 1150 1948 1154 1952
rect 1118 1738 1122 1742
rect 1102 1728 1106 1732
rect 1094 1628 1098 1632
rect 1086 1588 1090 1592
rect 1094 1588 1098 1592
rect 1078 1568 1082 1572
rect 1142 1568 1146 1572
rect 1102 1318 1106 1322
rect 1046 1028 1050 1032
rect 1050 903 1054 907
rect 1057 903 1058 907
rect 1058 903 1061 907
rect 1062 758 1066 762
rect 1046 738 1050 742
rect 1050 703 1054 707
rect 1057 703 1058 707
rect 1058 703 1061 707
rect 1134 1408 1138 1412
rect 1110 1238 1114 1242
rect 1094 1058 1098 1062
rect 1086 918 1090 922
rect 1086 848 1090 852
rect 1094 728 1098 732
rect 1070 568 1074 572
rect 1070 518 1074 522
rect 1050 503 1054 507
rect 1057 503 1058 507
rect 1058 503 1061 507
rect 1038 478 1042 482
rect 1126 1268 1130 1272
rect 1102 638 1106 642
rect 1158 1928 1162 1932
rect 1182 2008 1186 2012
rect 1174 1878 1178 1882
rect 1166 1818 1170 1822
rect 1174 1748 1178 1752
rect 1182 1698 1186 1702
rect 1158 1678 1162 1682
rect 1174 1568 1178 1572
rect 1174 1468 1178 1472
rect 1166 1438 1170 1442
rect 1246 2658 1250 2662
rect 1254 2628 1258 2632
rect 1246 2558 1250 2562
rect 1230 2548 1234 2552
rect 1230 2508 1234 2512
rect 1230 2488 1234 2492
rect 1214 2418 1218 2422
rect 1230 2418 1234 2422
rect 1222 2358 1226 2362
rect 1230 2348 1234 2352
rect 1214 2278 1218 2282
rect 1214 1748 1218 1752
rect 1198 1468 1202 1472
rect 1190 1458 1194 1462
rect 1190 1438 1194 1442
rect 1198 1438 1202 1442
rect 1134 518 1138 522
rect 1198 1368 1202 1372
rect 1198 1288 1202 1292
rect 1198 1258 1202 1262
rect 1198 1208 1202 1212
rect 1214 1538 1218 1542
rect 1230 1878 1234 1882
rect 1270 2498 1274 2502
rect 1254 2438 1258 2442
rect 1246 2358 1250 2362
rect 1262 2348 1266 2352
rect 1254 2288 1258 2292
rect 1246 2268 1250 2272
rect 1254 2268 1258 2272
rect 1230 1718 1234 1722
rect 1238 1708 1242 1712
rect 1222 1478 1226 1482
rect 1230 1448 1234 1452
rect 1214 1428 1218 1432
rect 1230 1428 1234 1432
rect 1246 1648 1250 1652
rect 1230 1358 1234 1362
rect 1238 1328 1242 1332
rect 1350 4748 1354 4752
rect 1310 4638 1314 4642
rect 1334 4678 1338 4682
rect 1382 4658 1386 4662
rect 1382 4548 1386 4552
rect 1374 4168 1378 4172
rect 1310 3708 1314 3712
rect 1318 3598 1322 3602
rect 1310 3568 1314 3572
rect 1302 3538 1306 3542
rect 1318 3548 1322 3552
rect 1294 3338 1298 3342
rect 1294 3308 1298 3312
rect 1294 3038 1298 3042
rect 1286 2908 1290 2912
rect 1326 3538 1330 3542
rect 1326 3478 1330 3482
rect 1358 3678 1362 3682
rect 1334 3428 1338 3432
rect 1562 4803 1566 4807
rect 1569 4803 1570 4807
rect 1570 4803 1573 4807
rect 1502 4748 1506 4752
rect 1630 4748 1634 4752
rect 1622 4738 1626 4742
rect 1542 4648 1546 4652
rect 1494 4538 1498 4542
rect 1446 4528 1450 4532
rect 1454 4418 1458 4422
rect 1462 4338 1466 4342
rect 1494 4318 1498 4322
rect 1414 4228 1418 4232
rect 1398 4148 1402 4152
rect 1406 4148 1410 4152
rect 1406 4058 1410 4062
rect 1374 3418 1378 3422
rect 1350 3308 1354 3312
rect 1326 3218 1330 3222
rect 1310 2958 1314 2962
rect 1318 2958 1322 2962
rect 1302 2948 1306 2952
rect 1310 2938 1314 2942
rect 1310 2888 1314 2892
rect 1302 2678 1306 2682
rect 1286 2568 1290 2572
rect 1278 2438 1282 2442
rect 1278 2368 1282 2372
rect 1294 2338 1298 2342
rect 1270 2068 1274 2072
rect 1286 2068 1290 2072
rect 1278 1968 1282 1972
rect 1286 1968 1290 1972
rect 1270 1698 1274 1702
rect 1270 1648 1274 1652
rect 1262 1368 1266 1372
rect 1246 1318 1250 1322
rect 1230 1308 1234 1312
rect 1214 1148 1218 1152
rect 1190 528 1194 532
rect 1238 1138 1242 1142
rect 1238 818 1242 822
rect 1246 648 1250 652
rect 1390 3458 1394 3462
rect 1406 3628 1410 3632
rect 1534 4528 1538 4532
rect 1562 4603 1566 4607
rect 1569 4603 1570 4607
rect 1570 4603 1573 4607
rect 1574 4518 1578 4522
rect 1562 4403 1566 4407
rect 1569 4403 1570 4407
rect 1570 4403 1573 4407
rect 1598 4448 1602 4452
rect 1590 4418 1594 4422
rect 1494 4158 1498 4162
rect 1510 4138 1514 4142
rect 1446 3938 1450 3942
rect 1446 3908 1450 3912
rect 1438 3718 1442 3722
rect 1478 3898 1482 3902
rect 1422 3548 1426 3552
rect 1414 3518 1418 3522
rect 1430 3518 1434 3522
rect 1454 3498 1458 3502
rect 1414 3478 1418 3482
rect 1398 3438 1402 3442
rect 1382 3168 1386 3172
rect 1374 3118 1378 3122
rect 1366 3108 1370 3112
rect 1350 3028 1354 3032
rect 1334 2988 1338 2992
rect 1318 2568 1322 2572
rect 1318 2538 1322 2542
rect 1350 2938 1354 2942
rect 1342 2768 1346 2772
rect 1374 2978 1378 2982
rect 1366 2668 1370 2672
rect 1366 2638 1370 2642
rect 1326 2468 1330 2472
rect 1318 2418 1322 2422
rect 1318 2388 1322 2392
rect 1318 2138 1322 2142
rect 1358 2458 1362 2462
rect 1350 2438 1354 2442
rect 1334 2218 1338 2222
rect 1326 2108 1330 2112
rect 1310 1928 1314 1932
rect 1302 1858 1306 1862
rect 1302 1788 1306 1792
rect 1302 1518 1306 1522
rect 1318 1838 1322 1842
rect 1334 2088 1338 2092
rect 1406 3328 1410 3332
rect 1470 3468 1474 3472
rect 1414 3058 1418 3062
rect 1390 2978 1394 2982
rect 1374 2498 1378 2502
rect 1430 2978 1434 2982
rect 1422 2788 1426 2792
rect 1398 2678 1402 2682
rect 1462 3328 1466 3332
rect 1454 3218 1458 3222
rect 1446 3008 1450 3012
rect 1438 2948 1442 2952
rect 1494 3538 1498 3542
rect 1486 3528 1490 3532
rect 1526 4038 1530 4042
rect 1510 3718 1514 3722
rect 1518 3458 1522 3462
rect 1510 3418 1514 3422
rect 1486 3398 1490 3402
rect 1486 3358 1490 3362
rect 1502 3298 1506 3302
rect 1494 3248 1498 3252
rect 1478 3228 1482 3232
rect 1494 3198 1498 3202
rect 1494 3148 1498 3152
rect 1486 3138 1490 3142
rect 1438 2808 1442 2812
rect 1422 2708 1426 2712
rect 1414 2688 1418 2692
rect 1414 2588 1418 2592
rect 1462 2838 1466 2842
rect 1454 2758 1458 2762
rect 1430 2598 1434 2602
rect 1478 2638 1482 2642
rect 1398 2548 1402 2552
rect 1446 2548 1450 2552
rect 1390 2458 1394 2462
rect 1358 2188 1362 2192
rect 1350 1968 1354 1972
rect 1342 1948 1346 1952
rect 1326 1828 1330 1832
rect 1326 1648 1330 1652
rect 1326 1558 1330 1562
rect 1326 1448 1330 1452
rect 1358 1768 1362 1772
rect 1358 1488 1362 1492
rect 1342 1468 1346 1472
rect 1342 1318 1346 1322
rect 1326 1258 1330 1262
rect 1334 1188 1338 1192
rect 1350 1308 1354 1312
rect 1374 1578 1378 1582
rect 1366 1358 1370 1362
rect 1254 538 1258 542
rect 1286 678 1290 682
rect 1050 303 1054 307
rect 1057 303 1058 307
rect 1058 303 1061 307
rect 1078 278 1082 282
rect 1062 238 1066 242
rect 1270 378 1274 382
rect 1326 368 1330 372
rect 1350 338 1354 342
rect 1390 2148 1394 2152
rect 1406 2318 1410 2322
rect 1406 2308 1410 2312
rect 1398 2118 1402 2122
rect 1398 1878 1402 1882
rect 1398 1868 1402 1872
rect 1390 1508 1394 1512
rect 1390 1378 1394 1382
rect 1430 2408 1434 2412
rect 1430 2388 1434 2392
rect 1430 2048 1434 2052
rect 1422 1928 1426 1932
rect 1414 1918 1418 1922
rect 1430 1798 1434 1802
rect 1430 1748 1434 1752
rect 1406 1578 1410 1582
rect 1422 1528 1426 1532
rect 1422 1468 1426 1472
rect 1422 1408 1426 1412
rect 1398 1348 1402 1352
rect 1382 1298 1386 1302
rect 1406 1248 1410 1252
rect 1414 968 1418 972
rect 1462 2458 1466 2462
rect 1454 2438 1458 2442
rect 1462 2358 1466 2362
rect 1462 2248 1466 2252
rect 1454 1748 1458 1752
rect 1470 2138 1474 2142
rect 1446 1658 1450 1662
rect 1430 838 1434 842
rect 1414 808 1418 812
rect 1422 778 1426 782
rect 1494 2818 1498 2822
rect 1486 2628 1490 2632
rect 1562 4203 1566 4207
rect 1569 4203 1570 4207
rect 1570 4203 1573 4207
rect 1562 4003 1566 4007
rect 1569 4003 1570 4007
rect 1570 4003 1573 4007
rect 1534 3678 1538 3682
rect 1534 3468 1538 3472
rect 1518 2978 1522 2982
rect 1510 2958 1514 2962
rect 1510 2928 1514 2932
rect 1518 2918 1522 2922
rect 1510 2838 1514 2842
rect 1510 2658 1514 2662
rect 1502 2648 1506 2652
rect 1510 2648 1514 2652
rect 1502 2338 1506 2342
rect 1494 2318 1498 2322
rect 1486 2308 1490 2312
rect 1486 2038 1490 2042
rect 1510 2278 1514 2282
rect 1502 2198 1506 2202
rect 1502 2078 1506 2082
rect 1494 1998 1498 2002
rect 1486 1988 1490 1992
rect 1502 1958 1506 1962
rect 1510 1938 1514 1942
rect 1478 1798 1482 1802
rect 1478 1738 1482 1742
rect 1478 1718 1482 1722
rect 1494 1748 1498 1752
rect 1534 3048 1538 3052
rect 1526 2898 1530 2902
rect 1566 3868 1570 3872
rect 1630 4538 1634 4542
rect 1558 3848 1562 3852
rect 1562 3803 1566 3807
rect 1569 3803 1570 3807
rect 1570 3803 1573 3807
rect 1590 3708 1594 3712
rect 1598 3688 1602 3692
rect 1622 4048 1626 4052
rect 1630 4048 1634 4052
rect 1562 3603 1566 3607
rect 1569 3603 1570 3607
rect 1570 3603 1573 3607
rect 1606 3588 1610 3592
rect 1562 3403 1566 3407
rect 1569 3403 1570 3407
rect 1570 3403 1573 3407
rect 1562 3203 1566 3207
rect 1569 3203 1570 3207
rect 1570 3203 1573 3207
rect 1598 3508 1602 3512
rect 1590 3268 1594 3272
rect 1582 3198 1586 3202
rect 1550 3158 1554 3162
rect 1630 3578 1634 3582
rect 1638 3558 1642 3562
rect 1630 3548 1634 3552
rect 1630 3468 1634 3472
rect 1622 3458 1626 3462
rect 1562 3003 1566 3007
rect 1569 3003 1570 3007
rect 1570 3003 1573 3007
rect 1582 2998 1586 3002
rect 1534 2868 1538 2872
rect 1550 2808 1554 2812
rect 1562 2803 1566 2807
rect 1569 2803 1570 2807
rect 1570 2803 1573 2807
rect 1582 2798 1586 2802
rect 1566 2618 1570 2622
rect 1550 2608 1554 2612
rect 1526 2588 1530 2592
rect 1542 2568 1546 2572
rect 1526 2538 1530 2542
rect 1534 2288 1538 2292
rect 1534 1908 1538 1912
rect 1518 1868 1522 1872
rect 1510 1828 1514 1832
rect 1502 1738 1506 1742
rect 1534 1818 1538 1822
rect 1526 1758 1530 1762
rect 1518 1638 1522 1642
rect 1486 1548 1490 1552
rect 1562 2603 1566 2607
rect 1569 2603 1570 2607
rect 1570 2603 1573 2607
rect 1590 2608 1594 2612
rect 1590 2528 1594 2532
rect 1582 2458 1586 2462
rect 1582 2448 1586 2452
rect 1562 2403 1566 2407
rect 1569 2403 1570 2407
rect 1570 2403 1573 2407
rect 1630 3308 1634 3312
rect 1638 3278 1642 3282
rect 1630 3268 1634 3272
rect 1614 3048 1618 3052
rect 1622 2898 1626 2902
rect 1630 2888 1634 2892
rect 1606 2838 1610 2842
rect 1630 2838 1634 2842
rect 1622 2758 1626 2762
rect 1630 2628 1634 2632
rect 1606 2438 1610 2442
rect 1606 2408 1610 2412
rect 1606 2368 1610 2372
rect 1582 2218 1586 2222
rect 1562 2203 1566 2207
rect 1569 2203 1570 2207
rect 1570 2203 1573 2207
rect 1558 2128 1562 2132
rect 1582 2078 1586 2082
rect 1550 2058 1554 2062
rect 1550 2038 1554 2042
rect 1566 2028 1570 2032
rect 1562 2003 1566 2007
rect 1569 2003 1570 2007
rect 1570 2003 1573 2007
rect 1542 1678 1546 1682
rect 1478 1488 1482 1492
rect 1502 1488 1506 1492
rect 1470 1438 1474 1442
rect 1446 1398 1450 1402
rect 1462 1278 1466 1282
rect 1446 1248 1450 1252
rect 1462 1218 1466 1222
rect 1454 1068 1458 1072
rect 1462 958 1466 962
rect 1414 768 1418 772
rect 1398 458 1402 462
rect 1398 388 1402 392
rect 1446 538 1450 542
rect 1422 358 1426 362
rect 1050 103 1054 107
rect 1057 103 1058 107
rect 1058 103 1061 107
rect 350 68 354 72
rect 974 68 978 72
rect 1478 1148 1482 1152
rect 1614 2288 1618 2292
rect 1622 2268 1626 2272
rect 1606 2258 1610 2262
rect 1654 3418 1658 3422
rect 1702 4738 1706 4742
rect 1678 4728 1682 4732
rect 1718 4528 1722 4532
rect 1678 4318 1682 4322
rect 1670 3748 1674 3752
rect 1670 3728 1674 3732
rect 1718 4148 1722 4152
rect 1710 4128 1714 4132
rect 1694 3748 1698 3752
rect 1670 3718 1674 3722
rect 1670 3598 1674 3602
rect 1686 3718 1690 3722
rect 1678 3468 1682 3472
rect 1646 2878 1650 2882
rect 1662 3088 1666 3092
rect 1750 4178 1754 4182
rect 1726 4068 1730 4072
rect 1718 3808 1722 3812
rect 1710 3768 1714 3772
rect 1686 3298 1690 3302
rect 1718 3688 1722 3692
rect 1710 3558 1714 3562
rect 1718 3458 1722 3462
rect 1710 3378 1714 3382
rect 1718 3358 1722 3362
rect 1702 3338 1706 3342
rect 1718 3338 1722 3342
rect 1694 3288 1698 3292
rect 1718 3208 1722 3212
rect 1670 3058 1674 3062
rect 1670 2958 1674 2962
rect 1662 2848 1666 2852
rect 1654 2698 1658 2702
rect 1646 2668 1650 2672
rect 1662 2628 1666 2632
rect 1646 2588 1650 2592
rect 1654 2518 1658 2522
rect 1654 2398 1658 2402
rect 1670 2388 1674 2392
rect 1654 2368 1658 2372
rect 1638 2178 1642 2182
rect 1630 2078 1634 2082
rect 1606 2008 1610 2012
rect 1606 1938 1610 1942
rect 1562 1803 1566 1807
rect 1569 1803 1570 1807
rect 1570 1803 1573 1807
rect 1562 1603 1566 1607
rect 1569 1603 1570 1607
rect 1570 1603 1573 1607
rect 1558 1558 1562 1562
rect 1574 1558 1578 1562
rect 1550 1448 1554 1452
rect 1566 1448 1570 1452
rect 1562 1403 1566 1407
rect 1569 1403 1570 1407
rect 1570 1403 1573 1407
rect 1558 1348 1562 1352
rect 1606 1868 1610 1872
rect 1590 1598 1594 1602
rect 1598 1548 1602 1552
rect 1562 1203 1566 1207
rect 1569 1203 1570 1207
rect 1570 1203 1573 1207
rect 1558 1118 1562 1122
rect 1542 1058 1546 1062
rect 1526 1038 1530 1042
rect 1486 948 1490 952
rect 1526 888 1530 892
rect 1582 1008 1586 1012
rect 1562 1003 1566 1007
rect 1569 1003 1570 1007
rect 1570 1003 1573 1007
rect 1562 803 1566 807
rect 1569 803 1570 807
rect 1570 803 1573 807
rect 1654 2218 1658 2222
rect 1742 3938 1746 3942
rect 1734 3678 1738 3682
rect 1726 3158 1730 3162
rect 1694 3078 1698 3082
rect 1694 3048 1698 3052
rect 1694 3028 1698 3032
rect 1694 2778 1698 2782
rect 1702 2738 1706 2742
rect 1718 2908 1722 2912
rect 2030 4728 2034 4732
rect 1750 3718 1754 3722
rect 1758 3688 1762 3692
rect 1750 3678 1754 3682
rect 1750 3618 1754 3622
rect 1822 4258 1826 4262
rect 1806 4018 1810 4022
rect 1766 3658 1770 3662
rect 1750 3578 1754 3582
rect 1758 3558 1762 3562
rect 1758 3548 1762 3552
rect 1742 3118 1746 3122
rect 1742 3108 1746 3112
rect 1734 3048 1738 3052
rect 1734 3038 1738 3042
rect 1726 2778 1730 2782
rect 1726 2748 1730 2752
rect 1694 2638 1698 2642
rect 1718 2608 1722 2612
rect 1710 2578 1714 2582
rect 1694 2558 1698 2562
rect 1686 2548 1690 2552
rect 1750 2748 1754 2752
rect 1750 2728 1754 2732
rect 1750 2628 1754 2632
rect 1750 2518 1754 2522
rect 1702 2438 1706 2442
rect 1734 2438 1738 2442
rect 1686 2418 1690 2422
rect 1670 2278 1674 2282
rect 1662 2088 1666 2092
rect 1622 1438 1626 1442
rect 1630 1438 1634 1442
rect 1646 1718 1650 1722
rect 1638 1398 1642 1402
rect 1646 1388 1650 1392
rect 1622 1198 1626 1202
rect 1598 978 1602 982
rect 1614 978 1618 982
rect 1694 2268 1698 2272
rect 1734 2388 1738 2392
rect 1710 2348 1714 2352
rect 1702 2238 1706 2242
rect 1694 2108 1698 2112
rect 1702 2098 1706 2102
rect 1694 2068 1698 2072
rect 1710 2038 1714 2042
rect 1678 2018 1682 2022
rect 1702 1998 1706 2002
rect 1670 1618 1674 1622
rect 1702 1578 1706 1582
rect 1678 1498 1682 1502
rect 1686 1498 1690 1502
rect 1646 1078 1650 1082
rect 1654 998 1658 1002
rect 1630 858 1634 862
rect 1646 848 1650 852
rect 1622 818 1626 822
rect 1606 798 1610 802
rect 1590 758 1594 762
rect 1478 738 1482 742
rect 1534 728 1538 732
rect 1454 148 1458 152
rect 1518 618 1522 622
rect 1518 448 1522 452
rect 1686 818 1690 822
rect 1686 788 1690 792
rect 1562 603 1566 607
rect 1569 603 1570 607
rect 1570 603 1573 607
rect 1542 568 1546 572
rect 1562 403 1566 407
rect 1569 403 1570 407
rect 1570 403 1573 407
rect 1526 278 1530 282
rect 1562 203 1566 207
rect 1569 203 1570 207
rect 1570 203 1573 207
rect 1486 148 1490 152
rect 1678 748 1682 752
rect 1750 2468 1754 2472
rect 1750 2398 1754 2402
rect 1750 2318 1754 2322
rect 1726 2108 1730 2112
rect 1750 2118 1754 2122
rect 1774 3528 1778 3532
rect 1782 3418 1786 3422
rect 1814 3828 1818 3832
rect 1814 3648 1818 3652
rect 1790 3038 1794 3042
rect 1846 4388 1850 4392
rect 2074 4703 2078 4707
rect 2081 4703 2082 4707
rect 2082 4703 2085 4707
rect 1958 4648 1962 4652
rect 1854 4368 1858 4372
rect 1838 3998 1842 4002
rect 1918 4478 1922 4482
rect 1862 3888 1866 3892
rect 1910 4188 1914 4192
rect 1902 4058 1906 4062
rect 1894 4028 1898 4032
rect 1894 3878 1898 3882
rect 1862 3798 1866 3802
rect 1854 3788 1858 3792
rect 1830 3498 1834 3502
rect 1822 3288 1826 3292
rect 1822 3278 1826 3282
rect 1806 2808 1810 2812
rect 1774 2768 1778 2772
rect 1766 2448 1770 2452
rect 1798 2608 1802 2612
rect 1798 2538 1802 2542
rect 1806 2478 1810 2482
rect 1774 2128 1778 2132
rect 1766 2058 1770 2062
rect 1742 2038 1746 2042
rect 1774 1938 1778 1942
rect 1758 1838 1762 1842
rect 1774 1878 1778 1882
rect 1734 1828 1738 1832
rect 1766 1828 1770 1832
rect 1750 1778 1754 1782
rect 1734 1758 1738 1762
rect 1758 1758 1762 1762
rect 1750 1698 1754 1702
rect 1718 1528 1722 1532
rect 1702 1478 1706 1482
rect 1702 1148 1706 1152
rect 1710 1108 1714 1112
rect 1678 658 1682 662
rect 1750 1638 1754 1642
rect 1790 2398 1794 2402
rect 1790 2148 1794 2152
rect 1806 2298 1810 2302
rect 1782 1758 1786 1762
rect 1774 1708 1778 1712
rect 1766 1508 1770 1512
rect 1710 688 1714 692
rect 1686 548 1690 552
rect 1694 368 1698 372
rect 1726 858 1730 862
rect 1830 2878 1834 2882
rect 1910 3758 1914 3762
rect 1862 3448 1866 3452
rect 1830 2578 1834 2582
rect 1854 2818 1858 2822
rect 1854 2678 1858 2682
rect 1822 2548 1826 2552
rect 1830 2478 1834 2482
rect 1822 2318 1826 2322
rect 1878 2928 1882 2932
rect 1870 2658 1874 2662
rect 1870 2618 1874 2622
rect 1838 2428 1842 2432
rect 1846 2428 1850 2432
rect 1830 2228 1834 2232
rect 1838 2218 1842 2222
rect 1838 2208 1842 2212
rect 1822 2178 1826 2182
rect 1846 2078 1850 2082
rect 1830 1948 1834 1952
rect 1822 1938 1826 1942
rect 1838 1898 1842 1902
rect 1806 1888 1810 1892
rect 1854 2028 1858 2032
rect 1806 1848 1810 1852
rect 1814 1718 1818 1722
rect 1822 1658 1826 1662
rect 1806 1618 1810 1622
rect 1814 1618 1818 1622
rect 1822 1618 1826 1622
rect 1782 1448 1786 1452
rect 1774 978 1778 982
rect 1758 648 1762 652
rect 1798 1408 1802 1412
rect 1798 1128 1802 1132
rect 1806 1038 1810 1042
rect 1838 1848 1842 1852
rect 1838 1758 1842 1762
rect 1902 3668 1906 3672
rect 1974 4378 1978 4382
rect 1966 4018 1970 4022
rect 1942 3638 1946 3642
rect 1926 3628 1930 3632
rect 1910 3218 1914 3222
rect 1910 3158 1914 3162
rect 1918 3118 1922 3122
rect 1910 2908 1914 2912
rect 1918 2768 1922 2772
rect 1902 2718 1906 2722
rect 1902 2698 1906 2702
rect 1886 2518 1890 2522
rect 1886 2498 1890 2502
rect 1886 2458 1890 2462
rect 1894 2458 1898 2462
rect 1894 2438 1898 2442
rect 1910 2438 1914 2442
rect 1910 2418 1914 2422
rect 1902 2408 1906 2412
rect 1950 3238 1954 3242
rect 1950 3138 1954 3142
rect 1942 3018 1946 3022
rect 1950 2998 1954 3002
rect 1942 2968 1946 2972
rect 1950 2928 1954 2932
rect 1934 2768 1938 2772
rect 1942 2728 1946 2732
rect 1934 2568 1938 2572
rect 1934 2478 1938 2482
rect 1926 2468 1930 2472
rect 1950 2568 1954 2572
rect 1966 3328 1970 3332
rect 2030 4468 2034 4472
rect 1982 3768 1986 3772
rect 2022 4038 2026 4042
rect 2006 3778 2010 3782
rect 1990 3718 1994 3722
rect 1990 3448 1994 3452
rect 1998 3248 2002 3252
rect 1974 3158 1978 3162
rect 1982 3158 1986 3162
rect 1974 3128 1978 3132
rect 1982 3118 1986 3122
rect 1974 3058 1978 3062
rect 1974 3028 1978 3032
rect 1966 2918 1970 2922
rect 1982 2998 1986 3002
rect 1974 2828 1978 2832
rect 1974 2818 1978 2822
rect 1966 2738 1970 2742
rect 1974 2678 1978 2682
rect 1958 2558 1962 2562
rect 1950 2538 1954 2542
rect 1966 2518 1970 2522
rect 1958 2508 1962 2512
rect 1942 2448 1946 2452
rect 1926 2438 1930 2442
rect 1910 2348 1914 2352
rect 1918 2318 1922 2322
rect 1878 2288 1882 2292
rect 1894 2278 1898 2282
rect 1910 2278 1914 2282
rect 1886 2208 1890 2212
rect 1878 2188 1882 2192
rect 1894 2168 1898 2172
rect 1910 2168 1914 2172
rect 1894 2148 1898 2152
rect 1886 2118 1890 2122
rect 1870 1798 1874 1802
rect 1870 1718 1874 1722
rect 1854 1688 1858 1692
rect 1838 1128 1842 1132
rect 1830 958 1834 962
rect 1822 888 1826 892
rect 1894 1848 1898 1852
rect 1886 1808 1890 1812
rect 1886 1738 1890 1742
rect 1934 2188 1938 2192
rect 1926 2158 1930 2162
rect 1966 2398 1970 2402
rect 1950 2318 1954 2322
rect 1958 2288 1962 2292
rect 1966 2278 1970 2282
rect 1950 2198 1954 2202
rect 1958 2178 1962 2182
rect 1958 2128 1962 2132
rect 1950 2108 1954 2112
rect 1958 2098 1962 2102
rect 1918 1888 1922 1892
rect 1878 1658 1882 1662
rect 1886 1588 1890 1592
rect 1886 1568 1890 1572
rect 1894 1468 1898 1472
rect 1878 1268 1882 1272
rect 1910 1668 1914 1672
rect 1934 1598 1938 1602
rect 1910 1518 1914 1522
rect 1902 1348 1906 1352
rect 1894 1248 1898 1252
rect 1902 1138 1906 1142
rect 1902 1038 1906 1042
rect 1878 1018 1882 1022
rect 1774 478 1778 482
rect 1750 378 1754 382
rect 1766 138 1770 142
rect 1966 1928 1970 1932
rect 1950 1568 1954 1572
rect 1958 1548 1962 1552
rect 1942 1508 1946 1512
rect 1958 1368 1962 1372
rect 1942 1298 1946 1302
rect 2074 4503 2078 4507
rect 2081 4503 2082 4507
rect 2082 4503 2085 4507
rect 2070 4448 2074 4452
rect 2074 4303 2078 4307
rect 2081 4303 2082 4307
rect 2082 4303 2085 4307
rect 2134 4278 2138 4282
rect 2134 4268 2138 4272
rect 2074 4103 2078 4107
rect 2081 4103 2082 4107
rect 2082 4103 2085 4107
rect 2030 3778 2034 3782
rect 2030 3748 2034 3752
rect 2030 3718 2034 3722
rect 2074 3903 2078 3907
rect 2081 3903 2082 3907
rect 2082 3903 2085 3907
rect 2062 3898 2066 3902
rect 2094 3708 2098 3712
rect 2074 3703 2078 3707
rect 2081 3703 2082 3707
rect 2082 3703 2085 3707
rect 2134 4048 2138 4052
rect 2054 3558 2058 3562
rect 2006 3088 2010 3092
rect 2022 3138 2026 3142
rect 2022 3128 2026 3132
rect 2006 2938 2010 2942
rect 1998 2758 2002 2762
rect 1990 2678 1994 2682
rect 1998 2488 2002 2492
rect 2014 2808 2018 2812
rect 2038 3358 2042 3362
rect 2074 3503 2078 3507
rect 2081 3503 2082 3507
rect 2082 3503 2085 3507
rect 2078 3448 2082 3452
rect 2046 3348 2050 3352
rect 2074 3303 2078 3307
rect 2081 3303 2082 3307
rect 2082 3303 2085 3307
rect 2126 3898 2130 3902
rect 2118 3458 2122 3462
rect 2102 3438 2106 3442
rect 2110 3438 2114 3442
rect 2126 3298 2130 3302
rect 2110 3268 2114 3272
rect 2126 3238 2130 3242
rect 2094 3178 2098 3182
rect 2062 3148 2066 3152
rect 2054 3118 2058 3122
rect 2074 3103 2078 3107
rect 2081 3103 2082 3107
rect 2082 3103 2085 3107
rect 2046 3068 2050 3072
rect 2038 2938 2042 2942
rect 2046 2908 2050 2912
rect 2062 3088 2066 3092
rect 2054 2888 2058 2892
rect 2046 2868 2050 2872
rect 2046 2848 2050 2852
rect 2014 2578 2018 2582
rect 2014 2518 2018 2522
rect 2006 2478 2010 2482
rect 2006 2438 2010 2442
rect 1990 2378 1994 2382
rect 2006 2348 2010 2352
rect 1998 2298 2002 2302
rect 1998 2238 2002 2242
rect 1990 2228 1994 2232
rect 1990 2208 1994 2212
rect 1990 1838 1994 1842
rect 1974 1478 1978 1482
rect 1942 828 1946 832
rect 1934 778 1938 782
rect 1934 718 1938 722
rect 1934 548 1938 552
rect 1926 448 1930 452
rect 2014 2028 2018 2032
rect 2014 1978 2018 1982
rect 2030 2108 2034 2112
rect 2054 2688 2058 2692
rect 2046 2668 2050 2672
rect 2074 2903 2078 2907
rect 2081 2903 2082 2907
rect 2082 2903 2085 2907
rect 2086 2788 2090 2792
rect 2102 3108 2106 3112
rect 2174 4348 2178 4352
rect 2166 3998 2170 4002
rect 2166 3928 2170 3932
rect 2150 3778 2154 3782
rect 2142 3318 2146 3322
rect 2102 3098 2106 3102
rect 2134 3098 2138 3102
rect 2126 2888 2130 2892
rect 2102 2828 2106 2832
rect 2118 2798 2122 2802
rect 2110 2778 2114 2782
rect 2094 2728 2098 2732
rect 2074 2703 2078 2707
rect 2081 2703 2082 2707
rect 2082 2703 2085 2707
rect 2086 2658 2090 2662
rect 2062 2618 2066 2622
rect 2046 2588 2050 2592
rect 2046 2558 2050 2562
rect 2046 2428 2050 2432
rect 2086 2568 2090 2572
rect 2070 2538 2074 2542
rect 2074 2503 2078 2507
rect 2081 2503 2082 2507
rect 2082 2503 2085 2507
rect 2062 2418 2066 2422
rect 2054 2388 2058 2392
rect 2046 2358 2050 2362
rect 2054 2308 2058 2312
rect 2086 2378 2090 2382
rect 2074 2303 2078 2307
rect 2081 2303 2082 2307
rect 2082 2303 2085 2307
rect 2046 2198 2050 2202
rect 2046 2078 2050 2082
rect 2102 2708 2106 2712
rect 2102 2328 2106 2332
rect 2070 2218 2074 2222
rect 2062 2208 2066 2212
rect 2062 2188 2066 2192
rect 2102 2168 2106 2172
rect 2074 2103 2078 2107
rect 2081 2103 2082 2107
rect 2082 2103 2085 2107
rect 2078 2078 2082 2082
rect 2054 2008 2058 2012
rect 2046 1898 2050 1902
rect 2022 1838 2026 1842
rect 2038 1738 2042 1742
rect 1990 1168 1994 1172
rect 1982 778 1986 782
rect 2022 1358 2026 1362
rect 2022 1328 2026 1332
rect 2014 1048 2018 1052
rect 1998 718 2002 722
rect 2006 678 2010 682
rect 2070 1978 2074 1982
rect 2118 2268 2122 2272
rect 2118 2248 2122 2252
rect 2118 2158 2122 2162
rect 2086 1968 2090 1972
rect 2094 1968 2098 1972
rect 2070 1928 2074 1932
rect 2062 1908 2066 1912
rect 2094 1908 2098 1912
rect 2074 1903 2078 1907
rect 2081 1903 2082 1907
rect 2082 1903 2085 1907
rect 2094 1898 2098 1902
rect 2062 1818 2066 1822
rect 2054 1548 2058 1552
rect 2046 1358 2050 1362
rect 2078 1798 2082 1802
rect 2070 1748 2074 1752
rect 2086 1748 2090 1752
rect 2074 1703 2078 1707
rect 2081 1703 2082 1707
rect 2082 1703 2085 1707
rect 2086 1678 2090 1682
rect 2102 1718 2106 1722
rect 2094 1558 2098 1562
rect 2074 1503 2078 1507
rect 2081 1503 2082 1507
rect 2082 1503 2085 1507
rect 2086 1398 2090 1402
rect 2074 1303 2078 1307
rect 2081 1303 2082 1307
rect 2082 1303 2085 1307
rect 2070 1268 2074 1272
rect 2086 1268 2090 1272
rect 2054 1138 2058 1142
rect 2046 1128 2050 1132
rect 2062 1118 2066 1122
rect 2046 888 2050 892
rect 2030 568 2034 572
rect 2014 388 2018 392
rect 1886 258 1890 262
rect 806 58 810 62
rect 934 58 938 62
rect 1926 138 1930 142
rect 2074 1103 2078 1107
rect 2081 1103 2082 1107
rect 2082 1103 2085 1107
rect 2118 2038 2122 2042
rect 2182 4308 2186 4312
rect 2182 4258 2186 4262
rect 2182 3928 2186 3932
rect 2182 3868 2186 3872
rect 2246 4518 2250 4522
rect 2254 4468 2258 4472
rect 2238 4458 2242 4462
rect 2270 4418 2274 4422
rect 2214 4098 2218 4102
rect 2222 4058 2226 4062
rect 2166 3498 2170 3502
rect 2158 3218 2162 3222
rect 2190 3238 2194 3242
rect 2182 3048 2186 3052
rect 2166 2998 2170 3002
rect 2174 2918 2178 2922
rect 2174 2898 2178 2902
rect 2150 2738 2154 2742
rect 2150 2658 2154 2662
rect 2142 2618 2146 2622
rect 2150 2608 2154 2612
rect 2150 2518 2154 2522
rect 2142 2298 2146 2302
rect 2166 2698 2170 2702
rect 2182 2498 2186 2502
rect 2174 2458 2178 2462
rect 2166 2398 2170 2402
rect 2174 2398 2178 2402
rect 2150 2278 2154 2282
rect 2150 2258 2154 2262
rect 2166 2198 2170 2202
rect 2150 2168 2154 2172
rect 2142 2068 2146 2072
rect 2150 1928 2154 1932
rect 2134 1858 2138 1862
rect 2126 1808 2130 1812
rect 2118 1708 2122 1712
rect 2142 1788 2146 1792
rect 2150 1748 2154 1752
rect 2134 1638 2138 1642
rect 2118 1508 2122 1512
rect 2086 958 2090 962
rect 2118 1128 2122 1132
rect 2118 1028 2122 1032
rect 2074 903 2078 907
rect 2081 903 2082 907
rect 2082 903 2085 907
rect 2086 838 2090 842
rect 2074 703 2078 707
rect 2081 703 2082 707
rect 2082 703 2085 707
rect 2062 558 2066 562
rect 2074 503 2078 507
rect 2081 503 2082 507
rect 2082 503 2085 507
rect 2102 888 2106 892
rect 2134 1398 2138 1402
rect 2182 2088 2186 2092
rect 2174 1848 2178 1852
rect 2166 1598 2170 1602
rect 2158 1488 2162 1492
rect 2166 1458 2170 1462
rect 2158 1428 2162 1432
rect 2142 1308 2146 1312
rect 2158 1258 2162 1262
rect 2134 1108 2138 1112
rect 2150 1168 2154 1172
rect 2134 858 2138 862
rect 2110 658 2114 662
rect 2102 648 2106 652
rect 2142 618 2146 622
rect 2074 303 2078 307
rect 2081 303 2082 307
rect 2082 303 2085 307
rect 2182 1758 2186 1762
rect 2198 2898 2202 2902
rect 2214 3218 2218 3222
rect 2198 2768 2202 2772
rect 2198 2598 2202 2602
rect 2238 3808 2242 3812
rect 2230 3688 2234 3692
rect 2238 3418 2242 3422
rect 2230 3038 2234 3042
rect 2222 2948 2226 2952
rect 2230 2948 2234 2952
rect 2222 2858 2226 2862
rect 2198 2498 2202 2502
rect 2198 2348 2202 2352
rect 2206 2288 2210 2292
rect 2206 2208 2210 2212
rect 2206 2018 2210 2022
rect 2198 1928 2202 1932
rect 2198 1848 2202 1852
rect 2190 1738 2194 1742
rect 2182 1718 2186 1722
rect 2190 1718 2194 1722
rect 2190 1698 2194 1702
rect 2206 1558 2210 1562
rect 2198 1488 2202 1492
rect 2190 1468 2194 1472
rect 2190 1458 2194 1462
rect 2198 1288 2202 1292
rect 2262 3958 2266 3962
rect 2294 4238 2298 4242
rect 2326 4178 2330 4182
rect 2294 3908 2298 3912
rect 2254 3688 2258 3692
rect 2246 3268 2250 3272
rect 2278 3688 2282 3692
rect 2374 4858 2378 4862
rect 2342 4328 2346 4332
rect 2374 4448 2378 4452
rect 2366 4428 2370 4432
rect 2390 4358 2394 4362
rect 2374 4288 2378 4292
rect 2350 4178 2354 4182
rect 2358 4068 2362 4072
rect 2342 4058 2346 4062
rect 2326 3918 2330 3922
rect 2318 3838 2322 3842
rect 2294 3608 2298 3612
rect 2286 3348 2290 3352
rect 2278 3288 2282 3292
rect 2286 3288 2290 3292
rect 2270 3218 2274 3222
rect 2294 3088 2298 3092
rect 2294 3048 2298 3052
rect 2262 2988 2266 2992
rect 2246 2748 2250 2752
rect 2246 2708 2250 2712
rect 2270 2668 2274 2672
rect 2246 2548 2250 2552
rect 2238 2538 2242 2542
rect 2230 2518 2234 2522
rect 2238 2468 2242 2472
rect 2230 2378 2234 2382
rect 2246 2358 2250 2362
rect 2238 2308 2242 2312
rect 2238 2278 2242 2282
rect 2262 2578 2266 2582
rect 2278 2628 2282 2632
rect 2278 2538 2282 2542
rect 2262 2348 2266 2352
rect 2254 2268 2258 2272
rect 2254 2068 2258 2072
rect 2246 2058 2250 2062
rect 2230 1888 2234 1892
rect 2246 1838 2250 1842
rect 2238 1768 2242 1772
rect 2246 1768 2250 1772
rect 2270 2278 2274 2282
rect 2270 2218 2274 2222
rect 2270 2108 2274 2112
rect 2294 2628 2298 2632
rect 2318 3808 2322 3812
rect 2350 3968 2354 3972
rect 2326 3798 2330 3802
rect 2318 3268 2322 3272
rect 2318 3168 2322 3172
rect 2334 3208 2338 3212
rect 2358 3668 2362 3672
rect 2350 3608 2354 3612
rect 2350 3538 2354 3542
rect 2318 2898 2322 2902
rect 2334 2858 2338 2862
rect 2310 2848 2314 2852
rect 2358 2988 2362 2992
rect 2358 2738 2362 2742
rect 2334 2608 2338 2612
rect 2318 2548 2322 2552
rect 2342 2508 2346 2512
rect 2318 2468 2322 2472
rect 2294 2328 2298 2332
rect 2310 2328 2314 2332
rect 2318 2188 2322 2192
rect 2262 1588 2266 1592
rect 2214 1218 2218 1222
rect 2246 1428 2250 1432
rect 2278 2008 2282 2012
rect 2286 1888 2290 1892
rect 2286 1618 2290 1622
rect 2278 1568 2282 1572
rect 2278 1528 2282 1532
rect 2286 1478 2290 1482
rect 2246 1408 2250 1412
rect 2270 1288 2274 1292
rect 2246 1148 2250 1152
rect 2222 1018 2226 1022
rect 2254 888 2258 892
rect 2270 848 2274 852
rect 2246 538 2250 542
rect 2310 2098 2314 2102
rect 2310 2078 2314 2082
rect 2310 1958 2314 1962
rect 2334 2388 2338 2392
rect 2334 2308 2338 2312
rect 2334 2228 2338 2232
rect 2350 2178 2354 2182
rect 2326 1938 2330 1942
rect 2302 1548 2306 1552
rect 2302 1418 2306 1422
rect 2310 1348 2314 1352
rect 2302 558 2306 562
rect 2334 1858 2338 1862
rect 2326 1628 2330 1632
rect 2326 1278 2330 1282
rect 2358 1848 2362 1852
rect 2358 1818 2362 1822
rect 2374 3838 2378 3842
rect 2390 4118 2394 4122
rect 2422 4478 2426 4482
rect 2586 4803 2590 4807
rect 2593 4803 2594 4807
rect 2594 4803 2597 4807
rect 2494 4528 2498 4532
rect 2502 4528 2506 4532
rect 2422 4138 2426 4142
rect 2422 4068 2426 4072
rect 2422 3868 2426 3872
rect 2438 4068 2442 4072
rect 2422 3858 2426 3862
rect 2406 3808 2410 3812
rect 2390 3768 2394 3772
rect 2430 3768 2434 3772
rect 2438 3738 2442 3742
rect 2398 3528 2402 3532
rect 2390 3478 2394 3482
rect 2390 3458 2394 3462
rect 2382 3368 2386 3372
rect 2382 3188 2386 3192
rect 2398 2928 2402 2932
rect 2398 2888 2402 2892
rect 2422 3518 2426 3522
rect 2422 3168 2426 3172
rect 2438 3538 2442 3542
rect 2494 3688 2498 3692
rect 2478 3668 2482 3672
rect 2478 3618 2482 3622
rect 2502 3568 2506 3572
rect 2478 3488 2482 3492
rect 2462 3338 2466 3342
rect 2486 3338 2490 3342
rect 2446 3188 2450 3192
rect 2414 3118 2418 3122
rect 2398 2568 2402 2572
rect 2406 2488 2410 2492
rect 2390 2458 2394 2462
rect 2398 2458 2402 2462
rect 2374 2408 2378 2412
rect 2374 2388 2378 2392
rect 2406 2398 2410 2402
rect 2438 3048 2442 3052
rect 2438 2968 2442 2972
rect 2430 2798 2434 2802
rect 2422 2518 2426 2522
rect 2422 2478 2426 2482
rect 2414 2358 2418 2362
rect 2414 2258 2418 2262
rect 2414 2168 2418 2172
rect 2398 2088 2402 2092
rect 2390 1878 2394 1882
rect 2374 1858 2378 1862
rect 2366 1668 2370 1672
rect 2390 1628 2394 1632
rect 2366 1588 2370 1592
rect 2414 1978 2418 1982
rect 2430 1898 2434 1902
rect 2430 1728 2434 1732
rect 2414 1718 2418 1722
rect 2462 3258 2466 3262
rect 2470 3118 2474 3122
rect 2454 2818 2458 2822
rect 2454 2668 2458 2672
rect 2486 3068 2490 3072
rect 2502 3348 2506 3352
rect 2662 4738 2666 4742
rect 2550 4688 2554 4692
rect 2534 4348 2538 4352
rect 2586 4603 2590 4607
rect 2593 4603 2594 4607
rect 2594 4603 2597 4607
rect 2566 4538 2570 4542
rect 2614 4408 2618 4412
rect 2586 4403 2590 4407
rect 2593 4403 2594 4407
rect 2594 4403 2597 4407
rect 2550 4348 2554 4352
rect 2586 4203 2590 4207
rect 2593 4203 2594 4207
rect 2594 4203 2597 4207
rect 2550 4058 2554 4062
rect 2518 3488 2522 3492
rect 2510 3258 2514 3262
rect 2510 3128 2514 3132
rect 2566 3668 2570 3672
rect 2558 3498 2562 3502
rect 2550 3348 2554 3352
rect 2558 3318 2562 3322
rect 2518 3108 2522 3112
rect 2534 3088 2538 3092
rect 2502 3078 2506 3082
rect 2526 3078 2530 3082
rect 2518 3068 2522 3072
rect 2502 3048 2506 3052
rect 2510 2898 2514 2902
rect 2510 2818 2514 2822
rect 2478 2808 2482 2812
rect 2470 2768 2474 2772
rect 2462 2508 2466 2512
rect 2462 2458 2466 2462
rect 2446 2198 2450 2202
rect 2446 1688 2450 1692
rect 2438 1678 2442 1682
rect 2446 1638 2450 1642
rect 2406 1418 2410 1422
rect 2398 1398 2402 1402
rect 2374 998 2378 1002
rect 2390 1338 2394 1342
rect 2374 928 2378 932
rect 2414 718 2418 722
rect 2422 648 2426 652
rect 2422 638 2426 642
rect 2398 588 2402 592
rect 2342 518 2346 522
rect 2398 518 2402 522
rect 2182 348 2186 352
rect 2166 268 2170 272
rect 2238 268 2242 272
rect 2206 258 2210 262
rect 2462 2238 2466 2242
rect 2502 2698 2506 2702
rect 2486 2678 2490 2682
rect 2494 2508 2498 2512
rect 2478 2438 2482 2442
rect 2510 2678 2514 2682
rect 2518 2598 2522 2602
rect 2502 2358 2506 2362
rect 2486 2218 2490 2222
rect 2494 2058 2498 2062
rect 2486 1968 2490 1972
rect 2510 2148 2514 2152
rect 2470 1938 2474 1942
rect 2494 1738 2498 1742
rect 2486 1728 2490 1732
rect 2462 1548 2466 1552
rect 2486 1578 2490 1582
rect 2478 1228 2482 1232
rect 2478 1008 2482 1012
rect 2470 888 2474 892
rect 2534 3038 2538 3042
rect 2534 2938 2538 2942
rect 2534 2878 2538 2882
rect 2542 2868 2546 2872
rect 2558 2868 2562 2872
rect 2558 2738 2562 2742
rect 2542 2638 2546 2642
rect 2558 2618 2562 2622
rect 2526 2358 2530 2362
rect 2518 2028 2522 2032
rect 2586 4003 2590 4007
rect 2593 4003 2594 4007
rect 2594 4003 2597 4007
rect 2606 3998 2610 4002
rect 2598 3918 2602 3922
rect 2586 3803 2590 3807
rect 2593 3803 2594 3807
rect 2594 3803 2597 3807
rect 2630 4258 2634 4262
rect 2622 3868 2626 3872
rect 2630 3778 2634 3782
rect 2586 3603 2590 3607
rect 2593 3603 2594 3607
rect 2594 3603 2597 3607
rect 2614 3588 2618 3592
rect 2574 3528 2578 3532
rect 2614 3518 2618 3522
rect 2586 3403 2590 3407
rect 2593 3403 2594 3407
rect 2594 3403 2597 3407
rect 2586 3203 2590 3207
rect 2593 3203 2594 3207
rect 2594 3203 2597 3207
rect 2614 3168 2618 3172
rect 2574 3088 2578 3092
rect 2542 2528 2546 2532
rect 2550 2458 2554 2462
rect 2534 2148 2538 2152
rect 2558 2228 2562 2232
rect 2542 2018 2546 2022
rect 2534 1908 2538 1912
rect 2542 1908 2546 1912
rect 2526 1658 2530 1662
rect 2510 1238 2514 1242
rect 2662 4218 2666 4222
rect 2654 4008 2658 4012
rect 2646 3798 2650 3802
rect 2646 3758 2650 3762
rect 2670 3648 2674 3652
rect 2630 3298 2634 3302
rect 2622 3118 2626 3122
rect 2614 3028 2618 3032
rect 2606 3008 2610 3012
rect 2586 3003 2590 3007
rect 2593 3003 2594 3007
rect 2594 3003 2597 3007
rect 2606 2918 2610 2922
rect 2586 2803 2590 2807
rect 2593 2803 2594 2807
rect 2594 2803 2597 2807
rect 3006 4738 3010 4742
rect 3098 4703 3102 4707
rect 3105 4703 3106 4707
rect 3106 4703 3109 4707
rect 2718 4658 2722 4662
rect 2710 4468 2714 4472
rect 2734 4448 2738 4452
rect 2686 3758 2690 3762
rect 2678 3478 2682 3482
rect 2678 3348 2682 3352
rect 2654 3278 2658 3282
rect 2654 3208 2658 3212
rect 2630 2938 2634 2942
rect 2622 2918 2626 2922
rect 2630 2848 2634 2852
rect 2622 2798 2626 2802
rect 2622 2638 2626 2642
rect 2606 2618 2610 2622
rect 2586 2603 2590 2607
rect 2593 2603 2594 2607
rect 2594 2603 2597 2607
rect 2614 2608 2618 2612
rect 2606 2488 2610 2492
rect 2586 2403 2590 2407
rect 2593 2403 2594 2407
rect 2594 2403 2597 2407
rect 2582 2368 2586 2372
rect 2574 2238 2578 2242
rect 2586 2203 2590 2207
rect 2593 2203 2594 2207
rect 2594 2203 2597 2207
rect 2582 2088 2586 2092
rect 2586 2003 2590 2007
rect 2593 2003 2594 2007
rect 2594 2003 2597 2007
rect 2558 1378 2562 1382
rect 2526 1138 2530 1142
rect 2518 1088 2522 1092
rect 2510 1028 2514 1032
rect 2542 1328 2546 1332
rect 2586 1803 2590 1807
rect 2593 1803 2594 1807
rect 2594 1803 2597 1807
rect 2574 1658 2578 1662
rect 2586 1603 2590 1607
rect 2593 1603 2594 1607
rect 2594 1603 2597 1607
rect 2586 1403 2590 1407
rect 2593 1403 2594 1407
rect 2594 1403 2597 1407
rect 2574 1388 2578 1392
rect 2582 1278 2586 1282
rect 2574 1268 2578 1272
rect 2586 1203 2590 1207
rect 2593 1203 2594 1207
rect 2594 1203 2597 1207
rect 2646 2958 2650 2962
rect 2646 2928 2650 2932
rect 2726 3898 2730 3902
rect 2702 3848 2706 3852
rect 2662 3138 2666 3142
rect 2686 3048 2690 3052
rect 2662 2998 2666 3002
rect 2662 2978 2666 2982
rect 2662 2938 2666 2942
rect 2662 2868 2666 2872
rect 2654 2718 2658 2722
rect 2702 2708 2706 2712
rect 2702 2688 2706 2692
rect 2694 2648 2698 2652
rect 2702 2648 2706 2652
rect 2638 2538 2642 2542
rect 2638 2528 2642 2532
rect 2646 2518 2650 2522
rect 2638 2498 2642 2502
rect 2630 2488 2634 2492
rect 2654 2468 2658 2472
rect 2630 2348 2634 2352
rect 2670 2348 2674 2352
rect 2678 2328 2682 2332
rect 2630 2228 2634 2232
rect 2614 2008 2618 2012
rect 2614 1888 2618 1892
rect 2630 1928 2634 1932
rect 2646 1878 2650 1882
rect 2622 1868 2626 1872
rect 2670 2078 2674 2082
rect 2678 2078 2682 2082
rect 2590 1118 2594 1122
rect 2590 1078 2594 1082
rect 2606 1078 2610 1082
rect 2586 1003 2590 1007
rect 2593 1003 2594 1007
rect 2594 1003 2597 1007
rect 2622 1178 2626 1182
rect 2638 1258 2642 1262
rect 2654 1168 2658 1172
rect 2622 1058 2626 1062
rect 2654 1058 2658 1062
rect 2670 1668 2674 1672
rect 2606 978 2610 982
rect 2662 978 2666 982
rect 2558 968 2562 972
rect 2566 968 2570 972
rect 2654 948 2658 952
rect 2638 918 2642 922
rect 2586 803 2590 807
rect 2593 803 2594 807
rect 2594 803 2597 807
rect 2614 778 2618 782
rect 2526 748 2530 752
rect 2454 738 2458 742
rect 2630 678 2634 682
rect 2654 658 2658 662
rect 2586 603 2590 607
rect 2593 603 2594 607
rect 2594 603 2597 607
rect 2878 4428 2882 4432
rect 2766 4228 2770 4232
rect 2798 4338 2802 4342
rect 2830 4338 2834 4342
rect 2846 4318 2850 4322
rect 2806 4188 2810 4192
rect 2782 4098 2786 4102
rect 2774 4078 2778 4082
rect 2758 3918 2762 3922
rect 2750 3688 2754 3692
rect 2758 3378 2762 3382
rect 2766 3378 2770 3382
rect 2742 3288 2746 3292
rect 2750 3198 2754 3202
rect 2726 3018 2730 3022
rect 2734 3018 2738 3022
rect 2718 2718 2722 2722
rect 2710 2608 2714 2612
rect 2710 2598 2714 2602
rect 2702 2548 2706 2552
rect 2702 2468 2706 2472
rect 2702 2368 2706 2372
rect 2694 2358 2698 2362
rect 2694 2208 2698 2212
rect 2710 2128 2714 2132
rect 2702 1858 2706 1862
rect 2702 1828 2706 1832
rect 2702 1748 2706 1752
rect 2694 1488 2698 1492
rect 2678 1138 2682 1142
rect 2678 948 2682 952
rect 2702 1468 2706 1472
rect 2702 1168 2706 1172
rect 2726 2578 2730 2582
rect 2758 3038 2762 3042
rect 2742 2808 2746 2812
rect 2822 4148 2826 4152
rect 2830 4068 2834 4072
rect 2830 4058 2834 4062
rect 2846 4138 2850 4142
rect 2846 3998 2850 4002
rect 2846 3958 2850 3962
rect 2822 3918 2826 3922
rect 2862 3918 2866 3922
rect 3038 4658 3042 4662
rect 3030 4648 3034 4652
rect 2998 4538 3002 4542
rect 2990 4528 2994 4532
rect 2966 4278 2970 4282
rect 2894 4058 2898 4062
rect 2878 3958 2882 3962
rect 2886 3928 2890 3932
rect 2926 4218 2930 4222
rect 2902 3828 2906 3832
rect 2814 3468 2818 3472
rect 2814 3338 2818 3342
rect 2814 3218 2818 3222
rect 2798 2858 2802 2862
rect 2854 3548 2858 3552
rect 2822 2828 2826 2832
rect 2758 2578 2762 2582
rect 2742 2498 2746 2502
rect 2742 2488 2746 2492
rect 2750 2408 2754 2412
rect 2734 2368 2738 2372
rect 2726 2008 2730 2012
rect 2726 1838 2730 1842
rect 2830 2788 2834 2792
rect 2814 2628 2818 2632
rect 2822 2578 2826 2582
rect 2798 2428 2802 2432
rect 2814 2478 2818 2482
rect 2822 2458 2826 2462
rect 2822 2348 2826 2352
rect 2814 2198 2818 2202
rect 2886 3458 2890 3462
rect 2902 3348 2906 3352
rect 2894 3318 2898 3322
rect 2950 4158 2954 4162
rect 2950 3958 2954 3962
rect 2934 3768 2938 3772
rect 2942 3358 2946 3362
rect 2870 3248 2874 3252
rect 2862 3048 2866 3052
rect 2854 2718 2858 2722
rect 2846 2708 2850 2712
rect 2846 2668 2850 2672
rect 2886 2948 2890 2952
rect 2878 2908 2882 2912
rect 2870 2658 2874 2662
rect 2846 2568 2850 2572
rect 2846 2538 2850 2542
rect 2838 2428 2842 2432
rect 2790 2058 2794 2062
rect 2782 1918 2786 1922
rect 2758 1678 2762 1682
rect 2734 1568 2738 1572
rect 2782 1678 2786 1682
rect 2774 1598 2778 1602
rect 2758 1528 2762 1532
rect 2774 1498 2778 1502
rect 2726 1068 2730 1072
rect 2718 1058 2722 1062
rect 2734 1018 2738 1022
rect 2742 988 2746 992
rect 2694 728 2698 732
rect 2646 468 2650 472
rect 2438 278 2442 282
rect 2586 403 2590 407
rect 2593 403 2594 407
rect 2594 403 2597 407
rect 2670 368 2674 372
rect 2686 348 2690 352
rect 2518 148 2522 152
rect 2374 118 2378 122
rect 2074 103 2078 107
rect 2081 103 2082 107
rect 2082 103 2085 107
rect 2766 1198 2770 1202
rect 2766 788 2770 792
rect 2806 1888 2810 1892
rect 2838 1738 2842 1742
rect 2886 2478 2890 2482
rect 2934 3148 2938 3152
rect 2918 3108 2922 3112
rect 2902 2778 2906 2782
rect 2902 2668 2906 2672
rect 2894 2438 2898 2442
rect 2918 2888 2922 2892
rect 2998 4018 3002 4022
rect 2990 3968 2994 3972
rect 3030 4278 3034 4282
rect 2958 3528 2962 3532
rect 2918 2328 2922 2332
rect 2878 2268 2882 2272
rect 2854 1848 2858 1852
rect 2870 1788 2874 1792
rect 2854 1758 2858 1762
rect 2830 1648 2834 1652
rect 2862 1648 2866 1652
rect 2806 1468 2810 1472
rect 2782 1038 2786 1042
rect 2798 798 2802 802
rect 2798 768 2802 772
rect 2798 548 2802 552
rect 2846 1578 2850 1582
rect 2870 1618 2874 1622
rect 2854 1538 2858 1542
rect 2838 1378 2842 1382
rect 2830 1208 2834 1212
rect 2838 958 2842 962
rect 2586 203 2590 207
rect 2593 203 2594 207
rect 2594 203 2597 207
rect 2782 268 2786 272
rect 2830 448 2834 452
rect 2590 128 2594 132
rect 2726 128 2730 132
rect 2750 118 2754 122
rect 2862 1508 2866 1512
rect 2902 1918 2906 1922
rect 2894 1618 2898 1622
rect 2934 2508 2938 2512
rect 2998 3658 3002 3662
rect 3610 4803 3614 4807
rect 3617 4803 3618 4807
rect 3618 4803 3621 4807
rect 3294 4638 3298 4642
rect 3046 3948 3050 3952
rect 3038 3808 3042 3812
rect 3014 3538 3018 3542
rect 2966 3478 2970 3482
rect 2966 3388 2970 3392
rect 2966 3178 2970 3182
rect 2974 3178 2978 3182
rect 2966 3148 2970 3152
rect 2974 3138 2978 3142
rect 2974 2948 2978 2952
rect 2998 3148 3002 3152
rect 2990 3098 2994 3102
rect 2982 2838 2986 2842
rect 2950 2528 2954 2532
rect 2958 2378 2962 2382
rect 2966 2348 2970 2352
rect 2966 2298 2970 2302
rect 2950 2258 2954 2262
rect 2966 2228 2970 2232
rect 2958 2208 2962 2212
rect 2966 2208 2970 2212
rect 2966 2178 2970 2182
rect 2926 2128 2930 2132
rect 2894 1518 2898 1522
rect 2902 1518 2906 1522
rect 2862 1328 2866 1332
rect 2846 858 2850 862
rect 2878 1258 2882 1262
rect 2894 858 2898 862
rect 2926 1628 2930 1632
rect 2942 1708 2946 1712
rect 2942 1628 2946 1632
rect 2918 1408 2922 1412
rect 2910 758 2914 762
rect 2926 1328 2930 1332
rect 2950 1368 2954 1372
rect 2942 1248 2946 1252
rect 2934 1148 2938 1152
rect 2982 2548 2986 2552
rect 3046 3658 3050 3662
rect 3022 3268 3026 3272
rect 3262 4548 3266 4552
rect 3098 4503 3102 4507
rect 3105 4503 3106 4507
rect 3106 4503 3109 4507
rect 3098 4303 3102 4307
rect 3105 4303 3106 4307
rect 3106 4303 3109 4307
rect 3406 4648 3410 4652
rect 3494 4548 3498 4552
rect 3198 4438 3202 4442
rect 3150 4418 3154 4422
rect 3198 4408 3202 4412
rect 3174 4338 3178 4342
rect 3150 4318 3154 4322
rect 3142 4238 3146 4242
rect 3134 4208 3138 4212
rect 3126 4148 3130 4152
rect 3126 4128 3130 4132
rect 3098 4103 3102 4107
rect 3105 4103 3106 4107
rect 3106 4103 3109 4107
rect 3078 3908 3082 3912
rect 3098 3903 3102 3907
rect 3105 3903 3106 3907
rect 3106 3903 3109 3907
rect 3070 3818 3074 3822
rect 3086 3748 3090 3752
rect 3098 3703 3102 3707
rect 3105 3703 3106 3707
rect 3106 3703 3109 3707
rect 3086 3698 3090 3702
rect 3118 3668 3122 3672
rect 3134 3918 3138 3922
rect 3182 4068 3186 4072
rect 3150 3598 3154 3602
rect 3134 3588 3138 3592
rect 3182 3568 3186 3572
rect 3098 3503 3102 3507
rect 3105 3503 3106 3507
rect 3106 3503 3109 3507
rect 3102 3478 3106 3482
rect 3054 3298 3058 3302
rect 3062 3258 3066 3262
rect 3046 3118 3050 3122
rect 3006 3078 3010 3082
rect 3046 3068 3050 3072
rect 3030 2978 3034 2982
rect 3014 2848 3018 2852
rect 3098 3303 3102 3307
rect 3105 3303 3106 3307
rect 3106 3303 3109 3307
rect 3078 3048 3082 3052
rect 3046 2838 3050 2842
rect 3118 3188 3122 3192
rect 3098 3103 3102 3107
rect 3105 3103 3106 3107
rect 3106 3103 3109 3107
rect 3110 2928 3114 2932
rect 3098 2903 3102 2907
rect 3105 2903 3106 2907
rect 3106 2903 3109 2907
rect 3214 4288 3218 4292
rect 3550 4658 3554 4662
rect 3542 4528 3546 4532
rect 3526 4518 3530 4522
rect 3518 4468 3522 4472
rect 3366 4378 3370 4382
rect 3318 4338 3322 4342
rect 3326 4338 3330 4342
rect 3278 4258 3282 4262
rect 3238 4078 3242 4082
rect 3230 4058 3234 4062
rect 3214 3718 3218 3722
rect 3222 3718 3226 3722
rect 3214 3568 3218 3572
rect 3206 3548 3210 3552
rect 3150 3448 3154 3452
rect 3142 3318 3146 3322
rect 3142 3298 3146 3302
rect 3102 2858 3106 2862
rect 3062 2798 3066 2802
rect 3038 2768 3042 2772
rect 3054 2708 3058 2712
rect 3006 2518 3010 2522
rect 3006 2498 3010 2502
rect 3006 2458 3010 2462
rect 2998 2368 3002 2372
rect 2990 2328 2994 2332
rect 2990 2278 2994 2282
rect 2998 2178 3002 2182
rect 2982 2118 2986 2122
rect 2998 2108 3002 2112
rect 2982 1948 2986 1952
rect 3022 2468 3026 2472
rect 3022 2228 3026 2232
rect 3022 2168 3026 2172
rect 3014 2088 3018 2092
rect 3006 1928 3010 1932
rect 3006 1578 3010 1582
rect 2998 1388 3002 1392
rect 3070 2698 3074 2702
rect 3070 2688 3074 2692
rect 3062 2318 3066 2322
rect 3078 2678 3082 2682
rect 3110 2848 3114 2852
rect 3126 2788 3130 2792
rect 3118 2708 3122 2712
rect 3098 2703 3102 2707
rect 3105 2703 3106 2707
rect 3106 2703 3109 2707
rect 3118 2678 3122 2682
rect 3126 2618 3130 2622
rect 3086 2608 3090 2612
rect 3134 2578 3138 2582
rect 3062 2238 3066 2242
rect 3054 2148 3058 2152
rect 3038 2098 3042 2102
rect 3030 1748 3034 1752
rect 2990 1078 2994 1082
rect 2974 918 2978 922
rect 2950 878 2954 882
rect 2966 818 2970 822
rect 2926 648 2930 652
rect 2910 478 2914 482
rect 2966 578 2970 582
rect 3038 1528 3042 1532
rect 3054 2118 3058 2122
rect 3078 2138 3082 2142
rect 3118 2508 3122 2512
rect 3098 2503 3102 2507
rect 3105 2503 3106 2507
rect 3106 2503 3109 2507
rect 3142 2518 3146 2522
rect 3142 2478 3146 2482
rect 3118 2428 3122 2432
rect 3126 2428 3130 2432
rect 3134 2408 3138 2412
rect 3110 2368 3114 2372
rect 3098 2303 3102 2307
rect 3105 2303 3106 2307
rect 3106 2303 3109 2307
rect 3118 2268 3122 2272
rect 3110 2218 3114 2222
rect 3098 2103 3102 2107
rect 3105 2103 3106 2107
rect 3106 2103 3109 2107
rect 3126 2098 3130 2102
rect 3118 2038 3122 2042
rect 3086 2018 3090 2022
rect 3098 1903 3102 1907
rect 3105 1903 3106 1907
rect 3106 1903 3109 1907
rect 3078 1898 3082 1902
rect 3070 1718 3074 1722
rect 3062 1528 3066 1532
rect 3054 1498 3058 1502
rect 3126 1908 3130 1912
rect 3158 2838 3162 2842
rect 3150 2458 3154 2462
rect 3158 2388 3162 2392
rect 3150 2188 3154 2192
rect 3174 2728 3178 2732
rect 3198 3258 3202 3262
rect 3190 3068 3194 3072
rect 3190 2998 3194 3002
rect 3190 2458 3194 2462
rect 3182 2408 3186 2412
rect 3254 4058 3258 4062
rect 3254 3668 3258 3672
rect 3246 3328 3250 3332
rect 3206 2808 3210 2812
rect 3206 2698 3210 2702
rect 3230 2598 3234 2602
rect 3214 2568 3218 2572
rect 3214 2478 3218 2482
rect 3206 2398 3210 2402
rect 3294 4218 3298 4222
rect 3278 3978 3282 3982
rect 3270 3208 3274 3212
rect 3342 4008 3346 4012
rect 3430 4248 3434 4252
rect 3406 4138 3410 4142
rect 3390 3918 3394 3922
rect 3366 3868 3370 3872
rect 3342 3858 3346 3862
rect 3334 3828 3338 3832
rect 3302 3548 3306 3552
rect 3310 3548 3314 3552
rect 3294 3478 3298 3482
rect 3342 3628 3346 3632
rect 3326 3458 3330 3462
rect 3326 3228 3330 3232
rect 3326 3058 3330 3062
rect 3326 2978 3330 2982
rect 3334 2848 3338 2852
rect 3262 2698 3266 2702
rect 3262 2638 3266 2642
rect 3254 2548 3258 2552
rect 3310 2588 3314 2592
rect 3254 2358 3258 2362
rect 3238 2298 3242 2302
rect 3214 2218 3218 2222
rect 3166 2038 3170 2042
rect 3206 2038 3210 2042
rect 3174 2028 3178 2032
rect 3238 2118 3242 2122
rect 3206 1968 3210 1972
rect 3182 1928 3186 1932
rect 3150 1918 3154 1922
rect 3086 1718 3090 1722
rect 3098 1703 3102 1707
rect 3105 1703 3106 1707
rect 3106 1703 3109 1707
rect 3086 1678 3090 1682
rect 3094 1678 3098 1682
rect 3142 1738 3146 1742
rect 3134 1638 3138 1642
rect 3094 1608 3098 1612
rect 3098 1503 3102 1507
rect 3105 1503 3106 1507
rect 3106 1503 3109 1507
rect 3190 1858 3194 1862
rect 3158 1788 3162 1792
rect 3166 1648 3170 1652
rect 3150 1528 3154 1532
rect 3118 1488 3122 1492
rect 3078 1458 3082 1462
rect 3126 1448 3130 1452
rect 3102 1418 3106 1422
rect 3110 1418 3114 1422
rect 3086 1398 3090 1402
rect 3038 1278 3042 1282
rect 3078 1098 3082 1102
rect 3070 1048 3074 1052
rect 2998 528 3002 532
rect 2990 338 2994 342
rect 2870 258 2874 262
rect 2838 138 2842 142
rect 2374 68 2378 72
rect 2686 68 2690 72
rect 2286 58 2290 62
rect 2750 58 2754 62
rect 3014 588 3018 592
rect 3070 748 3074 752
rect 3102 1348 3106 1352
rect 3142 1468 3146 1472
rect 3190 1728 3194 1732
rect 3198 1648 3202 1652
rect 3182 1488 3186 1492
rect 3182 1468 3186 1472
rect 3166 1308 3170 1312
rect 3098 1303 3102 1307
rect 3105 1303 3106 1307
rect 3106 1303 3109 1307
rect 3134 1298 3138 1302
rect 3110 1238 3114 1242
rect 3126 1118 3130 1122
rect 3098 1103 3102 1107
rect 3105 1103 3106 1107
rect 3106 1103 3109 1107
rect 3182 1258 3186 1262
rect 3150 1108 3154 1112
rect 3098 903 3102 907
rect 3105 903 3106 907
rect 3106 903 3109 907
rect 3094 718 3098 722
rect 3098 703 3102 707
rect 3105 703 3106 707
rect 3106 703 3109 707
rect 3062 658 3066 662
rect 3098 503 3102 507
rect 3105 503 3106 507
rect 3106 503 3109 507
rect 3142 928 3146 932
rect 3134 768 3138 772
rect 3182 1168 3186 1172
rect 3174 1158 3178 1162
rect 3134 688 3138 692
rect 3174 848 3178 852
rect 3158 658 3162 662
rect 3214 1648 3218 1652
rect 3214 1538 3218 1542
rect 3222 1498 3226 1502
rect 3214 1488 3218 1492
rect 3246 2108 3250 2112
rect 3262 2058 3266 2062
rect 3238 1498 3242 1502
rect 3214 1228 3218 1232
rect 3214 798 3218 802
rect 3206 728 3210 732
rect 3198 668 3202 672
rect 3098 303 3102 307
rect 3105 303 3106 307
rect 3106 303 3109 307
rect 3098 103 3102 107
rect 3105 103 3106 107
rect 3106 103 3109 107
rect 2654 48 2658 52
rect 2822 48 2826 52
rect 3254 1318 3258 1322
rect 3246 1298 3250 1302
rect 3254 1258 3258 1262
rect 3238 888 3242 892
rect 3230 738 3234 742
rect 3302 2448 3306 2452
rect 3302 2388 3306 2392
rect 3310 2368 3314 2372
rect 3310 2348 3314 2352
rect 3302 2208 3306 2212
rect 3286 2198 3290 2202
rect 3286 2158 3290 2162
rect 3318 2308 3322 2312
rect 3334 2548 3338 2552
rect 3350 2748 3354 2752
rect 3350 2678 3354 2682
rect 3350 2558 3354 2562
rect 3382 3838 3386 3842
rect 3390 3688 3394 3692
rect 3382 3508 3386 3512
rect 3382 3398 3386 3402
rect 3406 3578 3410 3582
rect 3374 3158 3378 3162
rect 3382 2548 3386 2552
rect 3374 2518 3378 2522
rect 3342 2418 3346 2422
rect 3350 2418 3354 2422
rect 3286 2098 3290 2102
rect 3278 1658 3282 1662
rect 3302 1948 3306 1952
rect 3302 1688 3306 1692
rect 3286 1248 3290 1252
rect 3382 2508 3386 2512
rect 3430 4108 3434 4112
rect 3430 3878 3434 3882
rect 3454 3968 3458 3972
rect 3446 3668 3450 3672
rect 3470 4088 3474 4092
rect 3470 3998 3474 4002
rect 3486 4038 3490 4042
rect 3478 3858 3482 3862
rect 3454 3638 3458 3642
rect 3454 3278 3458 3282
rect 3478 3588 3482 3592
rect 3470 3488 3474 3492
rect 3478 3488 3482 3492
rect 3446 3208 3450 3212
rect 3534 4478 3538 4482
rect 3534 3958 3538 3962
rect 3566 4128 3570 4132
rect 3610 4603 3614 4607
rect 3617 4603 3618 4607
rect 3618 4603 3621 4607
rect 3558 4108 3562 4112
rect 3518 3758 3522 3762
rect 3526 3728 3530 3732
rect 3542 3638 3546 3642
rect 3542 3598 3546 3602
rect 3494 3348 3498 3352
rect 3494 3328 3498 3332
rect 3518 3258 3522 3262
rect 3470 3168 3474 3172
rect 3430 3138 3434 3142
rect 3446 3138 3450 3142
rect 3462 3138 3466 3142
rect 3462 3128 3466 3132
rect 3430 3108 3434 3112
rect 3438 3058 3442 3062
rect 3430 2488 3434 2492
rect 3406 2438 3410 2442
rect 3414 2438 3418 2442
rect 3422 2428 3426 2432
rect 3454 2728 3458 2732
rect 3462 2528 3466 2532
rect 3462 2508 3466 2512
rect 3526 3068 3530 3072
rect 3502 2988 3506 2992
rect 3470 2448 3474 2452
rect 3478 2428 3482 2432
rect 3446 2418 3450 2422
rect 3438 2388 3442 2392
rect 3382 2358 3386 2362
rect 3422 2348 3426 2352
rect 3358 2238 3362 2242
rect 3350 2138 3354 2142
rect 3446 2308 3450 2312
rect 3422 2228 3426 2232
rect 3414 2218 3418 2222
rect 3422 2138 3426 2142
rect 3414 2068 3418 2072
rect 3326 2048 3330 2052
rect 3430 2068 3434 2072
rect 3358 2008 3362 2012
rect 3342 1998 3346 2002
rect 3350 1998 3354 2002
rect 3430 1998 3434 2002
rect 3414 1978 3418 1982
rect 3358 1958 3362 1962
rect 3382 1948 3386 1952
rect 3342 1638 3346 1642
rect 3318 1618 3322 1622
rect 3334 1608 3338 1612
rect 3326 1338 3330 1342
rect 3310 1298 3314 1302
rect 3294 1208 3298 1212
rect 3302 1188 3306 1192
rect 3294 1158 3298 1162
rect 3294 958 3298 962
rect 3294 908 3298 912
rect 3278 868 3282 872
rect 3270 848 3274 852
rect 3262 758 3266 762
rect 3342 1528 3346 1532
rect 3350 1528 3354 1532
rect 3358 1358 3362 1362
rect 3342 1188 3346 1192
rect 3342 1038 3346 1042
rect 3430 1948 3434 1952
rect 3430 1928 3434 1932
rect 3406 1848 3410 1852
rect 3382 1808 3386 1812
rect 3382 1778 3386 1782
rect 3406 1758 3410 1762
rect 3382 1668 3386 1672
rect 3414 1688 3418 1692
rect 3374 1238 3378 1242
rect 3374 1198 3378 1202
rect 3382 1168 3386 1172
rect 3366 1158 3370 1162
rect 3366 1058 3370 1062
rect 3374 948 3378 952
rect 3350 868 3354 872
rect 3350 858 3354 862
rect 3382 858 3386 862
rect 3358 738 3362 742
rect 3302 488 3306 492
rect 3254 338 3258 342
rect 3478 2298 3482 2302
rect 3462 2218 3466 2222
rect 3478 2128 3482 2132
rect 3454 2118 3458 2122
rect 3518 3008 3522 3012
rect 3526 2858 3530 2862
rect 3502 2388 3506 2392
rect 3494 2368 3498 2372
rect 3566 3988 3570 3992
rect 3566 3848 3570 3852
rect 3558 3798 3562 3802
rect 3550 2988 3554 2992
rect 3610 4403 3614 4407
rect 3617 4403 3618 4407
rect 3618 4403 3621 4407
rect 3598 4228 3602 4232
rect 3610 4203 3614 4207
rect 3617 4203 3618 4207
rect 3618 4203 3621 4207
rect 3630 4188 3634 4192
rect 3582 3728 3586 3732
rect 3590 3608 3594 3612
rect 3582 3528 3586 3532
rect 3574 3418 3578 3422
rect 3590 3198 3594 3202
rect 3574 3128 3578 3132
rect 3582 2898 3586 2902
rect 3574 2878 3578 2882
rect 3566 2828 3570 2832
rect 3558 2818 3562 2822
rect 3534 2748 3538 2752
rect 3518 2528 3522 2532
rect 3526 2468 3530 2472
rect 3526 2338 3530 2342
rect 3518 2318 3522 2322
rect 3518 2308 3522 2312
rect 3510 2198 3514 2202
rect 3454 2068 3458 2072
rect 3534 2138 3538 2142
rect 3510 2068 3514 2072
rect 3470 2028 3474 2032
rect 3446 1818 3450 1822
rect 3478 1878 3482 1882
rect 3486 1868 3490 1872
rect 3470 1848 3474 1852
rect 3446 1548 3450 1552
rect 3430 1408 3434 1412
rect 3414 1378 3418 1382
rect 3446 1438 3450 1442
rect 3470 1588 3474 1592
rect 3454 1398 3458 1402
rect 3438 1068 3442 1072
rect 3414 958 3418 962
rect 3430 888 3434 892
rect 3422 528 3426 532
rect 3438 838 3442 842
rect 3502 1728 3506 1732
rect 3558 2348 3562 2352
rect 3610 4003 3614 4007
rect 3617 4003 3618 4007
rect 3618 4003 3621 4007
rect 3614 3988 3618 3992
rect 3630 3938 3634 3942
rect 3614 3818 3618 3822
rect 3610 3803 3614 3807
rect 3617 3803 3618 3807
rect 3618 3803 3621 3807
rect 3610 3603 3614 3607
rect 3617 3603 3618 3607
rect 3618 3603 3621 3607
rect 3610 3403 3614 3407
rect 3617 3403 3618 3407
rect 3618 3403 3621 3407
rect 3622 3328 3626 3332
rect 3610 3203 3614 3207
rect 3617 3203 3618 3207
rect 3618 3203 3621 3207
rect 3610 3003 3614 3007
rect 3617 3003 3618 3007
rect 3618 3003 3621 3007
rect 3614 2968 3618 2972
rect 3606 2948 3610 2952
rect 3670 4018 3674 4022
rect 3662 3968 3666 3972
rect 3638 3688 3642 3692
rect 3710 4158 3714 4162
rect 3670 3788 3674 3792
rect 3662 3558 3666 3562
rect 3646 3278 3650 3282
rect 3638 2938 3642 2942
rect 3598 2838 3602 2842
rect 3610 2803 3614 2807
rect 3617 2803 3618 2807
rect 3618 2803 3621 2807
rect 3614 2788 3618 2792
rect 3598 2758 3602 2762
rect 3582 2658 3586 2662
rect 3574 2548 3578 2552
rect 3566 2338 3570 2342
rect 3566 2288 3570 2292
rect 3694 3858 3698 3862
rect 3726 4148 3730 4152
rect 3766 4338 3770 4342
rect 3790 4278 3794 4282
rect 3790 4228 3794 4232
rect 3822 4438 3826 4442
rect 3742 4038 3746 4042
rect 3750 3978 3754 3982
rect 3718 3888 3722 3892
rect 3702 3678 3706 3682
rect 3678 3268 3682 3272
rect 3662 2938 3666 2942
rect 3654 2908 3658 2912
rect 3630 2618 3634 2622
rect 3610 2603 3614 2607
rect 3617 2603 3618 2607
rect 3618 2603 3621 2607
rect 3622 2548 3626 2552
rect 3614 2538 3618 2542
rect 3622 2478 3626 2482
rect 3614 2418 3618 2422
rect 3610 2403 3614 2407
rect 3617 2403 3618 2407
rect 3618 2403 3621 2407
rect 3622 2368 3626 2372
rect 3614 2278 3618 2282
rect 3630 2258 3634 2262
rect 3574 2228 3578 2232
rect 3598 2228 3602 2232
rect 3558 2188 3562 2192
rect 3550 2178 3554 2182
rect 3566 2078 3570 2082
rect 3610 2203 3614 2207
rect 3617 2203 3618 2207
rect 3618 2203 3621 2207
rect 3630 2198 3634 2202
rect 3598 2128 3602 2132
rect 3582 2058 3586 2062
rect 3574 2008 3578 2012
rect 3558 1948 3562 1952
rect 3574 1898 3578 1902
rect 3610 2003 3614 2007
rect 3617 2003 3618 2007
rect 3618 2003 3621 2007
rect 3606 1908 3610 1912
rect 3630 1878 3634 1882
rect 3582 1808 3586 1812
rect 3550 1768 3554 1772
rect 3610 1803 3614 1807
rect 3617 1803 3618 1807
rect 3618 1803 3621 1807
rect 3518 1708 3522 1712
rect 3502 1658 3506 1662
rect 3486 1458 3490 1462
rect 3486 1078 3490 1082
rect 3566 1638 3570 1642
rect 3518 1258 3522 1262
rect 3526 1248 3530 1252
rect 3518 1128 3522 1132
rect 3518 798 3522 802
rect 3518 628 3522 632
rect 3454 538 3458 542
rect 3598 1748 3602 1752
rect 3598 1618 3602 1622
rect 3610 1603 3614 1607
rect 3617 1603 3618 1607
rect 3618 1603 3621 1607
rect 3598 1598 3602 1602
rect 3622 1568 3626 1572
rect 3630 1558 3634 1562
rect 3582 1538 3586 1542
rect 3558 1218 3562 1222
rect 3574 1448 3578 1452
rect 3534 558 3538 562
rect 3558 558 3562 562
rect 3486 148 3490 152
rect 3406 138 3410 142
rect 3590 1528 3594 1532
rect 3610 1403 3614 1407
rect 3617 1403 3618 1407
rect 3618 1403 3621 1407
rect 3622 1328 3626 1332
rect 3622 1268 3626 1272
rect 3610 1203 3614 1207
rect 3617 1203 3618 1207
rect 3618 1203 3621 1207
rect 3654 2148 3658 2152
rect 3646 1828 3650 1832
rect 3734 3778 3738 3782
rect 3718 3688 3722 3692
rect 3734 3668 3738 3672
rect 3742 3448 3746 3452
rect 3718 3248 3722 3252
rect 3742 3318 3746 3322
rect 3766 3628 3770 3632
rect 3790 4048 3794 4052
rect 3806 4028 3810 4032
rect 3790 3498 3794 3502
rect 3782 3438 3786 3442
rect 3758 3248 3762 3252
rect 3750 3138 3754 3142
rect 3726 3008 3730 3012
rect 3710 2958 3714 2962
rect 3718 2948 3722 2952
rect 3718 2838 3722 2842
rect 3702 2758 3706 2762
rect 3750 2948 3754 2952
rect 3750 2848 3754 2852
rect 3766 2848 3770 2852
rect 3814 3528 3818 3532
rect 3814 3508 3818 3512
rect 3878 4268 3882 4272
rect 3830 3638 3834 3642
rect 3798 3378 3802 3382
rect 3830 3088 3834 3092
rect 3806 3078 3810 3082
rect 3838 3068 3842 3072
rect 3822 3048 3826 3052
rect 3838 3038 3842 3042
rect 3790 2898 3794 2902
rect 3782 2888 3786 2892
rect 3790 2858 3794 2862
rect 3774 2828 3778 2832
rect 3750 2808 3754 2812
rect 3766 2788 3770 2792
rect 3782 2788 3786 2792
rect 3742 2728 3746 2732
rect 3686 2718 3690 2722
rect 3726 2708 3730 2712
rect 3694 2698 3698 2702
rect 3686 2678 3690 2682
rect 3670 2238 3674 2242
rect 3662 2068 3666 2072
rect 3702 2478 3706 2482
rect 3718 2468 3722 2472
rect 3702 2448 3706 2452
rect 3694 2338 3698 2342
rect 3646 1578 3650 1582
rect 3638 1188 3642 1192
rect 3610 1003 3614 1007
rect 3617 1003 3618 1007
rect 3618 1003 3621 1007
rect 3630 978 3634 982
rect 3610 803 3614 807
rect 3617 803 3618 807
rect 3618 803 3621 807
rect 3610 603 3614 607
rect 3617 603 3618 607
rect 3618 603 3621 607
rect 3678 1778 3682 1782
rect 3670 1578 3674 1582
rect 3694 2158 3698 2162
rect 3694 1858 3698 1862
rect 3686 1758 3690 1762
rect 3686 1668 3690 1672
rect 3678 1178 3682 1182
rect 3670 1098 3674 1102
rect 3574 548 3578 552
rect 3646 518 3650 522
rect 3610 403 3614 407
rect 3617 403 3618 407
rect 3618 403 3621 407
rect 3646 368 3650 372
rect 3718 2248 3722 2252
rect 3710 2218 3714 2222
rect 3734 2238 3738 2242
rect 3766 2428 3770 2432
rect 3750 2368 3754 2372
rect 3758 2298 3762 2302
rect 3742 2208 3746 2212
rect 3750 2188 3754 2192
rect 3758 2188 3762 2192
rect 3742 2178 3746 2182
rect 3734 2118 3738 2122
rect 3726 1988 3730 1992
rect 3710 1608 3714 1612
rect 3774 2268 3778 2272
rect 3806 2798 3810 2802
rect 3822 2768 3826 2772
rect 3806 2718 3810 2722
rect 3806 2528 3810 2532
rect 3806 2468 3810 2472
rect 3790 2458 3794 2462
rect 3798 2378 3802 2382
rect 3806 2368 3810 2372
rect 3814 2348 3818 2352
rect 3782 2258 3786 2262
rect 3758 2008 3762 2012
rect 3790 2018 3794 2022
rect 3774 1808 3778 1812
rect 3758 1798 3762 1802
rect 3742 1768 3746 1772
rect 3766 1718 3770 1722
rect 3774 1638 3778 1642
rect 3758 1598 3762 1602
rect 3718 1448 3722 1452
rect 3742 1388 3746 1392
rect 3758 1348 3762 1352
rect 3726 1238 3730 1242
rect 3750 1148 3754 1152
rect 3798 1778 3802 1782
rect 3790 1688 3794 1692
rect 3798 1568 3802 1572
rect 3798 1358 3802 1362
rect 3878 4018 3882 4022
rect 3918 4458 3922 4462
rect 3942 4348 3946 4352
rect 3902 4238 3906 4242
rect 3942 4248 3946 4252
rect 3918 3968 3922 3972
rect 3942 4058 3946 4062
rect 3958 4058 3962 4062
rect 3878 3648 3882 3652
rect 3902 3758 3906 3762
rect 3894 3468 3898 3472
rect 3862 3378 3866 3382
rect 3894 3238 3898 3242
rect 3910 3508 3914 3512
rect 3910 3328 3914 3332
rect 3902 3128 3906 3132
rect 3862 2928 3866 2932
rect 3838 2878 3842 2882
rect 3854 2878 3858 2882
rect 3846 2858 3850 2862
rect 3862 2758 3866 2762
rect 3846 2648 3850 2652
rect 3830 2358 3834 2362
rect 3846 2358 3850 2362
rect 3830 2338 3834 2342
rect 3814 1878 3818 1882
rect 3830 1748 3834 1752
rect 3814 1738 3818 1742
rect 3822 1678 3826 1682
rect 3814 1438 3818 1442
rect 3862 2528 3866 2532
rect 3862 2458 3866 2462
rect 3934 3348 3938 3352
rect 3926 3328 3930 3332
rect 3910 3068 3914 3072
rect 3878 2728 3882 2732
rect 3870 2338 3874 2342
rect 3854 2248 3858 2252
rect 3870 2248 3874 2252
rect 3854 2168 3858 2172
rect 3870 2218 3874 2222
rect 3862 2098 3866 2102
rect 3854 1948 3858 1952
rect 3854 1698 3858 1702
rect 3838 1658 3842 1662
rect 3838 1548 3842 1552
rect 3814 1308 3818 1312
rect 3806 1158 3810 1162
rect 3798 1148 3802 1152
rect 3830 1258 3834 1262
rect 3806 908 3810 912
rect 3782 848 3786 852
rect 3838 1238 3842 1242
rect 3830 1148 3834 1152
rect 3830 788 3834 792
rect 3726 748 3730 752
rect 3718 738 3722 742
rect 3862 1528 3866 1532
rect 3958 3898 3962 3902
rect 3950 3578 3954 3582
rect 3950 3448 3954 3452
rect 3926 2768 3930 2772
rect 3926 2738 3930 2742
rect 3918 2678 3922 2682
rect 3910 2558 3914 2562
rect 3910 2488 3914 2492
rect 3902 2368 3906 2372
rect 3902 2078 3906 2082
rect 3886 2048 3890 2052
rect 3894 2048 3898 2052
rect 3878 1568 3882 1572
rect 3878 1458 3882 1462
rect 3870 1298 3874 1302
rect 3878 1248 3882 1252
rect 3910 2038 3914 2042
rect 3894 1938 3898 1942
rect 3902 1918 3906 1922
rect 3894 1538 3898 1542
rect 3910 1498 3914 1502
rect 3926 2638 3930 2642
rect 3934 2508 3938 2512
rect 3926 1958 3930 1962
rect 3990 4308 3994 4312
rect 4022 4328 4026 4332
rect 3990 4138 3994 4142
rect 3990 4118 3994 4122
rect 3990 4088 3994 4092
rect 4006 4088 4010 4092
rect 3990 3658 3994 3662
rect 3998 3598 4002 3602
rect 3982 3448 3986 3452
rect 3966 3338 3970 3342
rect 3966 3298 3970 3302
rect 3966 3268 3970 3272
rect 3966 3248 3970 3252
rect 3966 2908 3970 2912
rect 3990 3278 3994 3282
rect 3990 3168 3994 3172
rect 4022 4248 4026 4252
rect 4022 3598 4026 3602
rect 4022 3158 4026 3162
rect 4014 3148 4018 3152
rect 4014 3108 4018 3112
rect 4014 3078 4018 3082
rect 3990 2988 3994 2992
rect 3974 2728 3978 2732
rect 3958 2568 3962 2572
rect 3950 2478 3954 2482
rect 3950 2458 3954 2462
rect 3942 2088 3946 2092
rect 3942 2058 3946 2062
rect 3942 2048 3946 2052
rect 3934 1758 3938 1762
rect 3846 1158 3850 1162
rect 3862 1058 3866 1062
rect 3846 828 3850 832
rect 3774 718 3778 722
rect 3686 368 3690 372
rect 3610 203 3614 207
rect 3617 203 3618 207
rect 3618 203 3621 207
rect 3870 348 3874 352
rect 3918 948 3922 952
rect 3934 1418 3938 1422
rect 3966 2498 3970 2502
rect 3974 2438 3978 2442
rect 3982 2428 3986 2432
rect 3990 2418 3994 2422
rect 3974 2248 3978 2252
rect 3982 2178 3986 2182
rect 3990 2178 3994 2182
rect 4022 2998 4026 3002
rect 4014 2688 4018 2692
rect 4014 2668 4018 2672
rect 4006 2208 4010 2212
rect 3998 2128 4002 2132
rect 4038 4278 4042 4282
rect 4046 4258 4050 4262
rect 4038 4248 4042 4252
rect 4114 4703 4118 4707
rect 4121 4703 4122 4707
rect 4122 4703 4125 4707
rect 4086 4458 4090 4462
rect 4086 4348 4090 4352
rect 4062 4268 4066 4272
rect 4046 4048 4050 4052
rect 4038 3948 4042 3952
rect 4070 4128 4074 4132
rect 4062 3868 4066 3872
rect 4046 3728 4050 3732
rect 4038 3298 4042 3302
rect 4038 3278 4042 3282
rect 4038 3128 4042 3132
rect 4062 3578 4066 3582
rect 4038 2918 4042 2922
rect 4114 4503 4118 4507
rect 4121 4503 4122 4507
rect 4122 4503 4125 4507
rect 4150 4428 4154 4432
rect 4114 4303 4118 4307
rect 4121 4303 4122 4307
rect 4122 4303 4125 4307
rect 4070 3108 4074 3112
rect 4054 2718 4058 2722
rect 4046 2698 4050 2702
rect 4038 2218 4042 2222
rect 4038 2158 4042 2162
rect 4030 2038 4034 2042
rect 4022 2018 4026 2022
rect 4014 1978 4018 1982
rect 4022 1968 4026 1972
rect 4022 1948 4026 1952
rect 3974 1858 3978 1862
rect 3966 1718 3970 1722
rect 3958 1518 3962 1522
rect 3950 1278 3954 1282
rect 3934 1038 3938 1042
rect 3926 888 3930 892
rect 3934 838 3938 842
rect 4006 1878 4010 1882
rect 3990 1758 3994 1762
rect 3998 1708 4002 1712
rect 3998 1688 4002 1692
rect 3990 1678 3994 1682
rect 3982 1308 3986 1312
rect 3998 1288 4002 1292
rect 3990 948 3994 952
rect 4030 1908 4034 1912
rect 4038 1838 4042 1842
rect 4038 1598 4042 1602
rect 4062 2698 4066 2702
rect 4054 2628 4058 2632
rect 4078 2968 4082 2972
rect 4114 4103 4118 4107
rect 4121 4103 4122 4107
rect 4122 4103 4125 4107
rect 4094 4078 4098 4082
rect 4094 4048 4098 4052
rect 4114 3903 4118 3907
rect 4121 3903 4122 3907
rect 4122 3903 4125 3907
rect 4158 4278 4162 4282
rect 4206 4648 4210 4652
rect 4174 4038 4178 4042
rect 4150 3958 4154 3962
rect 4230 4058 4234 4062
rect 4222 3978 4226 3982
rect 4182 3888 4186 3892
rect 4114 3703 4118 3707
rect 4121 3703 4122 3707
rect 4122 3703 4125 3707
rect 4102 3638 4106 3642
rect 4118 3538 4122 3542
rect 4114 3503 4118 3507
rect 4121 3503 4122 3507
rect 4122 3503 4125 3507
rect 4114 3303 4118 3307
rect 4121 3303 4122 3307
rect 4122 3303 4125 3307
rect 4198 3858 4202 3862
rect 4190 3688 4194 3692
rect 4102 3108 4106 3112
rect 4078 2728 4082 2732
rect 4078 2588 4082 2592
rect 4070 2328 4074 2332
rect 4054 2118 4058 2122
rect 4054 2068 4058 2072
rect 4062 1928 4066 1932
rect 4114 3103 4118 3107
rect 4121 3103 4122 3107
rect 4122 3103 4125 3107
rect 4150 3328 4154 3332
rect 4142 3058 4146 3062
rect 4126 2938 4130 2942
rect 4114 2903 4118 2907
rect 4121 2903 4122 2907
rect 4122 2903 4125 2907
rect 4134 2768 4138 2772
rect 4114 2703 4118 2707
rect 4121 2703 4122 2707
rect 4122 2703 4125 2707
rect 4126 2518 4130 2522
rect 4102 2508 4106 2512
rect 4114 2503 4118 2507
rect 4121 2503 4122 2507
rect 4122 2503 4125 2507
rect 4114 2303 4118 2307
rect 4121 2303 4122 2307
rect 4122 2303 4125 2307
rect 4118 2268 4122 2272
rect 4086 2218 4090 2222
rect 4094 2118 4098 2122
rect 4094 1978 4098 1982
rect 4086 1958 4090 1962
rect 4086 1898 4090 1902
rect 4078 1788 4082 1792
rect 4078 1768 4082 1772
rect 4078 1688 4082 1692
rect 4078 1638 4082 1642
rect 4062 1568 4066 1572
rect 4078 1578 4082 1582
rect 4070 1558 4074 1562
rect 4062 1508 4066 1512
rect 4046 1368 4050 1372
rect 4054 1328 4058 1332
rect 4014 958 4018 962
rect 3998 588 4002 592
rect 3958 348 3962 352
rect 3670 78 3674 82
rect 3950 68 3954 72
rect 3414 58 3418 62
rect 3510 58 3514 62
rect 4030 558 4034 562
rect 4030 458 4034 462
rect 4054 1168 4058 1172
rect 4078 1108 4082 1112
rect 4114 2103 4118 2107
rect 4121 2103 4122 2107
rect 4122 2103 4125 2107
rect 4134 2058 4138 2062
rect 4118 2028 4122 2032
rect 4110 1998 4114 2002
rect 4114 1903 4118 1907
rect 4121 1903 4122 1907
rect 4122 1903 4125 1907
rect 4118 1868 4122 1872
rect 4114 1703 4118 1707
rect 4121 1703 4122 1707
rect 4122 1703 4125 1707
rect 4102 1578 4106 1582
rect 4114 1503 4118 1507
rect 4121 1503 4122 1507
rect 4122 1503 4125 1507
rect 4126 1478 4130 1482
rect 4158 3038 4162 3042
rect 4150 2648 4154 2652
rect 4222 3958 4226 3962
rect 4230 3928 4234 3932
rect 4222 3848 4226 3852
rect 4206 3298 4210 3302
rect 4182 2928 4186 2932
rect 4166 2888 4170 2892
rect 4182 2888 4186 2892
rect 4174 2858 4178 2862
rect 4190 2858 4194 2862
rect 4182 2848 4186 2852
rect 4190 2848 4194 2852
rect 4158 2538 4162 2542
rect 4206 3018 4210 3022
rect 4206 2678 4210 2682
rect 4222 3268 4226 3272
rect 4262 4258 4266 4262
rect 4310 4528 4314 4532
rect 4398 4418 4402 4422
rect 4278 4338 4282 4342
rect 4254 3878 4258 3882
rect 4262 3828 4266 3832
rect 4238 3348 4242 3352
rect 4238 3218 4242 3222
rect 4246 3188 4250 3192
rect 4230 2878 4234 2882
rect 4230 2738 4234 2742
rect 4214 2528 4218 2532
rect 4174 2468 4178 2472
rect 4190 2448 4194 2452
rect 4174 2348 4178 2352
rect 4182 2258 4186 2262
rect 4166 2098 4170 2102
rect 4174 2048 4178 2052
rect 4150 2028 4154 2032
rect 4166 1938 4170 1942
rect 4246 2338 4250 2342
rect 4222 2228 4226 2232
rect 4206 2188 4210 2192
rect 4214 2128 4218 2132
rect 4190 1938 4194 1942
rect 4166 1848 4170 1852
rect 4174 1818 4178 1822
rect 4158 1648 4162 1652
rect 4166 1528 4170 1532
rect 4134 1368 4138 1372
rect 4114 1303 4118 1307
rect 4121 1303 4122 1307
rect 4122 1303 4125 1307
rect 4118 1128 4122 1132
rect 4114 1103 4118 1107
rect 4121 1103 4122 1107
rect 4122 1103 4125 1107
rect 4182 1498 4186 1502
rect 4114 903 4118 907
rect 4121 903 4122 907
rect 4122 903 4125 907
rect 4086 748 4090 752
rect 4062 678 4066 682
rect 4054 658 4058 662
rect 4054 538 4058 542
rect 4114 703 4118 707
rect 4121 703 4122 707
rect 4122 703 4125 707
rect 4126 518 4130 522
rect 4114 503 4118 507
rect 4121 503 4122 507
rect 4122 503 4125 507
rect 4142 348 4146 352
rect 4114 303 4118 307
rect 4121 303 4122 307
rect 4122 303 4125 307
rect 4198 1848 4202 1852
rect 4318 4068 4322 4072
rect 4294 3968 4298 3972
rect 4262 3308 4266 3312
rect 4270 3148 4274 3152
rect 4262 3068 4266 3072
rect 4318 3848 4322 3852
rect 4318 3738 4322 3742
rect 4310 3568 4314 3572
rect 4302 3508 4306 3512
rect 4286 3008 4290 3012
rect 4278 2558 4282 2562
rect 4254 2228 4258 2232
rect 4238 1978 4242 1982
rect 4230 1968 4234 1972
rect 4222 1738 4226 1742
rect 4230 1688 4234 1692
rect 4182 968 4186 972
rect 4206 1588 4210 1592
rect 4254 1758 4258 1762
rect 4254 1468 4258 1472
rect 4230 1138 4234 1142
rect 4206 468 4210 472
rect 4174 268 4178 272
rect 4198 348 4202 352
rect 4038 138 4042 142
rect 4114 103 4118 107
rect 4121 103 4122 107
rect 4122 103 4125 107
rect 4254 838 4258 842
rect 4318 3118 4322 3122
rect 4286 2258 4290 2262
rect 4294 2068 4298 2072
rect 4278 1888 4282 1892
rect 4294 1888 4298 1892
rect 4278 1548 4282 1552
rect 4294 1758 4298 1762
rect 4302 1748 4306 1752
rect 4286 1348 4290 1352
rect 4398 3958 4402 3962
rect 4358 3838 4362 3842
rect 4358 3648 4362 3652
rect 4342 3468 4346 3472
rect 4342 3058 4346 3062
rect 4334 2938 4338 2942
rect 4334 2808 4338 2812
rect 4350 2848 4354 2852
rect 4350 2808 4354 2812
rect 4366 3468 4370 3472
rect 4478 4538 4482 4542
rect 4430 4528 4434 4532
rect 4558 4578 4562 4582
rect 4518 4538 4522 4542
rect 4494 4518 4498 4522
rect 4446 4368 4450 4372
rect 4542 4408 4546 4412
rect 4446 3858 4450 3862
rect 4454 3608 4458 3612
rect 4398 3458 4402 3462
rect 4382 3258 4386 3262
rect 4390 3228 4394 3232
rect 4374 2828 4378 2832
rect 4366 2588 4370 2592
rect 4358 2478 4362 2482
rect 4350 2368 4354 2372
rect 4350 2348 4354 2352
rect 4358 2308 4362 2312
rect 4342 2148 4346 2152
rect 4342 2138 4346 2142
rect 4334 1938 4338 1942
rect 4350 1888 4354 1892
rect 4334 1648 4338 1652
rect 4318 1488 4322 1492
rect 4342 1598 4346 1602
rect 4350 1578 4354 1582
rect 4430 3528 4434 3532
rect 4494 3808 4498 3812
rect 4606 4458 4610 4462
rect 4558 4328 4562 4332
rect 4606 4268 4610 4272
rect 4542 4158 4546 4162
rect 4534 4148 4538 4152
rect 4550 4128 4554 4132
rect 4510 3718 4514 3722
rect 4470 3518 4474 3522
rect 4422 3298 4426 3302
rect 4438 3288 4442 3292
rect 4406 2858 4410 2862
rect 4390 2568 4394 2572
rect 4382 2448 4386 2452
rect 4382 2438 4386 2442
rect 4366 2168 4370 2172
rect 4390 2298 4394 2302
rect 4390 2228 4394 2232
rect 4382 2128 4386 2132
rect 4366 2118 4370 2122
rect 4374 1948 4378 1952
rect 4398 2198 4402 2202
rect 4382 1868 4386 1872
rect 4374 1818 4378 1822
rect 4374 1748 4378 1752
rect 4374 1658 4378 1662
rect 4358 1478 4362 1482
rect 4366 1468 4370 1472
rect 4430 2828 4434 2832
rect 4414 2248 4418 2252
rect 4414 2058 4418 2062
rect 4414 1958 4418 1962
rect 4406 1708 4410 1712
rect 4398 1548 4402 1552
rect 4390 1358 4394 1362
rect 4342 1258 4346 1262
rect 4342 1168 4346 1172
rect 4326 968 4330 972
rect 4326 828 4330 832
rect 4270 738 4274 742
rect 4310 758 4314 762
rect 4358 1178 4362 1182
rect 4358 1018 4362 1022
rect 4358 928 4362 932
rect 4310 468 4314 472
rect 4510 3358 4514 3362
rect 4598 4168 4602 4172
rect 4558 3868 4562 3872
rect 4550 3848 4554 3852
rect 4518 3328 4522 3332
rect 4550 3528 4554 3532
rect 4542 3278 4546 3282
rect 4534 3148 4538 3152
rect 4454 2978 4458 2982
rect 4462 2978 4466 2982
rect 4486 3038 4490 3042
rect 4470 2968 4474 2972
rect 4462 2958 4466 2962
rect 4462 2898 4466 2902
rect 4438 2738 4442 2742
rect 4462 2728 4466 2732
rect 4446 2718 4450 2722
rect 4430 2488 4434 2492
rect 4438 2468 4442 2472
rect 4446 2288 4450 2292
rect 4470 2538 4474 2542
rect 4494 2988 4498 2992
rect 4494 2528 4498 2532
rect 4478 2398 4482 2402
rect 4470 2338 4474 2342
rect 4470 2218 4474 2222
rect 4486 2178 4490 2182
rect 4470 2078 4474 2082
rect 4430 1958 4434 1962
rect 4486 2028 4490 2032
rect 4462 1888 4466 1892
rect 4454 1858 4458 1862
rect 4438 1748 4442 1752
rect 4446 1698 4450 1702
rect 4430 1478 4434 1482
rect 4422 1128 4426 1132
rect 4430 1028 4434 1032
rect 4470 1788 4474 1792
rect 4470 1668 4474 1672
rect 4470 1598 4474 1602
rect 4486 1218 4490 1222
rect 4486 938 4490 942
rect 4406 548 4410 552
rect 4382 468 4386 472
rect 4286 258 4290 262
rect 4366 258 4370 262
rect 4214 138 4218 142
rect 4230 138 4234 142
rect 4206 78 4210 82
rect 4398 78 4402 82
rect 4478 538 4482 542
rect 4526 3048 4530 3052
rect 4526 2838 4530 2842
rect 4526 2538 4530 2542
rect 4574 3858 4578 3862
rect 4574 3748 4578 3752
rect 4566 3368 4570 3372
rect 4550 2858 4554 2862
rect 4510 2068 4514 2072
rect 4502 1648 4506 1652
rect 4502 1488 4506 1492
rect 4542 2358 4546 2362
rect 4518 1338 4522 1342
rect 4574 3338 4578 3342
rect 4606 3868 4610 3872
rect 4590 3368 4594 3372
rect 4590 3358 4594 3362
rect 4590 3278 4594 3282
rect 4582 3038 4586 3042
rect 4590 2968 4594 2972
rect 4598 2958 4602 2962
rect 4574 2428 4578 2432
rect 4566 2228 4570 2232
rect 4550 2128 4554 2132
rect 4542 1848 4546 1852
rect 4550 1808 4554 1812
rect 4542 1668 4546 1672
rect 4550 1638 4554 1642
rect 4550 1348 4554 1352
rect 4526 1198 4530 1202
rect 4534 1168 4538 1172
rect 4542 1158 4546 1162
rect 4502 778 4506 782
rect 4510 748 4514 752
rect 4494 548 4498 552
rect 4486 348 4490 352
rect 4086 68 4090 72
rect 4582 2158 4586 2162
rect 4574 1998 4578 2002
rect 4574 1798 4578 1802
rect 4574 1728 4578 1732
rect 4582 1678 4586 1682
rect 4566 1418 4570 1422
rect 4574 1268 4578 1272
rect 4534 718 4538 722
rect 4582 1198 4586 1202
rect 4526 348 4530 352
rect 4518 138 4522 142
rect 4566 138 4570 142
rect 4438 68 4442 72
rect 4542 68 4546 72
rect 4634 4803 4638 4807
rect 4641 4803 4642 4807
rect 4642 4803 4645 4807
rect 4622 4668 4626 4672
rect 4634 4603 4638 4607
rect 4641 4603 4642 4607
rect 4642 4603 4645 4607
rect 4750 4548 4754 4552
rect 4634 4403 4638 4407
rect 4641 4403 4642 4407
rect 4642 4403 4645 4407
rect 4634 4203 4638 4207
rect 4641 4203 4642 4207
rect 4642 4203 4645 4207
rect 4622 4188 4626 4192
rect 4646 4158 4650 4162
rect 4622 4148 4626 4152
rect 4654 4088 4658 4092
rect 4634 4003 4638 4007
rect 4641 4003 4642 4007
rect 4642 4003 4645 4007
rect 4678 4218 4682 4222
rect 4694 4168 4698 4172
rect 4734 4078 4738 4082
rect 4678 4058 4682 4062
rect 4662 3988 4666 3992
rect 4702 3978 4706 3982
rect 4694 3928 4698 3932
rect 4634 3803 4638 3807
rect 4641 3803 4642 3807
rect 4642 3803 4645 3807
rect 4634 3603 4638 3607
rect 4641 3603 4642 3607
rect 4642 3603 4645 3607
rect 4634 3403 4638 3407
rect 4641 3403 4642 3407
rect 4642 3403 4645 3407
rect 4634 3203 4638 3207
rect 4641 3203 4642 3207
rect 4642 3203 4645 3207
rect 4614 2958 4618 2962
rect 4634 3003 4638 3007
rect 4641 3003 4642 3007
rect 4642 3003 4645 3007
rect 4630 2938 4634 2942
rect 4622 2868 4626 2872
rect 4634 2803 4638 2807
rect 4641 2803 4642 2807
rect 4642 2803 4645 2807
rect 4646 2788 4650 2792
rect 4710 3658 4714 3662
rect 4710 3548 4714 3552
rect 4710 3468 4714 3472
rect 4678 3448 4682 3452
rect 4718 3448 4722 3452
rect 4670 3298 4674 3302
rect 4662 3188 4666 3192
rect 4686 3138 4690 3142
rect 4686 2898 4690 2902
rect 4662 2788 4666 2792
rect 4634 2603 4638 2607
rect 4641 2603 4642 2607
rect 4642 2603 4645 2607
rect 4622 2568 4626 2572
rect 4654 2518 4658 2522
rect 4634 2403 4638 2407
rect 4641 2403 4642 2407
rect 4642 2403 4645 2407
rect 4654 2388 4658 2392
rect 4646 2308 4650 2312
rect 4638 2278 4642 2282
rect 4634 2203 4638 2207
rect 4641 2203 4642 2207
rect 4642 2203 4645 2207
rect 4634 2003 4638 2007
rect 4641 2003 4642 2007
rect 4642 2003 4645 2007
rect 4646 1968 4650 1972
rect 4662 2068 4666 2072
rect 4662 2018 4666 2022
rect 4654 1878 4658 1882
rect 4634 1803 4638 1807
rect 4641 1803 4642 1807
rect 4642 1803 4645 1807
rect 4614 1708 4618 1712
rect 4630 1678 4634 1682
rect 4614 1668 4618 1672
rect 4606 1588 4610 1592
rect 4598 1228 4602 1232
rect 4634 1603 4638 1607
rect 4641 1603 4642 1607
rect 4642 1603 4645 1607
rect 4654 1488 4658 1492
rect 4634 1403 4638 1407
rect 4641 1403 4642 1407
rect 4642 1403 4645 1407
rect 4634 1203 4638 1207
rect 4641 1203 4642 1207
rect 4642 1203 4645 1207
rect 4646 1148 4650 1152
rect 4634 1003 4638 1007
rect 4641 1003 4642 1007
rect 4642 1003 4645 1007
rect 4614 868 4618 872
rect 4634 803 4638 807
rect 4641 803 4642 807
rect 4642 803 4645 807
rect 4686 2558 4690 2562
rect 4678 2148 4682 2152
rect 4670 1918 4674 1922
rect 4702 2318 4706 2322
rect 4670 1668 4674 1672
rect 4686 1638 4690 1642
rect 4678 1268 4682 1272
rect 4630 768 4634 772
rect 4678 1088 4682 1092
rect 4670 958 4674 962
rect 4678 938 4682 942
rect 4634 603 4638 607
rect 4641 603 4642 607
rect 4642 603 4645 607
rect 4634 403 4638 407
rect 4641 403 4642 407
rect 4642 403 4645 407
rect 4702 2238 4706 2242
rect 4702 1958 4706 1962
rect 4758 4448 4762 4452
rect 4758 3938 4762 3942
rect 4758 3748 4762 3752
rect 4742 3488 4746 3492
rect 4750 3028 4754 3032
rect 4750 2858 4754 2862
rect 4758 2658 4762 2662
rect 4782 3358 4786 3362
rect 4862 4858 4866 4862
rect 4814 3958 4818 3962
rect 4854 4648 4858 4652
rect 4838 4318 4842 4322
rect 4766 2558 4770 2562
rect 4790 2548 4794 2552
rect 4742 2468 4746 2472
rect 4750 2268 4754 2272
rect 4734 1938 4738 1942
rect 4726 1878 4730 1882
rect 4718 1628 4722 1632
rect 4710 1588 4714 1592
rect 4726 1428 4730 1432
rect 4702 1178 4706 1182
rect 4694 1158 4698 1162
rect 4694 1018 4698 1022
rect 4694 938 4698 942
rect 4710 958 4714 962
rect 4710 938 4714 942
rect 4742 1488 4746 1492
rect 4766 2118 4770 2122
rect 4766 2108 4770 2112
rect 4766 1838 4770 1842
rect 4790 2158 4794 2162
rect 4758 1048 4762 1052
rect 4782 948 4786 952
rect 4766 858 4770 862
rect 4926 4858 4930 4862
rect 4886 4578 4890 4582
rect 4894 3338 4898 3342
rect 4894 3168 4898 3172
rect 4886 2948 4890 2952
rect 4830 2278 4834 2282
rect 4822 1878 4826 1882
rect 4750 668 4754 672
rect 4634 203 4638 207
rect 4641 203 4642 207
rect 4642 203 4645 207
rect 4814 1048 4818 1052
rect 4854 2468 4858 2472
rect 4862 1978 4866 1982
rect 4846 1868 4850 1872
rect 4846 1788 4850 1792
rect 4902 2888 4906 2892
rect 4894 2758 4898 2762
rect 4878 1918 4882 1922
rect 4870 1888 4874 1892
rect 4870 1868 4874 1872
rect 4870 1718 4874 1722
rect 4854 1698 4858 1702
rect 4862 1678 4866 1682
rect 4846 988 4850 992
rect 4838 938 4842 942
rect 4830 658 4834 662
rect 4598 108 4602 112
rect 4854 688 4858 692
rect 4862 258 4866 262
rect 4902 2148 4906 2152
rect 4910 2128 4914 2132
rect 4902 2098 4906 2102
rect 4982 4018 4986 4022
rect 4974 3358 4978 3362
rect 4966 3348 4970 3352
rect 4966 3338 4970 3342
rect 4942 3128 4946 3132
rect 4942 3078 4946 3082
rect 4918 1828 4922 1832
rect 4910 1758 4914 1762
rect 4918 1738 4922 1742
rect 4902 1568 4906 1572
rect 4942 2068 4946 2072
rect 4902 968 4906 972
rect 4942 888 4946 892
rect 4950 728 4954 732
rect 4974 1768 4978 1772
rect 4982 1728 4986 1732
rect 4966 728 4970 732
rect 4950 78 4954 82
rect 5030 4478 5034 4482
rect 5022 2918 5026 2922
rect 5030 2888 5034 2892
rect 5022 2778 5026 2782
rect 5054 4658 5058 4662
rect 5110 4858 5114 4862
rect 5070 4378 5074 4382
rect 5054 3348 5058 3352
rect 5086 4218 5090 4222
rect 5046 2638 5050 2642
rect 5014 2108 5018 2112
rect 5006 2088 5010 2092
rect 4998 2078 5002 2082
rect 4998 2058 5002 2062
rect 5014 1868 5018 1872
rect 5022 1718 5026 1722
rect 5014 1558 5018 1562
rect 5014 1238 5018 1242
rect 5078 2788 5082 2792
rect 5062 2308 5066 2312
rect 5062 2078 5066 2082
rect 5070 2068 5074 2072
rect 5166 3998 5170 4002
rect 5118 2958 5122 2962
rect 5110 2648 5114 2652
rect 5110 2628 5114 2632
rect 5094 2378 5098 2382
rect 5094 2358 5098 2362
rect 5126 2568 5130 2572
rect 5126 2548 5130 2552
rect 5118 2538 5122 2542
rect 5158 3048 5162 3052
rect 5142 2658 5146 2662
rect 5134 2468 5138 2472
rect 5134 2428 5138 2432
rect 5102 2338 5106 2342
rect 5054 1498 5058 1502
rect 5038 648 5042 652
rect 5006 578 5010 582
rect 5062 738 5066 742
rect 5086 1488 5090 1492
rect 5094 1258 5098 1262
rect 5142 2278 5146 2282
rect 5134 2038 5138 2042
rect 5166 2638 5170 2642
rect 5158 2418 5162 2422
rect 5150 2258 5154 2262
rect 5110 188 5114 192
rect 5014 88 5018 92
rect 5190 2758 5194 2762
rect 5182 2668 5186 2672
rect 5182 2648 5186 2652
rect 5166 2028 5170 2032
rect 5166 928 5170 932
rect 5190 2068 5194 2072
rect 5182 858 5186 862
rect 5182 288 5186 292
rect 4694 58 4698 62
rect 4758 58 4762 62
rect 5142 58 5146 62
rect 4046 48 4050 52
rect 4126 48 4130 52
rect 4558 48 4562 52
rect 4822 48 4826 52
rect 538 3 542 7
rect 545 3 546 7
rect 546 3 549 7
rect 1562 3 1566 7
rect 1569 3 1570 7
rect 1570 3 1573 7
rect 2586 3 2590 7
rect 2593 3 2594 7
rect 2594 3 2597 7
rect 3610 3 3614 7
rect 3617 3 3618 7
rect 3618 3 3621 7
rect 4634 3 4638 7
rect 4641 3 4642 7
rect 4642 3 4645 7
<< metal5 >>
rect 1054 4903 1057 4907
rect 1053 4902 1058 4903
rect 1063 4902 1064 4907
rect 2078 4903 2081 4907
rect 2077 4902 2082 4903
rect 2087 4902 2088 4907
rect 3102 4903 3105 4907
rect 3101 4902 3106 4903
rect 3111 4902 3112 4907
rect 4118 4903 4121 4907
rect 4117 4902 4122 4903
rect 4127 4902 4128 4907
rect 586 4858 766 4861
rect 770 4858 1246 4861
rect 1250 4858 1542 4861
rect 2378 4858 2381 4861
rect 4862 4852 4865 4858
rect 4926 4852 4929 4858
rect 5106 4858 5110 4861
rect 542 4803 545 4807
rect 541 4802 546 4803
rect 551 4802 552 4807
rect 1566 4803 1569 4807
rect 1565 4802 1570 4803
rect 1575 4802 1576 4807
rect 2590 4803 2593 4807
rect 2589 4802 2594 4803
rect 2599 4802 2600 4807
rect 3614 4803 3617 4807
rect 3613 4802 3618 4803
rect 3623 4802 3624 4807
rect 4638 4803 4641 4807
rect 4637 4802 4642 4803
rect 4647 4802 4648 4807
rect 674 4748 1222 4751
rect 1226 4748 1350 4751
rect 1506 4748 1630 4751
rect 1626 4738 1702 4741
rect 2666 4738 3006 4741
rect 1682 4728 2030 4731
rect 1054 4703 1057 4707
rect 1053 4702 1058 4703
rect 1063 4702 1064 4707
rect 2078 4703 2081 4707
rect 2077 4702 2082 4703
rect 2087 4702 2088 4707
rect 3102 4703 3105 4707
rect 3101 4702 3106 4703
rect 3111 4702 3112 4707
rect 4118 4703 4121 4707
rect 4117 4702 4122 4703
rect 4127 4702 4128 4707
rect 498 4688 1206 4691
rect 1210 4688 2550 4691
rect 1154 4678 1334 4681
rect 4626 4668 5057 4671
rect 5054 4662 5057 4668
rect 1202 4658 1382 4661
rect 2722 4658 3038 4661
rect 3042 4658 3550 4661
rect 154 4648 422 4651
rect 426 4648 1542 4651
rect 1962 4648 3030 4651
rect 3034 4648 3406 4651
rect 4210 4648 4854 4651
rect 1314 4638 1597 4641
rect 1602 4638 3294 4641
rect 542 4603 545 4607
rect 541 4602 546 4603
rect 551 4602 552 4607
rect 1566 4603 1569 4607
rect 1565 4602 1570 4603
rect 1575 4602 1576 4607
rect 2590 4603 2593 4607
rect 2589 4602 2594 4603
rect 2599 4602 2600 4607
rect 3614 4603 3617 4607
rect 3613 4602 3618 4603
rect 3623 4602 3624 4607
rect 4638 4603 4641 4607
rect 4637 4602 4642 4603
rect 4647 4602 4648 4607
rect 4562 4578 4886 4581
rect 1386 4548 3262 4551
rect 3498 4548 4750 4551
rect 746 4538 749 4541
rect 1498 4538 1630 4541
rect 2570 4538 2998 4541
rect 4482 4538 4518 4541
rect 866 4528 1278 4531
rect 1450 4528 1534 4531
rect 1634 4528 1718 4531
rect 1722 4528 2494 4531
rect 2506 4528 2990 4531
rect 3546 4528 4310 4531
rect 4314 4528 4430 4531
rect 322 4518 1190 4521
rect 1578 4518 2246 4521
rect 3530 4518 3549 4521
rect 3554 4518 4494 4521
rect 1054 4503 1057 4507
rect 1053 4502 1058 4503
rect 1063 4502 1064 4507
rect 2078 4503 2081 4507
rect 2077 4502 2082 4503
rect 2087 4502 2088 4507
rect 3102 4503 3105 4507
rect 3101 4502 3106 4503
rect 3111 4502 3112 4507
rect 4118 4503 4121 4507
rect 4117 4502 4122 4503
rect 4127 4502 4128 4507
rect 1922 4478 2422 4481
rect 3538 4478 5030 4481
rect 658 4468 2030 4471
rect 2258 4468 2710 4471
rect 3522 4468 4761 4471
rect 1170 4458 2238 4461
rect 2242 4458 3918 4461
rect 4090 4458 4606 4461
rect 4758 4461 4761 4468
rect 4754 4458 4761 4461
rect 4758 4452 4761 4458
rect 634 4448 1598 4451
rect 1602 4448 1661 4451
rect 2074 4448 2374 4451
rect 2734 4442 2737 4448
rect 3202 4438 3822 4441
rect 2338 4428 2366 4431
rect 2882 4428 4150 4431
rect 1458 4418 1590 4421
rect 1594 4418 2270 4421
rect 2274 4418 3150 4421
rect 4398 4412 4401 4418
rect 2618 4408 3198 4411
rect 542 4403 545 4407
rect 541 4402 546 4403
rect 551 4402 552 4407
rect 1566 4403 1569 4407
rect 1565 4402 1570 4403
rect 1575 4402 1576 4407
rect 2590 4403 2593 4407
rect 2589 4402 2594 4403
rect 2599 4402 2600 4407
rect 3614 4403 3617 4407
rect 3613 4402 3618 4403
rect 3623 4402 3624 4407
rect 4542 4402 4545 4408
rect 4638 4403 4641 4407
rect 4637 4402 4642 4403
rect 4647 4402 4648 4407
rect 1810 4388 1846 4391
rect 1850 4388 3549 4391
rect 1978 4378 3366 4381
rect 5070 4372 5073 4378
rect 1858 4368 2717 4371
rect 2738 4368 4446 4371
rect 1090 4358 2390 4361
rect 282 4348 493 4351
rect 498 4348 2174 4351
rect 2538 4348 2550 4351
rect 3946 4348 4086 4351
rect 1466 4338 2798 4341
rect 2834 4338 3174 4341
rect 3178 4338 3318 4341
rect 3330 4338 3766 4341
rect 3770 4338 4278 4341
rect 4558 4332 4561 4337
rect 714 4328 998 4331
rect 1002 4328 2342 4331
rect 2722 4328 4022 4331
rect 554 4318 781 4321
rect 786 4318 1494 4321
rect 1498 4318 1678 4321
rect 1682 4318 2846 4321
rect 3154 4318 4838 4321
rect 2186 4308 2189 4311
rect 3938 4308 3990 4311
rect 1054 4303 1057 4307
rect 1053 4302 1058 4303
rect 1063 4302 1064 4307
rect 2078 4303 2081 4307
rect 2077 4302 2082 4303
rect 2087 4302 2088 4307
rect 3102 4303 3105 4307
rect 3101 4302 3106 4303
rect 3111 4302 3112 4307
rect 4118 4303 4121 4307
rect 4117 4302 4122 4303
rect 4127 4302 4128 4307
rect 634 4288 1150 4291
rect 2378 4288 3214 4291
rect 1178 4278 2134 4281
rect 2970 4278 3030 4281
rect 3034 4278 3790 4281
rect 4042 4278 4158 4281
rect 2138 4268 3533 4271
rect 3882 4268 4049 4271
rect 4066 4268 4606 4271
rect 4046 4262 4049 4268
rect 818 4258 1822 4261
rect 2182 4251 2185 4258
rect 2562 4258 2630 4261
rect 3282 4258 4041 4261
rect 4266 4258 4269 4261
rect 4038 4252 4041 4258
rect 266 4248 2185 4251
rect 2482 4248 3430 4251
rect 3538 4248 3942 4251
rect 4018 4248 4022 4251
rect 858 4238 1006 4241
rect 1010 4238 2294 4241
rect 3146 4238 3902 4241
rect 1418 4228 2477 4231
rect 2770 4228 3598 4231
rect 3794 4228 4397 4231
rect 2666 4218 2926 4221
rect 3298 4218 4045 4221
rect 4050 4218 4678 4221
rect 4682 4218 5086 4221
rect 542 4203 545 4207
rect 541 4202 546 4203
rect 551 4202 552 4207
rect 1566 4203 1569 4207
rect 1565 4202 1570 4203
rect 1575 4202 1576 4207
rect 2590 4203 2593 4207
rect 2589 4202 2594 4203
rect 2599 4202 2600 4207
rect 3134 4202 3137 4208
rect 3614 4203 3617 4207
rect 3613 4202 3618 4203
rect 3623 4202 3624 4207
rect 4638 4203 4641 4207
rect 4637 4202 4642 4203
rect 4647 4202 4648 4207
rect 1914 4188 2806 4191
rect 2946 4188 3437 4191
rect 3442 4188 3630 4191
rect 4622 4182 4625 4188
rect 370 4178 1750 4181
rect 2354 4178 3133 4181
rect 1378 4168 2173 4171
rect 2326 4171 2329 4178
rect 2178 4168 2329 4171
rect 4602 4168 4694 4171
rect 1498 4158 2941 4161
rect 2954 4158 3710 4161
rect 4546 4158 4646 4161
rect 794 4148 1398 4151
rect 1410 4148 1718 4151
rect 2422 4148 2822 4151
rect 3130 4148 3726 4151
rect 4538 4148 4622 4151
rect 2422 4142 2425 4148
rect 426 4138 1510 4141
rect 2850 4138 3406 4141
rect 3986 4138 3990 4141
rect 4530 4138 4553 4141
rect 4550 4132 4553 4138
rect 898 4128 1710 4131
rect 3130 4128 3566 4131
rect 3570 4128 4070 4131
rect 1234 4118 1261 4121
rect 2394 4118 3990 4121
rect 306 4108 966 4111
rect 3434 4108 3558 4111
rect 1054 4103 1057 4107
rect 1053 4102 1058 4103
rect 1063 4102 1064 4107
rect 2078 4103 2081 4107
rect 2077 4102 2082 4103
rect 2087 4102 2088 4107
rect 3102 4103 3105 4107
rect 3101 4102 3106 4103
rect 3111 4102 3112 4107
rect 4118 4103 4121 4107
rect 4117 4102 4122 4103
rect 4127 4102 4128 4107
rect 2218 4098 2782 4101
rect 3474 4088 3990 4091
rect 4010 4088 4654 4091
rect 394 4078 1214 4081
rect 1234 4078 2425 4081
rect 2778 4078 3238 4081
rect 4098 4078 4734 4081
rect 2422 4072 2425 4078
rect 790 4068 798 4071
rect 802 4068 966 4071
rect 1162 4068 1726 4071
rect 2442 4068 2830 4071
rect 3186 4068 4318 4071
rect 322 4058 1406 4061
rect 1906 4058 2222 4061
rect 2226 4058 2342 4061
rect 2358 4061 2361 4068
rect 2358 4058 2365 4061
rect 2554 4058 2830 4061
rect 2898 4058 3230 4061
rect 3258 4058 3942 4061
rect 3962 4058 4230 4061
rect 4234 4058 4678 4061
rect 906 4048 1622 4051
rect 1634 4048 2134 4051
rect 2138 4048 3790 4051
rect 4050 4048 4061 4051
rect 4098 4048 4101 4051
rect 930 4038 1526 4041
rect 2026 4038 2829 4041
rect 2834 4038 3486 4041
rect 3746 4038 4174 4041
rect 570 4028 878 4031
rect 1258 4028 1270 4031
rect 1274 4028 1894 4031
rect 2370 4028 3806 4031
rect 386 4018 1806 4021
rect 1970 4018 2998 4021
rect 3674 4018 3878 4021
rect 4978 4018 4982 4021
rect 2658 4008 3342 4011
rect 542 4003 545 4007
rect 541 4002 546 4003
rect 551 4002 552 4007
rect 1566 4003 1569 4007
rect 1565 4002 1570 4003
rect 1575 4002 1576 4007
rect 2590 4003 2593 4007
rect 2589 4002 2594 4003
rect 2599 4002 2600 4007
rect 3614 4003 3617 4007
rect 3613 4002 3618 4003
rect 3623 4002 3624 4007
rect 4638 4003 4641 4007
rect 4637 4002 4642 4003
rect 4647 4002 4648 4007
rect 1842 3998 2166 4001
rect 2610 3998 2846 4001
rect 2994 3998 3470 4001
rect 5154 3998 5166 4001
rect 1026 3988 3566 3991
rect 3618 3988 4662 3991
rect 1082 3978 3278 3981
rect 3346 3978 3750 3981
rect 4226 3978 4702 3981
rect 594 3968 1158 3971
rect 1174 3968 1182 3971
rect 1186 3968 1214 3971
rect 1226 3968 2350 3971
rect 2994 3968 3454 3971
rect 3666 3968 3918 3971
rect 3922 3968 4294 3971
rect 274 3958 1214 3961
rect 1290 3958 2241 3961
rect 2266 3958 2493 3961
rect 2238 3951 2241 3958
rect 2850 3958 2878 3961
rect 2954 3958 3534 3961
rect 4154 3958 4222 3961
rect 4390 3958 4398 3961
rect 4402 3958 4814 3961
rect 2238 3948 3046 3951
rect 3298 3948 4038 3951
rect 722 3938 1446 3941
rect 1746 3938 3630 3941
rect 4762 3938 4765 3941
rect 1106 3928 2166 3931
rect 2186 3928 2873 3931
rect 2890 3928 4230 3931
rect 1098 3918 2326 3921
rect 2602 3918 2758 3921
rect 2826 3918 2862 3921
rect 2870 3921 2873 3928
rect 4578 3928 4694 3931
rect 2870 3918 3134 3921
rect 3390 3912 3393 3918
rect 1450 3908 2061 3911
rect 2298 3908 3078 3911
rect 1054 3903 1057 3907
rect 1053 3902 1058 3903
rect 1063 3902 1064 3907
rect 2078 3903 2081 3907
rect 2077 3902 2082 3903
rect 2087 3902 2088 3907
rect 3102 3903 3105 3907
rect 3101 3902 3106 3903
rect 3111 3902 3112 3907
rect 4118 3903 4121 3907
rect 4117 3902 4122 3903
rect 4127 3902 4128 3907
rect 1482 3898 2062 3901
rect 2130 3898 2726 3901
rect 3118 3898 3958 3901
rect 910 3892 913 3898
rect 1282 3888 1862 3891
rect 3118 3891 3121 3898
rect 2402 3888 3121 3891
rect 3722 3888 4182 3891
rect 1154 3878 1894 3881
rect 3434 3878 4254 3881
rect 418 3868 797 3871
rect 802 3868 1566 3871
rect 1574 3868 2182 3871
rect 2426 3868 2622 3871
rect 3370 3868 4062 3871
rect 4562 3868 4606 3871
rect 1574 3861 1577 3868
rect 282 3858 1577 3861
rect 2426 3858 3342 3861
rect 3482 3858 3694 3861
rect 4202 3858 4221 3861
rect 4450 3858 4574 3861
rect 1554 3848 1558 3851
rect 1562 3848 2702 3851
rect 3570 3848 4222 3851
rect 4322 3848 4550 3851
rect 674 3838 2318 3841
rect 2378 3838 3382 3841
rect 3410 3838 4285 3841
rect 4290 3838 4358 3841
rect 1818 3828 2902 3831
rect 3338 3828 4262 3831
rect 770 3818 2413 3821
rect 2418 3818 3070 3821
rect 3602 3818 3614 3821
rect 1722 3808 2238 3811
rect 2310 3808 2318 3811
rect 2322 3808 2406 3811
rect 3042 3808 3213 3811
rect 4498 3808 4509 3811
rect 542 3803 545 3807
rect 541 3802 546 3803
rect 551 3802 552 3807
rect 1566 3803 1569 3807
rect 1565 3802 1570 3803
rect 1575 3802 1576 3807
rect 2590 3803 2593 3807
rect 2589 3802 2594 3803
rect 2599 3802 2600 3807
rect 3614 3803 3617 3807
rect 3613 3802 3618 3803
rect 3623 3802 3624 3807
rect 4638 3803 4641 3807
rect 4637 3802 4642 3803
rect 4647 3802 4648 3807
rect 1866 3798 2326 3801
rect 2650 3798 3558 3801
rect 1858 3788 2157 3791
rect 2622 3788 3670 3791
rect 2010 3778 2030 3781
rect 2622 3781 2625 3788
rect 2154 3778 2625 3781
rect 2634 3778 3734 3781
rect 1714 3768 1725 3771
rect 1986 3768 2390 3771
rect 2434 3768 2934 3771
rect 1914 3758 2646 3761
rect 2690 3758 3485 3761
rect 3522 3758 3902 3761
rect 1674 3748 1694 3751
rect 3518 3751 3521 3758
rect 3090 3748 3521 3751
rect 4578 3748 4758 3751
rect 382 3742 385 3747
rect 2030 3742 2033 3748
rect 1186 3738 1933 3741
rect 2442 3738 4318 3741
rect 1674 3728 1949 3731
rect 1954 3728 2397 3731
rect 3530 3728 3533 3731
rect 3586 3728 4046 3731
rect 1410 3718 1438 3721
rect 1514 3718 1670 3721
rect 1690 3718 1750 3721
rect 1994 3718 2030 3721
rect 2066 3718 3214 3721
rect 3226 3718 3725 3721
rect 3730 3718 4510 3721
rect 1314 3708 1590 3711
rect 2098 3708 2221 3711
rect 2226 3708 2989 3711
rect 1054 3703 1057 3707
rect 1053 3702 1058 3703
rect 1063 3702 1064 3707
rect 2078 3703 2081 3707
rect 2077 3702 2082 3703
rect 2087 3702 2088 3707
rect 3102 3703 3105 3707
rect 3101 3702 3106 3703
rect 3111 3702 3112 3707
rect 4118 3703 4121 3707
rect 4117 3702 4122 3703
rect 4127 3702 4128 3707
rect 1034 3698 1037 3701
rect 670 3692 673 3698
rect 1714 3698 1721 3701
rect 1598 3692 1601 3697
rect 1718 3692 1721 3698
rect 2322 3698 3086 3701
rect 1762 3688 2230 3691
rect 2234 3688 2254 3691
rect 2282 3688 2494 3691
rect 3394 3688 3638 3691
rect 3722 3688 4190 3691
rect 2750 3682 2753 3688
rect 1362 3678 1534 3681
rect 1538 3678 1734 3681
rect 1754 3678 2317 3681
rect 478 3671 481 3678
rect 3490 3678 3702 3681
rect 478 3668 998 3671
rect 1202 3668 1902 3671
rect 2362 3668 2478 3671
rect 2570 3668 3118 3671
rect 3450 3668 3734 3671
rect 1770 3658 2998 3661
rect 3050 3658 3069 3661
rect 3254 3661 3257 3668
rect 3074 3658 3257 3661
rect 3954 3658 3990 3661
rect 4594 3658 4710 3661
rect 1146 3648 1814 3651
rect 1826 3648 2670 3651
rect 2674 3648 3878 3651
rect 3882 3648 4333 3651
rect 4338 3648 4358 3651
rect 1090 3638 1126 3641
rect 1130 3638 1942 3641
rect 3378 3638 3454 3641
rect 3546 3638 3830 3641
rect 4082 3638 4102 3641
rect 1114 3628 1406 3631
rect 1858 3628 1926 3631
rect 1930 3628 3342 3631
rect 3346 3628 3757 3631
rect 3762 3628 3766 3631
rect 1010 3618 1750 3621
rect 2482 3618 3405 3621
rect 2290 3608 2294 3611
rect 2354 3608 2477 3611
rect 3522 3608 3590 3611
rect 4458 3608 4573 3611
rect 542 3603 545 3607
rect 541 3602 546 3603
rect 551 3602 552 3607
rect 1566 3603 1569 3607
rect 1565 3602 1570 3603
rect 1575 3602 1576 3607
rect 2590 3603 2593 3607
rect 2589 3602 2594 3603
rect 2599 3602 2600 3607
rect 3614 3603 3617 3607
rect 3613 3602 3618 3603
rect 3623 3602 3624 3607
rect 4638 3603 4641 3607
rect 4637 3602 4642 3603
rect 4647 3602 4648 3607
rect 1074 3598 1230 3601
rect 1314 3598 1318 3601
rect 1674 3598 2093 3601
rect 3154 3598 3542 3601
rect 4002 3598 4022 3601
rect 1610 3588 2614 3591
rect 3138 3588 3478 3591
rect 3482 3588 4269 3591
rect 682 3578 1630 3581
rect 1746 3578 1750 3581
rect 2098 3578 3406 3581
rect 3954 3578 4062 3581
rect 834 3568 1310 3571
rect 2506 3568 3182 3571
rect 3218 3568 3421 3571
rect 3426 3568 4310 3571
rect 346 3558 358 3561
rect 362 3558 1638 3561
rect 1714 3558 1758 3561
rect 2058 3558 3645 3561
rect 3666 3558 3677 3561
rect 618 3548 686 3551
rect 690 3548 1318 3551
rect 1426 3548 1630 3551
rect 1762 3548 2441 3551
rect 2858 3548 3206 3551
rect 3210 3548 3302 3551
rect 3314 3548 4710 3551
rect 2438 3542 2441 3548
rect 1026 3538 1302 3541
rect 1330 3538 1494 3541
rect 1666 3538 2350 3541
rect 3018 3538 4118 3541
rect 1490 3528 1774 3531
rect 2402 3528 2574 3531
rect 2962 3528 3582 3531
rect 3818 3528 4430 3531
rect 4434 3528 4550 3531
rect 1418 3518 1430 3521
rect 1434 3518 1437 3521
rect 1458 3518 2422 3521
rect 2618 3518 4470 3521
rect 1266 3508 1598 3511
rect 3386 3508 3814 3511
rect 3914 3508 3917 3511
rect 4274 3508 4302 3511
rect 1054 3503 1057 3507
rect 1053 3502 1058 3503
rect 1063 3502 1064 3507
rect 2078 3503 2081 3507
rect 2077 3502 2082 3503
rect 2087 3502 2088 3507
rect 3102 3503 3105 3507
rect 3101 3502 3106 3503
rect 3111 3502 3112 3507
rect 4118 3503 4121 3507
rect 4117 3502 4122 3503
rect 4127 3502 4128 3507
rect 482 3498 502 3501
rect 1458 3498 1469 3501
rect 1474 3498 1830 3501
rect 2170 3498 2173 3501
rect 2546 3498 2558 3501
rect 3794 3498 3821 3501
rect 1122 3488 1821 3491
rect 1878 3488 2478 3491
rect 2522 3488 3470 3491
rect 3482 3488 4742 3491
rect 250 3478 446 3481
rect 450 3478 765 3481
rect 770 3478 1326 3481
rect 1878 3481 1881 3488
rect 1418 3478 1881 3481
rect 2394 3478 2678 3481
rect 2970 3478 3102 3481
rect 3106 3478 3294 3481
rect 1042 3468 1453 3471
rect 1474 3468 1534 3471
rect 1682 3468 2541 3471
rect 1002 3458 1069 3461
rect 1274 3458 1390 3461
rect 1522 3458 1622 3461
rect 1630 3461 1633 3468
rect 2818 3468 3629 3471
rect 3898 3468 4342 3471
rect 4370 3468 4373 3471
rect 4690 3468 4710 3471
rect 4398 3462 4401 3467
rect 1630 3458 1718 3461
rect 1722 3458 2118 3461
rect 2386 3458 2390 3461
rect 2890 3458 3326 3461
rect 682 3448 685 3451
rect 866 3448 1862 3451
rect 1994 3448 2078 3451
rect 3154 3448 3742 3451
rect 3954 3448 3982 3451
rect 4682 3448 4718 3451
rect 1402 3438 1917 3441
rect 1922 3438 2102 3441
rect 2114 3438 3782 3441
rect 1154 3428 1277 3431
rect 1338 3428 3597 3431
rect 722 3418 877 3421
rect 962 3418 1357 3421
rect 1378 3418 1510 3421
rect 1586 3418 1654 3421
rect 1786 3418 1789 3421
rect 2242 3418 3574 3421
rect 730 3408 733 3411
rect 1138 3408 1142 3411
rect 542 3403 545 3407
rect 541 3402 546 3403
rect 551 3402 552 3407
rect 1566 3403 1569 3407
rect 1565 3402 1570 3403
rect 1575 3402 1576 3407
rect 2590 3403 2593 3407
rect 2589 3402 2594 3403
rect 2599 3402 2600 3407
rect 3614 3403 3617 3407
rect 3613 3402 3618 3403
rect 3623 3402 3624 3407
rect 4638 3403 4641 3407
rect 4637 3402 4642 3403
rect 4647 3402 4648 3407
rect 690 3398 1486 3401
rect 3314 3398 3382 3401
rect 2970 3388 4557 3391
rect 1714 3378 2758 3381
rect 2770 3378 3798 3381
rect 3802 3378 3862 3381
rect 2386 3368 3293 3371
rect 4570 3368 4590 3371
rect 138 3358 550 3361
rect 698 3358 726 3361
rect 1490 3358 1718 3361
rect 2034 3358 2038 3361
rect 2946 3358 4510 3361
rect 4786 3358 4974 3361
rect 1274 3348 1629 3351
rect 1634 3348 2046 3351
rect 2290 3348 2502 3351
rect 2554 3348 2678 3351
rect 2906 3348 3494 3351
rect 3938 3348 4238 3351
rect 4590 3351 4593 3358
rect 4242 3348 4593 3351
rect 4970 3348 5054 3351
rect 1182 3338 1197 3341
rect 1182 3332 1185 3338
rect 1298 3338 1702 3341
rect 1722 3338 2462 3341
rect 2490 3338 2814 3341
rect 3970 3338 4477 3341
rect 4482 3338 4541 3341
rect 4546 3338 4574 3341
rect 4898 3338 4966 3341
rect 170 3328 518 3331
rect 522 3328 646 3331
rect 650 3328 990 3331
rect 1098 3328 1182 3331
rect 1258 3328 1406 3331
rect 1458 3328 1462 3331
rect 1970 3328 2029 3331
rect 2130 3328 3246 3331
rect 3498 3328 3622 3331
rect 3742 3328 3910 3331
rect 3930 3328 4150 3331
rect 4154 3328 4518 3331
rect 3742 3322 3745 3328
rect 434 3318 518 3321
rect 1650 3318 2142 3321
rect 2898 3318 3142 3321
rect 2558 3312 2561 3318
rect 1210 3308 1294 3311
rect 1298 3308 1350 3311
rect 1362 3308 1630 3311
rect 4210 3308 4262 3311
rect 1054 3303 1057 3307
rect 1053 3302 1058 3303
rect 1063 3302 1064 3307
rect 2078 3303 2081 3307
rect 2077 3302 2082 3303
rect 2087 3302 2088 3307
rect 3102 3303 3105 3307
rect 3101 3302 3106 3303
rect 3111 3302 3112 3307
rect 4118 3303 4121 3307
rect 4117 3302 4122 3303
rect 4127 3302 4128 3307
rect 1186 3298 1502 3301
rect 1690 3298 1757 3301
rect 2130 3298 2630 3301
rect 2634 3298 3054 3301
rect 3146 3298 3966 3301
rect 4034 3298 4038 3301
rect 4210 3298 4422 3301
rect 4426 3298 4670 3301
rect 946 3288 949 3291
rect 986 3288 1694 3291
rect 1826 3288 2278 3291
rect 2290 3288 2742 3291
rect 2746 3288 4438 3291
rect 274 3278 662 3281
rect 674 3278 1629 3281
rect 1642 3278 1822 3281
rect 1826 3278 2125 3281
rect 2658 3278 3197 3281
rect 3458 3278 3646 3281
rect 3986 3278 3990 3281
rect 4042 3278 4542 3281
rect 4546 3278 4590 3281
rect 890 3268 1590 3271
rect 1634 3268 2110 3271
rect 2250 3268 2318 3271
rect 2322 3268 3022 3271
rect 3090 3268 3678 3271
rect 3970 3268 4222 3271
rect 338 3258 925 3261
rect 1814 3258 2462 3261
rect 2514 3258 2669 3261
rect 1814 3251 1817 3258
rect 3066 3258 3198 3261
rect 3522 3258 4382 3261
rect 1498 3248 1817 3251
rect 2002 3248 2870 3251
rect 3042 3248 3718 3251
rect 3746 3248 3758 3251
rect 3762 3248 3966 3251
rect 770 3238 957 3241
rect 1954 3238 2013 3241
rect 2018 3238 2126 3241
rect 2194 3238 3894 3241
rect 858 3228 918 3231
rect 1138 3228 1341 3231
rect 1482 3228 1485 3231
rect 1634 3228 2701 3231
rect 3330 3228 4390 3231
rect 754 3218 910 3221
rect 1458 3218 1910 3221
rect 2162 3218 2214 3221
rect 2274 3218 2814 3221
rect 1326 3212 1329 3218
rect 3378 3218 4238 3221
rect 954 3208 1149 3211
rect 1714 3208 1718 3211
rect 1938 3208 2334 3211
rect 2658 3208 3270 3211
rect 3274 3208 3446 3211
rect 542 3203 545 3207
rect 541 3202 546 3203
rect 551 3202 552 3207
rect 1566 3203 1569 3207
rect 1565 3202 1570 3203
rect 1575 3202 1576 3207
rect 2590 3203 2593 3207
rect 2589 3202 2594 3203
rect 2599 3202 2600 3207
rect 3614 3203 3617 3207
rect 3613 3202 3618 3203
rect 3623 3202 3624 3207
rect 4638 3203 4641 3207
rect 4637 3202 4642 3203
rect 4647 3202 4648 3207
rect 578 3198 1494 3201
rect 1586 3198 2397 3201
rect 2754 3198 3590 3201
rect 474 3188 998 3191
rect 1098 3188 2382 3191
rect 2450 3188 3118 3191
rect 4250 3188 4662 3191
rect 778 3178 829 3181
rect 1074 3178 2094 3181
rect 2098 3178 2733 3181
rect 2738 3178 2966 3181
rect 2978 3178 4525 3181
rect 1130 3168 1158 3171
rect 1202 3168 1382 3171
rect 1394 3168 2318 3171
rect 2426 3168 2614 3171
rect 3994 3168 4894 3171
rect 3470 3162 3473 3168
rect 378 3158 774 3161
rect 994 3158 1134 3161
rect 1162 3158 1293 3161
rect 1298 3158 1550 3161
rect 1730 3158 1773 3161
rect 1914 3158 1974 3161
rect 1986 3158 2141 3161
rect 2510 3158 3374 3161
rect 26 3148 710 3151
rect 722 3148 734 3151
rect 738 3148 1494 3151
rect 1538 3148 1953 3151
rect 2510 3151 2513 3158
rect 4018 3158 4022 3161
rect 2066 3148 2513 3151
rect 3002 3148 3969 3151
rect 4018 3148 4270 3151
rect 1950 3142 1953 3148
rect 682 3138 990 3141
rect 1154 3138 1165 3141
rect 1178 3138 1486 3141
rect 2026 3138 2061 3141
rect 2114 3138 2662 3141
rect 2934 3141 2937 3148
rect 2966 3141 2969 3148
rect 2934 3138 2969 3141
rect 2978 3138 3430 3141
rect 3450 3138 3462 3141
rect 3586 3138 3750 3141
rect 3966 3141 3969 3148
rect 4530 3148 4534 3151
rect 3966 3138 4686 3141
rect 4690 3138 4733 3141
rect 818 3128 1421 3131
rect 1978 3128 2022 3131
rect 2026 3128 2510 3131
rect 3202 3128 3462 3131
rect 3578 3128 3902 3131
rect 4042 3128 4942 3131
rect 714 3118 1374 3121
rect 1746 3118 1837 3121
rect 1922 3118 1982 3121
rect 2058 3118 2285 3121
rect 2418 3118 2470 3121
rect 2626 3118 2685 3121
rect 3050 3118 3133 3121
rect 3138 3118 4318 3121
rect 818 3108 982 3111
rect 1370 3108 1742 3111
rect 2106 3108 2518 3111
rect 2626 3108 2918 3111
rect 2922 3108 2941 3111
rect 3434 3108 4014 3111
rect 4074 3108 4102 3111
rect 1054 3103 1057 3107
rect 1053 3102 1058 3103
rect 1063 3102 1064 3107
rect 2078 3103 2081 3107
rect 2077 3102 2082 3103
rect 2087 3102 2088 3107
rect 3102 3103 3105 3107
rect 3101 3102 3106 3103
rect 3111 3102 3112 3107
rect 4118 3103 4121 3107
rect 4117 3102 4122 3103
rect 4127 3102 4128 3107
rect 2106 3098 2134 3101
rect 2306 3098 2990 3101
rect 762 3088 1485 3091
rect 1666 3088 2001 3091
rect 2010 3088 2062 3091
rect 1002 3078 1694 3081
rect 1998 3081 2001 3088
rect 2274 3088 2294 3091
rect 2538 3088 2574 3091
rect 1998 3078 2502 3081
rect 2530 3078 3006 3081
rect 3830 3081 3833 3088
rect 3810 3078 3833 3081
rect 4018 3078 4942 3081
rect 178 3068 846 3071
rect 2050 3068 2486 3071
rect 2522 3068 3046 3071
rect 3186 3068 3190 3071
rect 3530 3068 3838 3071
rect 3914 3068 3917 3071
rect 3326 3062 3329 3067
rect 778 3058 1414 3061
rect 1602 3058 1670 3061
rect 1978 3058 2301 3061
rect 3442 3058 4142 3061
rect 4262 3061 4265 3068
rect 4262 3058 4342 3061
rect 978 3048 1534 3051
rect 1618 3048 1694 3051
rect 1738 3048 2182 3051
rect 2298 3048 2438 3051
rect 2506 3048 2686 3051
rect 2866 3048 3078 3051
rect 3826 3048 4526 3051
rect 5162 3048 5165 3051
rect 934 3038 1213 3041
rect 934 3032 937 3038
rect 1266 3038 1294 3041
rect 1730 3038 1734 3041
rect 1794 3038 2230 3041
rect 2538 3038 2758 3041
rect 3842 3038 4158 3041
rect 4490 3038 4582 3041
rect 946 3028 950 3031
rect 1354 3028 1357 3031
rect 1362 3028 1694 3031
rect 1698 3028 1974 3031
rect 2618 3028 4157 3031
rect 4162 3028 4750 3031
rect 1042 3018 1190 3021
rect 1218 3018 1929 3021
rect 1946 3018 1981 3021
rect 714 3008 1446 3011
rect 1926 3011 1929 3018
rect 2050 3018 2726 3021
rect 2738 3018 4093 3021
rect 4098 3018 4206 3021
rect 1926 3008 2221 3011
rect 2610 3008 2749 3011
rect 2754 3008 3518 3011
rect 3730 3008 4189 3011
rect 4194 3008 4286 3011
rect 542 3003 545 3007
rect 541 3002 546 3003
rect 551 3002 552 3007
rect 1566 3003 1569 3007
rect 1565 3002 1570 3003
rect 1575 3002 1576 3007
rect 2590 3003 2593 3007
rect 2589 3002 2594 3003
rect 2599 3002 2600 3007
rect 3614 3003 3617 3007
rect 3613 3002 3618 3003
rect 3623 3002 3624 3007
rect 4638 3003 4641 3007
rect 4637 3002 4642 3003
rect 4647 3002 4648 3007
rect 666 2998 1246 3001
rect 1586 2998 1950 3001
rect 1970 2998 1982 3001
rect 2170 2998 2573 3001
rect 2666 2998 3190 3001
rect 4026 2998 4045 3001
rect 1218 2988 1222 2991
rect 1338 2988 2262 2991
rect 2362 2988 3502 2991
rect 3554 2988 3933 2991
rect 3938 2988 3990 2991
rect 4258 2988 4494 2991
rect 946 2978 1014 2981
rect 1146 2978 1374 2981
rect 1394 2978 1430 2981
rect 1522 2978 1709 2981
rect 2578 2978 2662 2981
rect 3034 2978 3326 2981
rect 3650 2978 3869 2981
rect 3874 2978 4454 2981
rect 4462 2972 4465 2978
rect 778 2968 1942 2971
rect 2442 2968 3614 2971
rect 3618 2968 4078 2971
rect 4474 2968 4590 2971
rect 922 2958 1310 2961
rect 1322 2958 1510 2961
rect 1674 2958 2646 2961
rect 3714 2958 4462 2961
rect 4466 2958 4598 2961
rect 4602 2958 4614 2961
rect 5118 2952 5121 2958
rect 202 2948 694 2951
rect 866 2948 873 2951
rect 798 2942 801 2947
rect 870 2942 873 2948
rect 1306 2948 1438 2951
rect 1038 2942 1041 2948
rect 1906 2948 2222 2951
rect 2234 2948 2886 2951
rect 2978 2948 3549 2951
rect 3554 2948 3606 2951
rect 3634 2948 3718 2951
rect 3754 2948 4886 2951
rect 1130 2938 1310 2941
rect 1354 2938 2006 2941
rect 2042 2938 2534 2941
rect 2634 2938 2653 2941
rect 2666 2938 3638 2941
rect 3666 2938 4126 2941
rect 4338 2938 4630 2941
rect 970 2928 1238 2931
rect 1314 2928 1501 2931
rect 1514 2928 1878 2931
rect 1882 2928 1885 2931
rect 1954 2928 2398 2931
rect 2650 2928 3110 2931
rect 3866 2928 4073 2931
rect 1522 2918 1901 2921
rect 1182 2912 1185 2918
rect 1970 2918 2174 2921
rect 2178 2918 2606 2921
rect 2626 2918 4038 2921
rect 4070 2921 4073 2928
rect 4178 2928 4182 2931
rect 4070 2918 4093 2921
rect 5022 2912 5025 2918
rect 1290 2908 1718 2911
rect 1914 2908 2046 2911
rect 2130 2908 2878 2911
rect 3170 2908 3654 2911
rect 1054 2903 1057 2907
rect 1053 2902 1058 2903
rect 1063 2902 1064 2907
rect 2078 2903 2081 2907
rect 2077 2902 2082 2903
rect 2087 2902 2088 2907
rect 3102 2903 3105 2907
rect 3101 2902 3106 2903
rect 3111 2902 3112 2907
rect 3966 2902 3969 2908
rect 4118 2903 4121 2907
rect 4117 2902 4122 2903
rect 4127 2902 4128 2907
rect 1186 2898 1526 2901
rect 1626 2898 1645 2901
rect 1030 2891 1033 2898
rect 2178 2898 2198 2901
rect 2514 2898 2929 2901
rect 3586 2898 3790 2901
rect 2318 2892 2321 2898
rect 834 2888 1033 2891
rect 1090 2888 1150 2891
rect 1314 2888 1630 2891
rect 2058 2888 2126 2891
rect 2402 2888 2918 2891
rect 2926 2891 2929 2898
rect 4466 2898 4686 2901
rect 2926 2888 3405 2891
rect 3778 2888 3782 2891
rect 4002 2888 4166 2891
rect 4186 2888 4301 2891
rect 4306 2888 4902 2891
rect 5034 2888 5069 2891
rect 1026 2878 1373 2881
rect 1650 2878 1830 2881
rect 2162 2878 2534 2881
rect 3578 2878 3837 2881
rect 3858 2878 4230 2881
rect 2542 2872 2545 2877
rect 4622 2872 4625 2877
rect 578 2868 758 2871
rect 1010 2868 1021 2871
rect 1538 2868 2046 2871
rect 2562 2868 2662 2871
rect 3410 2868 3933 2871
rect 1218 2858 2222 2861
rect 2338 2858 2621 2861
rect 2802 2858 3102 2861
rect 3106 2858 3526 2861
rect 3530 2858 3790 2861
rect 3850 2858 4174 2861
rect 4194 2858 4406 2861
rect 4554 2858 4750 2861
rect 410 2848 790 2851
rect 938 2848 1662 2851
rect 2050 2848 2125 2851
rect 2314 2848 2630 2851
rect 3018 2848 3110 2851
rect 3338 2848 3750 2851
rect 3770 2848 4182 2851
rect 4194 2848 4350 2851
rect 1018 2838 1417 2841
rect 562 2828 1006 2831
rect 1414 2831 1417 2838
rect 1442 2838 1462 2841
rect 1514 2838 1606 2841
rect 1634 2838 2982 2841
rect 3050 2838 3158 2841
rect 3602 2838 3661 2841
rect 3722 2838 4526 2841
rect 1414 2828 1974 2831
rect 2106 2828 2822 2831
rect 3570 2828 3774 2831
rect 4378 2828 4430 2831
rect 786 2818 1038 2821
rect 1498 2818 1854 2821
rect 1978 2818 2454 2821
rect 3562 2818 4353 2821
rect 2510 2812 2513 2818
rect 4350 2812 4353 2818
rect 1442 2808 1550 2811
rect 1634 2808 1806 2811
rect 2018 2808 2478 2811
rect 2746 2808 3206 2811
rect 3754 2808 4334 2811
rect 4354 2808 4381 2811
rect 542 2803 545 2807
rect 541 2802 546 2803
rect 551 2802 552 2807
rect 1566 2803 1569 2807
rect 1565 2802 1570 2803
rect 1575 2802 1576 2807
rect 2590 2803 2593 2807
rect 2589 2802 2594 2803
rect 2599 2802 2600 2807
rect 3614 2803 3617 2807
rect 3613 2802 3618 2803
rect 3623 2802 3624 2807
rect 4638 2803 4641 2807
rect 4637 2802 4642 2803
rect 4647 2802 4648 2807
rect 1586 2798 1725 2801
rect 1730 2798 2118 2801
rect 2370 2798 2430 2801
rect 2626 2798 3062 2801
rect 3634 2798 3806 2801
rect 1426 2788 2086 2791
rect 2834 2788 3126 2791
rect 3618 2788 3766 2791
rect 3786 2788 4525 2791
rect 4650 2788 4662 2791
rect 5082 2788 5085 2791
rect 418 2778 653 2781
rect 658 2778 822 2781
rect 826 2778 1694 2781
rect 1730 2778 2110 2781
rect 2114 2778 2189 2781
rect 2194 2778 2902 2781
rect 2906 2778 3449 2781
rect 1346 2768 1774 2771
rect 1922 2768 1934 2771
rect 1990 2768 2198 2771
rect 2474 2768 3038 2771
rect 3446 2771 3449 2778
rect 3938 2778 5022 2781
rect 3446 2768 3822 2771
rect 3826 2768 3926 2771
rect 4138 2768 4141 2771
rect 314 2758 374 2761
rect 378 2758 510 2761
rect 514 2758 1454 2761
rect 1990 2761 1993 2768
rect 1626 2758 1993 2761
rect 2002 2758 3005 2761
rect 3602 2758 3702 2761
rect 3866 2758 3901 2761
rect 4530 2758 4894 2761
rect 4898 2758 5190 2761
rect 682 2748 701 2751
rect 746 2748 1629 2751
rect 1730 2748 1741 2751
rect 1754 2748 2246 2751
rect 2386 2748 3350 2751
rect 3538 2748 3885 2751
rect 1706 2738 1966 2741
rect 1970 2738 1981 2741
rect 2154 2738 2358 2741
rect 2562 2738 3693 2741
rect 3698 2738 3926 2741
rect 4234 2738 4438 2741
rect 954 2728 1750 2731
rect 1754 2728 1942 2731
rect 2098 2728 3174 2731
rect 3178 2728 3454 2731
rect 3458 2728 3742 2731
rect 3882 2728 3974 2731
rect 4082 2728 4462 2731
rect 1906 2718 2654 2721
rect 2658 2718 2718 2721
rect 2754 2718 2854 2721
rect 2858 2718 3629 2721
rect 3690 2718 3806 2721
rect 4058 2718 4446 2721
rect 1426 2708 1533 2711
rect 1650 2708 1805 2711
rect 2098 2708 2102 2711
rect 2250 2708 2702 2711
rect 2838 2708 2846 2711
rect 2850 2708 3054 2711
rect 3122 2708 3726 2711
rect 1054 2703 1057 2707
rect 1053 2702 1058 2703
rect 1063 2702 1064 2707
rect 2078 2703 2081 2707
rect 2077 2702 2082 2703
rect 2087 2702 2088 2707
rect 3102 2703 3105 2707
rect 3101 2702 3106 2703
rect 3111 2702 3112 2707
rect 4118 2703 4121 2707
rect 4117 2702 4122 2703
rect 4127 2702 4128 2707
rect 1658 2698 1902 2701
rect 2162 2698 2166 2701
rect 2506 2698 3070 2701
rect 3210 2698 3262 2701
rect 3698 2698 4046 2701
rect 4050 2698 4062 2701
rect 370 2688 574 2691
rect 1034 2688 1414 2691
rect 2058 2688 2637 2691
rect 2642 2688 2702 2691
rect 3074 2688 4014 2691
rect 4018 2688 4397 2691
rect 218 2678 686 2681
rect 842 2678 845 2681
rect 898 2678 998 2681
rect 1298 2678 1302 2681
rect 1402 2678 1854 2681
rect 1906 2678 1974 2681
rect 1994 2678 2381 2681
rect 2490 2678 2493 2681
rect 2514 2678 2913 2681
rect 3082 2678 3118 2681
rect 3354 2678 3686 2681
rect 3922 2678 4206 2681
rect 442 2668 758 2671
rect 762 2668 1182 2671
rect 1370 2668 1646 2671
rect 2050 2668 2205 2671
rect 2274 2668 2454 2671
rect 2850 2668 2902 2671
rect 2910 2671 2913 2678
rect 2910 2668 4014 2671
rect 5182 2662 5185 2668
rect 586 2658 838 2661
rect 1250 2658 1510 2661
rect 1538 2658 1581 2661
rect 1874 2658 1997 2661
rect 2090 2658 2150 2661
rect 2402 2658 2870 2661
rect 2874 2658 3582 2661
rect 4762 2658 5142 2661
rect 1002 2648 1502 2651
rect 1514 2648 2694 2651
rect 2706 2648 3846 2651
rect 3986 2648 4150 2651
rect 5114 2648 5182 2651
rect 650 2638 998 2641
rect 1226 2638 1366 2641
rect 1482 2638 1485 2641
rect 1698 2638 2542 2641
rect 2626 2638 3085 2641
rect 3266 2638 3926 2641
rect 5050 2638 5166 2641
rect 1662 2632 1665 2637
rect 698 2628 1254 2631
rect 1490 2628 1630 2631
rect 1746 2628 1750 2631
rect 1754 2628 2278 2631
rect 2298 2628 2301 2631
rect 2818 2628 4054 2631
rect 5106 2628 5110 2631
rect 330 2618 934 2621
rect 1570 2618 1661 2621
rect 1874 2618 1949 2621
rect 2066 2618 2142 2621
rect 2258 2618 2558 2621
rect 2610 2618 3126 2621
rect 3138 2618 3630 2621
rect 602 2608 1550 2611
rect 1594 2608 1677 2611
rect 1722 2608 1798 2611
rect 2154 2608 2334 2611
rect 2618 2608 2710 2611
rect 3090 2608 3373 2611
rect 542 2603 545 2607
rect 541 2602 546 2603
rect 551 2602 552 2607
rect 1566 2603 1569 2607
rect 1565 2602 1570 2603
rect 1575 2602 1576 2607
rect 2590 2603 2593 2607
rect 2589 2602 2594 2603
rect 2599 2602 2600 2607
rect 3614 2603 3617 2607
rect 3613 2602 3618 2603
rect 3623 2602 3624 2607
rect 4638 2603 4641 2607
rect 4637 2602 4642 2603
rect 4647 2602 4648 2607
rect 1162 2598 1206 2601
rect 1210 2598 1430 2601
rect 1918 2598 2198 2601
rect 2382 2598 2518 2601
rect 2714 2598 3230 2601
rect 1418 2588 1526 2591
rect 1918 2591 1921 2598
rect 1650 2588 1921 2591
rect 2382 2591 2385 2598
rect 2050 2588 2385 2591
rect 2478 2588 3310 2591
rect 786 2578 822 2581
rect 1154 2578 1710 2581
rect 1834 2578 1981 2581
rect 494 2572 497 2577
rect 574 2571 577 2578
rect 2018 2578 2045 2581
rect 2478 2581 2481 2588
rect 3842 2588 4078 2591
rect 4370 2588 4445 2591
rect 2266 2578 2481 2581
rect 2730 2578 2758 2581
rect 2826 2578 3134 2581
rect 574 2568 785 2571
rect 1290 2568 1318 2571
rect 1546 2568 1934 2571
rect 1954 2568 2086 2571
rect 2090 2568 2398 2571
rect 2850 2568 3133 2571
rect 782 2562 785 2568
rect 3218 2568 3469 2571
rect 3474 2568 3958 2571
rect 4394 2568 4622 2571
rect 1250 2558 1694 2561
rect 18 2548 414 2551
rect 1158 2551 1161 2558
rect 1954 2558 1958 2561
rect 2050 2558 3350 2561
rect 3914 2558 4278 2561
rect 4390 2561 4393 2568
rect 5106 2568 5126 2571
rect 4282 2558 4393 2561
rect 4690 2558 4766 2561
rect 5126 2558 5133 2561
rect 5126 2552 5129 2558
rect 1154 2548 1161 2551
rect 1210 2548 1213 2551
rect 1234 2548 1398 2551
rect 1450 2548 1686 2551
rect 1826 2548 2246 2551
rect 2322 2548 2702 2551
rect 2986 2548 3254 2551
rect 3338 2548 3382 2551
rect 3578 2548 3622 2551
rect 4526 2548 4790 2551
rect 4526 2542 4529 2548
rect 1322 2538 1526 2541
rect 1802 2538 1821 2541
rect 1954 2538 2070 2541
rect 2242 2538 2278 2541
rect 2402 2538 2638 2541
rect 2850 2538 3614 2541
rect 4162 2538 4470 2541
rect 5010 2538 5118 2541
rect 578 2528 846 2531
rect 930 2528 1590 2531
rect 1594 2528 2542 2531
rect 2642 2528 2950 2531
rect 3458 2528 3462 2531
rect 3522 2528 3806 2531
rect 3866 2528 4214 2531
rect 4218 2528 4494 2531
rect 10 2518 1654 2521
rect 1890 2518 1966 2521
rect 2018 2518 2109 2521
rect 1234 2508 1693 2511
rect 1750 2511 1753 2518
rect 2146 2518 2150 2521
rect 2234 2518 2345 2521
rect 2342 2512 2345 2518
rect 2354 2518 2422 2521
rect 2650 2518 3006 2521
rect 3146 2518 3374 2521
rect 4130 2518 4654 2521
rect 1714 2508 1753 2511
rect 1810 2508 1958 2511
rect 2466 2508 2494 2511
rect 3122 2508 3382 2511
rect 3466 2508 3934 2511
rect 1054 2503 1057 2507
rect 1053 2502 1058 2503
rect 1063 2502 1064 2507
rect 2078 2503 2081 2507
rect 2077 2502 2082 2503
rect 2087 2502 2088 2507
rect 634 2498 806 2501
rect 1074 2498 1270 2501
rect 1362 2498 1374 2501
rect 1890 2498 2045 2501
rect 2186 2498 2189 2501
rect 2202 2498 2333 2501
rect 2338 2498 2638 2501
rect 2934 2501 2937 2508
rect 3102 2503 3105 2507
rect 3101 2502 3106 2503
rect 3111 2502 3112 2507
rect 2746 2498 2937 2501
rect 122 2488 918 2491
rect 1018 2488 1230 2491
rect 2002 2488 2406 2491
rect 2610 2488 2630 2491
rect 2706 2488 2742 2491
rect 3006 2491 3009 2498
rect 3122 2498 3966 2501
rect 4102 2501 4105 2508
rect 4118 2503 4121 2507
rect 4117 2502 4122 2503
rect 4127 2502 4128 2507
rect 4082 2498 4105 2501
rect 3006 2488 3217 2491
rect 3434 2488 3910 2491
rect 3214 2482 3217 2488
rect 4082 2488 4430 2491
rect 546 2478 702 2481
rect 1018 2478 1030 2481
rect 1490 2478 1549 2481
rect 1810 2478 1830 2481
rect 2010 2478 2173 2481
rect 1934 2472 1937 2478
rect 2426 2478 2814 2481
rect 2890 2478 3142 2481
rect 3626 2478 3702 2481
rect 3954 2478 4205 2481
rect 1122 2468 1326 2471
rect 1754 2468 1926 2471
rect 354 2458 590 2461
rect 806 2461 809 2468
rect 2002 2468 2238 2471
rect 2322 2468 2654 2471
rect 2674 2468 2702 2471
rect 3026 2468 3117 2471
rect 3530 2468 3718 2471
rect 3810 2468 4174 2471
rect 4358 2471 4361 2478
rect 4178 2468 4361 2471
rect 4442 2468 4742 2471
rect 4858 2468 5134 2471
rect 806 2458 1174 2461
rect 1178 2458 1358 2461
rect 1394 2458 1462 2461
rect 1586 2458 1886 2461
rect 1898 2458 1953 2461
rect 590 2452 593 2458
rect 874 2448 1533 2451
rect 1538 2448 1549 2451
rect 1586 2448 1597 2451
rect 1770 2448 1942 2451
rect 1950 2451 1953 2458
rect 1986 2458 2174 2461
rect 2178 2458 2390 2461
rect 2402 2458 2462 2461
rect 2554 2458 2822 2461
rect 2974 2458 3006 2461
rect 3010 2458 3150 2461
rect 3194 2458 3790 2461
rect 2974 2451 2977 2458
rect 1950 2448 2977 2451
rect 3010 2448 3302 2451
rect 3306 2448 3470 2451
rect 3474 2448 3629 2451
rect 3862 2451 3865 2458
rect 3706 2448 3865 2451
rect 3950 2451 3953 2458
rect 3938 2448 3953 2451
rect 4194 2448 4382 2451
rect 18 2438 1254 2441
rect 1282 2438 1350 2441
rect 1458 2438 1597 2441
rect 1610 2438 1613 2441
rect 1706 2438 1734 2441
rect 1738 2438 1894 2441
rect 1906 2438 1910 2441
rect 1930 2438 2006 2441
rect 2050 2438 2478 2441
rect 2770 2438 2894 2441
rect 2898 2438 3117 2441
rect 3362 2438 3406 2441
rect 3418 2438 3974 2441
rect 4370 2438 4382 2441
rect 834 2428 1517 2431
rect 1538 2428 1838 2431
rect 1850 2428 1997 2431
rect 2050 2428 2798 2431
rect 2842 2428 3118 2431
rect 3130 2428 3422 2431
rect 3474 2428 3478 2431
rect 3570 2428 3766 2431
rect 3986 2428 4574 2431
rect 5138 2428 5149 2431
rect 666 2418 918 2421
rect 1114 2418 1214 2421
rect 1322 2418 1686 2421
rect 1230 2412 1233 2418
rect 1906 2418 1910 2421
rect 2066 2418 3342 2421
rect 3354 2418 3446 2421
rect 3618 2418 3990 2421
rect 5154 2418 5158 2421
rect 618 2408 894 2411
rect 1314 2408 1430 2411
rect 1610 2408 1902 2411
rect 2338 2408 2374 2411
rect 2754 2408 3134 2411
rect 3186 2408 3565 2411
rect 542 2403 545 2407
rect 541 2402 546 2403
rect 551 2402 552 2407
rect 1566 2403 1569 2407
rect 1565 2402 1570 2403
rect 1575 2402 1576 2407
rect 2590 2403 2593 2407
rect 2589 2402 2594 2403
rect 2599 2402 2600 2407
rect 3614 2403 3617 2407
rect 3613 2402 3618 2403
rect 3623 2402 3624 2407
rect 4638 2403 4641 2407
rect 4637 2402 4642 2403
rect 4647 2402 4648 2407
rect 1178 2398 1533 2401
rect 1602 2398 1654 2401
rect 1794 2398 1966 2401
rect 1974 2398 2166 2401
rect 2178 2398 2406 2401
rect 490 2388 622 2391
rect 898 2388 1318 2391
rect 1426 2388 1430 2391
rect 1434 2388 1670 2391
rect 1730 2388 1734 2391
rect 1750 2391 1753 2398
rect 1974 2391 1977 2398
rect 2914 2398 3206 2401
rect 4434 2398 4478 2401
rect 1750 2388 1977 2391
rect 2058 2388 2334 2391
rect 2378 2388 2381 2391
rect 2946 2388 3158 2391
rect 3306 2388 3438 2391
rect 3490 2388 3502 2391
rect 4578 2388 4654 2391
rect 946 2378 1158 2381
rect 1378 2378 1990 2381
rect 2090 2378 2093 2381
rect 2130 2378 2141 2381
rect 2146 2378 2230 2381
rect 2946 2378 2958 2381
rect 3122 2378 3798 2381
rect 4610 2378 5094 2381
rect 522 2368 1278 2371
rect 1602 2368 1606 2371
rect 1658 2368 2493 2371
rect 2586 2368 2702 2371
rect 2738 2368 2998 2371
rect 3114 2368 3305 2371
rect 3314 2368 3494 2371
rect 1226 2358 1246 2361
rect 1466 2358 2046 2361
rect 2250 2358 2414 2361
rect 2506 2358 2526 2361
rect 2698 2358 3254 2361
rect 3302 2361 3305 2368
rect 3602 2368 3622 2371
rect 3754 2368 3773 2371
rect 3810 2368 3902 2371
rect 3302 2358 3382 2361
rect 3806 2361 3809 2368
rect 4350 2362 4353 2368
rect 3386 2358 3809 2361
rect 3834 2358 3846 2361
rect 4546 2358 5094 2361
rect 18 2348 1230 2351
rect 1266 2348 1437 2351
rect 1522 2348 1710 2351
rect 1914 2348 2006 2351
rect 2050 2348 2198 2351
rect 2266 2348 2509 2351
rect 2514 2348 2630 2351
rect 2674 2348 2822 2351
rect 2970 2348 3165 2351
rect 3314 2348 3341 2351
rect 3426 2348 3558 2351
rect 3570 2348 3814 2351
rect 4178 2348 4350 2351
rect 1298 2338 1357 2341
rect 1506 2338 3526 2341
rect 3570 2338 3694 2341
rect 3834 2338 3870 2341
rect 3874 2338 4246 2341
rect 4474 2338 5102 2341
rect 18 2328 814 2331
rect 1266 2328 1409 2331
rect 1406 2322 1409 2328
rect 1458 2328 1725 2331
rect 1730 2328 2102 2331
rect 2210 2328 2294 2331
rect 2314 2328 2669 2331
rect 2682 2328 2918 2331
rect 2994 2328 4070 2331
rect 98 2318 1401 2321
rect 1498 2318 1750 2321
rect 1826 2318 1918 2321
rect 1954 2318 2337 2321
rect 3066 2318 3518 2321
rect 4358 2318 4702 2321
rect 1194 2308 1389 2311
rect 1398 2311 1401 2318
rect 2334 2312 2337 2318
rect 4358 2312 4361 2318
rect 1398 2308 1406 2311
rect 1490 2308 2054 2311
rect 2098 2308 2238 2311
rect 3298 2308 3318 2311
rect 3442 2308 3446 2311
rect 3522 2308 3581 2311
rect 4390 2308 4646 2311
rect 1054 2303 1057 2307
rect 1053 2302 1058 2303
rect 1063 2302 1064 2307
rect 2078 2303 2081 2307
rect 2077 2302 2082 2303
rect 2087 2302 2088 2307
rect 3102 2303 3105 2307
rect 3101 2302 3106 2303
rect 3111 2302 3112 2307
rect 4118 2303 4121 2307
rect 4117 2302 4122 2303
rect 4127 2302 4128 2307
rect 4390 2302 4393 2308
rect 4962 2308 5062 2311
rect 1202 2298 1806 2301
rect 1890 2298 1998 2301
rect 2146 2298 2157 2301
rect 2162 2298 2957 2301
rect 2962 2298 2966 2301
rect 3234 2298 3238 2301
rect 3482 2298 3758 2301
rect 1258 2288 1534 2291
rect 1618 2288 1878 2291
rect 1962 2288 2206 2291
rect 2338 2288 3566 2291
rect 3570 2288 4413 2291
rect 4418 2288 4446 2291
rect 386 2278 654 2281
rect 1218 2278 1510 2281
rect 1674 2278 1894 2281
rect 1914 2278 1966 2281
rect 2154 2278 2157 2281
rect 2194 2278 2238 2281
rect 2274 2278 2990 2281
rect 3618 2278 4638 2281
rect 4830 2272 4833 2278
rect 5138 2278 5142 2281
rect 482 2268 1246 2271
rect 1258 2268 1622 2271
rect 1698 2268 2093 2271
rect 2114 2268 2118 2271
rect 2258 2268 2878 2271
rect 3122 2268 3774 2271
rect 4122 2268 4541 2271
rect 4546 2268 4750 2271
rect 274 2258 945 2261
rect 1610 2258 1645 2261
rect 942 2252 945 2258
rect 1698 2258 2150 2261
rect 2418 2258 2813 2261
rect 2954 2258 3630 2261
rect 3786 2258 4182 2261
rect 4186 2258 4253 2261
rect 4286 2252 4289 2258
rect 5090 2258 5150 2261
rect 1410 2248 1462 2251
rect 1826 2248 1897 2251
rect 1138 2238 1373 2241
rect 1378 2238 1702 2241
rect 1894 2241 1897 2248
rect 1922 2248 1981 2251
rect 1986 2248 2118 2251
rect 2130 2248 2909 2251
rect 3722 2248 3854 2251
rect 3874 2248 3974 2251
rect 4418 2248 4573 2251
rect 1894 2238 1998 2241
rect 2034 2238 2462 2241
rect 2578 2238 3062 2241
rect 3066 2238 3358 2241
rect 3362 2238 3670 2241
rect 3738 2238 3773 2241
rect 3810 2238 4237 2241
rect 4242 2238 4702 2241
rect 2558 2232 2561 2237
rect 898 2228 909 2231
rect 1778 2228 1830 2231
rect 1994 2228 2125 2231
rect 2322 2228 2334 2231
rect 2634 2228 2966 2231
rect 3026 2228 3422 2231
rect 3442 2228 3574 2231
rect 3602 2228 4222 2231
rect 4226 2228 4254 2231
rect 4394 2228 4566 2231
rect 266 2218 470 2221
rect 474 2218 1334 2221
rect 1338 2218 1582 2221
rect 1658 2218 1838 2221
rect 2074 2218 2270 2221
rect 2490 2218 3110 2221
rect 3218 2218 3414 2221
rect 3466 2218 3710 2221
rect 3874 2218 4038 2221
rect 4090 2218 4470 2221
rect 962 2208 1006 2211
rect 1586 2208 1838 2211
rect 1890 2208 1990 2211
rect 2066 2208 2206 2211
rect 2698 2208 2958 2211
rect 2970 2208 3297 2211
rect 3306 2208 3309 2211
rect 542 2203 545 2207
rect 541 2202 546 2203
rect 551 2202 552 2207
rect 1566 2203 1569 2207
rect 1565 2202 1570 2203
rect 1575 2202 1576 2207
rect 2590 2203 2593 2207
rect 2589 2202 2594 2203
rect 2599 2202 2600 2207
rect 634 2198 1502 2201
rect 1842 2198 1950 2201
rect 2050 2198 2166 2201
rect 2242 2198 2446 2201
rect 2818 2198 3286 2201
rect 3294 2201 3297 2208
rect 3746 2208 4006 2211
rect 3614 2203 3617 2207
rect 3613 2202 3618 2203
rect 3623 2202 3624 2207
rect 4638 2203 4641 2207
rect 4637 2202 4642 2203
rect 4647 2202 4648 2207
rect 3294 2198 3510 2201
rect 3634 2198 4398 2201
rect 834 2188 854 2191
rect 1362 2188 1581 2191
rect 1882 2188 1934 2191
rect 2066 2188 2253 2191
rect 2322 2188 3150 2191
rect 3562 2188 3750 2191
rect 3762 2188 4206 2191
rect 594 2178 1629 2181
rect 1642 2178 1822 2181
rect 1962 2178 2350 2181
rect 2482 2178 2966 2181
rect 3002 2178 3037 2181
rect 3554 2178 3742 2181
rect 3746 2178 3981 2181
rect 3994 2178 4486 2181
rect 842 2168 1174 2171
rect 1898 2168 1901 2171
rect 1914 2168 2102 2171
rect 2418 2168 3022 2171
rect 3858 2168 4366 2171
rect 642 2158 654 2161
rect 930 2158 950 2161
rect 962 2158 1645 2161
rect 1930 2158 2118 2161
rect 2150 2161 2153 2168
rect 2150 2158 2269 2161
rect 2818 2158 3149 2161
rect 3290 2158 3689 2161
rect 3698 2158 4038 2161
rect 4586 2158 4749 2161
rect 1790 2152 1793 2157
rect 386 2148 878 2151
rect 1074 2148 1390 2151
rect 1898 2148 2510 2151
rect 2514 2148 2534 2151
rect 338 2138 694 2141
rect 910 2141 913 2148
rect 2546 2148 3054 2151
rect 3058 2148 3654 2151
rect 3686 2151 3689 2158
rect 4794 2158 4905 2161
rect 4902 2152 4905 2158
rect 3686 2148 4342 2151
rect 4346 2148 4525 2151
rect 4530 2148 4678 2151
rect 738 2138 913 2141
rect 962 2138 1118 2141
rect 1218 2138 1318 2141
rect 1474 2138 2317 2141
rect 2434 2138 2765 2141
rect 2850 2138 3078 2141
rect 3354 2138 3422 2141
rect 3538 2138 3805 2141
rect 4346 2138 4589 2141
rect 98 2128 1558 2131
rect 1778 2128 1889 2131
rect 1962 2128 2710 2131
rect 2930 2128 3478 2131
rect 3602 2128 3998 2131
rect 1886 2122 1889 2128
rect 4218 2128 4382 2131
rect 4554 2128 4910 2131
rect 4094 2122 4097 2127
rect 1034 2118 1398 2121
rect 1402 2118 1709 2121
rect 1754 2118 1773 2121
rect 1890 2118 2982 2121
rect 3058 2118 3238 2121
rect 3410 2118 3454 2121
rect 3738 2118 4054 2121
rect 4370 2118 4557 2121
rect 4562 2118 4766 2121
rect 690 2108 870 2111
rect 1330 2108 1694 2111
rect 1730 2108 1950 2111
rect 2034 2108 2045 2111
rect 2274 2108 2998 2111
rect 3250 2108 3481 2111
rect 4770 2108 5014 2111
rect 1054 2103 1057 2107
rect 1053 2102 1058 2103
rect 1063 2102 1064 2107
rect 2078 2103 2081 2107
rect 2077 2102 2082 2103
rect 2087 2102 2088 2107
rect 3102 2103 3105 2107
rect 3101 2102 3106 2103
rect 3111 2102 3112 2107
rect 1238 2098 1702 2101
rect 82 2088 166 2091
rect 1238 2091 1241 2098
rect 1714 2098 1958 2101
rect 2314 2098 3038 2101
rect 3130 2098 3286 2101
rect 3478 2101 3481 2108
rect 4118 2103 4121 2107
rect 4117 2102 4122 2103
rect 4127 2102 4128 2107
rect 3478 2098 3862 2101
rect 4170 2098 4902 2101
rect 986 2088 1241 2091
rect 1338 2088 1341 2091
rect 1666 2088 1805 2091
rect 1970 2088 2182 2091
rect 2302 2088 2398 2091
rect 2586 2088 2797 2091
rect 1042 2078 1046 2081
rect 1194 2078 1502 2081
rect 1586 2078 1630 2081
rect 1650 2078 1801 2081
rect 1850 2078 2046 2081
rect 2302 2081 2305 2088
rect 3018 2088 3942 2091
rect 4722 2088 5006 2091
rect 2082 2078 2305 2081
rect 2314 2078 2670 2081
rect 2682 2078 3566 2081
rect 626 2068 1270 2071
rect 1290 2068 1581 2071
rect 1798 2071 1801 2078
rect 3634 2078 3902 2081
rect 3906 2078 4093 2081
rect 4474 2078 4477 2081
rect 4594 2078 4998 2081
rect 5066 2078 5085 2081
rect 4510 2072 4513 2077
rect 1698 2068 1793 2071
rect 1798 2068 2142 2071
rect 2258 2068 2333 2071
rect 1098 2058 1121 2061
rect 1554 2058 1766 2061
rect 1790 2061 1793 2068
rect 3254 2068 3414 2071
rect 3434 2068 3437 2071
rect 1790 2058 2246 2061
rect 2498 2058 2790 2061
rect 1118 2052 1121 2058
rect 3254 2061 3257 2068
rect 2802 2058 3257 2061
rect 3430 2061 3433 2068
rect 3458 2068 3510 2071
rect 3666 2068 4054 2071
rect 4058 2068 4294 2071
rect 4666 2068 4669 2071
rect 4946 2068 5070 2071
rect 3266 2058 3433 2061
rect 3586 2058 3942 2061
rect 4138 2058 4157 2061
rect 4418 2058 4998 2061
rect 5190 2061 5193 2068
rect 5002 2058 5193 2061
rect 386 2048 478 2051
rect 1434 2048 3326 2051
rect 3330 2048 3886 2051
rect 3898 2048 3942 2051
rect 4178 2048 4189 2051
rect 658 2038 662 2041
rect 682 2038 1486 2041
rect 1554 2038 1710 2041
rect 1746 2038 1853 2041
rect 2050 2038 2105 2041
rect 690 2028 1069 2031
rect 1114 2028 1566 2031
rect 1634 2028 1854 2031
rect 1858 2028 2014 2031
rect 2102 2031 2105 2038
rect 2114 2038 2118 2041
rect 3122 2038 3166 2041
rect 3210 2038 3709 2041
rect 3914 2038 3933 2041
rect 4034 2038 5134 2041
rect 5166 2032 5169 2037
rect 2102 2028 2518 2031
rect 3178 2028 3181 2031
rect 3474 2028 4118 2031
rect 4154 2028 4486 2031
rect 986 2018 1678 2021
rect 1698 2018 2206 2021
rect 2514 2018 2542 2021
rect 3090 2018 3790 2021
rect 4026 2018 4662 2021
rect 914 2008 1182 2011
rect 1610 2008 2045 2011
rect 2058 2008 2278 2011
rect 2618 2008 2726 2011
rect 2730 2008 3358 2011
rect 3538 2008 3549 2011
rect 3578 2008 3581 2011
rect 3730 2008 3758 2011
rect 542 2003 545 2007
rect 541 2002 546 2003
rect 551 2002 552 2007
rect 1566 2003 1569 2007
rect 1565 2002 1570 2003
rect 1575 2002 1576 2007
rect 2590 2003 2593 2007
rect 2589 2002 2594 2003
rect 2599 2002 2600 2007
rect 3614 2003 3617 2007
rect 3613 2002 3618 2003
rect 3623 2002 3624 2007
rect 4638 2003 4641 2007
rect 4637 2002 4642 2003
rect 4647 2002 4648 2007
rect 746 1998 1494 2001
rect 1706 1998 2141 2001
rect 2674 1998 3342 2001
rect 3354 1998 3430 2001
rect 4114 1998 4574 2001
rect 1106 1988 1341 1991
rect 1490 1988 3726 1991
rect 4862 1982 4865 1987
rect 1146 1978 1149 1981
rect 1474 1978 2014 1981
rect 2074 1978 2414 1981
rect 2418 1978 3414 1981
rect 4018 1978 4094 1981
rect 4226 1978 4238 1981
rect 1074 1968 1278 1971
rect 1290 1968 1350 1971
rect 1442 1968 2086 1971
rect 2098 1968 2109 1971
rect 2490 1968 3206 1971
rect 3210 1968 4022 1971
rect 4234 1968 4646 1971
rect 618 1958 878 1961
rect 1506 1958 2310 1961
rect 3362 1958 3926 1961
rect 4418 1958 4430 1961
rect 298 1948 1134 1951
rect 1154 1948 1165 1951
rect 1346 1948 1830 1951
rect 2470 1948 2982 1951
rect 3306 1948 3382 1951
rect 2470 1942 2473 1948
rect 3426 1948 3430 1951
rect 3506 1948 3558 1951
rect 3858 1948 3869 1951
rect 4086 1951 4089 1958
rect 4026 1948 4089 1951
rect 4702 1951 4705 1958
rect 4378 1948 4705 1951
rect 946 1938 1161 1941
rect 862 1932 865 1937
rect 1158 1932 1161 1938
rect 1506 1938 1510 1941
rect 1610 1938 1774 1941
rect 1826 1938 2081 1941
rect 2330 1938 2333 1941
rect 1314 1928 1422 1931
rect 1970 1928 2070 1931
rect 2078 1931 2081 1938
rect 2498 1938 3894 1941
rect 3898 1938 4166 1941
rect 4178 1938 4190 1941
rect 4338 1938 4734 1941
rect 2078 1928 2150 1931
rect 2202 1928 2630 1931
rect 3010 1928 3182 1931
rect 3434 1928 4062 1931
rect 978 1918 1405 1921
rect 1418 1918 2749 1921
rect 2786 1918 2902 1921
rect 3154 1918 3309 1921
rect 3314 1918 3902 1921
rect 3906 1918 4670 1921
rect 4882 1918 4925 1921
rect 1538 1908 2062 1911
rect 2098 1908 2534 1911
rect 2546 1908 3053 1911
rect 3130 1908 3357 1911
rect 3522 1908 3597 1911
rect 3602 1908 3606 1911
rect 4034 1908 4061 1911
rect 1054 1903 1057 1907
rect 1053 1902 1058 1903
rect 1063 1902 1064 1907
rect 2078 1903 2081 1907
rect 2077 1902 2082 1903
rect 2087 1902 2088 1907
rect 3102 1903 3105 1907
rect 3101 1902 3106 1903
rect 3111 1902 3112 1907
rect 4118 1903 4121 1907
rect 4117 1902 4122 1903
rect 4127 1902 4128 1907
rect 650 1898 790 1901
rect 1410 1898 1838 1901
rect 1986 1898 2046 1901
rect 2098 1898 2413 1901
rect 2418 1898 2430 1901
rect 2434 1898 3078 1901
rect 3578 1898 4086 1901
rect 4350 1892 4353 1897
rect 394 1888 606 1891
rect 1090 1888 1785 1891
rect 1810 1888 1918 1891
rect 1922 1888 2230 1891
rect 2290 1888 2614 1891
rect 2618 1888 2806 1891
rect 1402 1878 1774 1881
rect 1782 1881 1785 1888
rect 3938 1888 4278 1891
rect 4298 1888 4301 1891
rect 4466 1888 4870 1891
rect 1782 1878 2390 1881
rect 2650 1878 2685 1881
rect 1082 1868 1165 1871
rect 1174 1871 1177 1878
rect 1230 1871 1233 1878
rect 2690 1878 3478 1881
rect 3634 1878 3757 1881
rect 3762 1878 3814 1881
rect 4010 1878 4654 1881
rect 4730 1878 4822 1881
rect 3486 1872 3489 1877
rect 1174 1868 1309 1871
rect 1402 1868 1518 1871
rect 1610 1868 1613 1871
rect 1666 1868 2189 1871
rect 2626 1868 3481 1871
rect 4122 1868 4301 1871
rect 994 1858 1293 1861
rect 1298 1858 1302 1861
rect 1618 1858 2134 1861
rect 2338 1858 2374 1861
rect 2706 1858 3190 1861
rect 3478 1861 3481 1868
rect 4306 1868 4382 1871
rect 4850 1868 4870 1871
rect 5018 1868 5021 1871
rect 3478 1858 3694 1861
rect 3978 1858 4454 1861
rect 4458 1858 4477 1861
rect 3470 1852 3473 1857
rect 1554 1848 1806 1851
rect 1842 1848 1894 1851
rect 1898 1848 2174 1851
rect 2202 1848 2358 1851
rect 2858 1848 3406 1851
rect 4170 1848 4198 1851
rect 4546 1848 4557 1851
rect 1010 1838 1318 1841
rect 1394 1838 1758 1841
rect 1994 1838 2013 1841
rect 2026 1838 2246 1841
rect 2730 1838 3933 1841
rect 4042 1838 4766 1841
rect 466 1828 1326 1831
rect 1514 1828 1734 1831
rect 1770 1828 2702 1831
rect 3650 1828 4749 1831
rect 4754 1828 4918 1831
rect 1170 1818 1534 1821
rect 1682 1818 2062 1821
rect 2362 1818 3446 1821
rect 3450 1818 3453 1821
rect 4178 1818 4374 1821
rect 1586 1808 1886 1811
rect 2130 1808 2429 1811
rect 3386 1808 3582 1811
rect 3778 1808 4550 1811
rect 542 1803 545 1807
rect 541 1802 546 1803
rect 551 1802 552 1807
rect 1566 1803 1569 1807
rect 1565 1802 1570 1803
rect 1575 1802 1576 1807
rect 2590 1803 2593 1807
rect 2589 1802 2594 1803
rect 2599 1802 2600 1807
rect 3614 1803 3617 1807
rect 3613 1802 3618 1803
rect 3623 1802 3624 1807
rect 4638 1803 4641 1807
rect 4637 1802 4642 1803
rect 4647 1802 4648 1807
rect 858 1798 1430 1801
rect 1474 1798 1478 1801
rect 1874 1798 2078 1801
rect 3762 1798 4574 1801
rect 242 1788 1241 1791
rect 1306 1788 2142 1791
rect 2874 1788 3158 1791
rect 4082 1788 4470 1791
rect 4474 1788 4846 1791
rect 1238 1781 1241 1788
rect 1238 1778 1750 1781
rect 1754 1778 3382 1781
rect 3394 1778 3678 1781
rect 3794 1778 3798 1781
rect 1362 1768 2238 1771
rect 2250 1768 3117 1771
rect 3474 1768 3550 1771
rect 3746 1768 4078 1771
rect 4818 1768 4974 1771
rect 1530 1758 1734 1761
rect 1762 1758 1782 1761
rect 1842 1758 2182 1761
rect 2858 1758 3085 1761
rect 3690 1758 3934 1761
rect 3994 1758 4254 1761
rect 4298 1758 4910 1761
rect 762 1748 1174 1751
rect 1202 1748 1214 1751
rect 1434 1748 1454 1751
rect 1498 1748 2070 1751
rect 2090 1748 2093 1751
rect 2154 1748 2541 1751
rect 2706 1748 3030 1751
rect 3406 1751 3409 1758
rect 3406 1748 3598 1751
rect 3834 1748 4302 1751
rect 4338 1748 4374 1751
rect 4434 1748 4438 1751
rect 1034 1738 1085 1741
rect 1122 1738 1478 1741
rect 1506 1738 1886 1741
rect 2042 1738 2190 1741
rect 2194 1738 2494 1741
rect 2498 1738 2838 1741
rect 2842 1738 3142 1741
rect 3818 1738 4222 1741
rect 4230 1738 4918 1741
rect 1106 1728 2430 1731
rect 2490 1728 3190 1731
rect 3194 1728 3277 1731
rect 4230 1731 4233 1738
rect 3506 1728 4233 1731
rect 4578 1728 4982 1731
rect 702 1722 705 1727
rect 1234 1718 1478 1721
rect 1650 1718 1814 1721
rect 1874 1718 2102 1721
rect 2162 1718 2182 1721
rect 2194 1718 2414 1721
rect 2770 1718 3070 1721
rect 3090 1718 3766 1721
rect 3970 1718 4870 1721
rect 5022 1712 5025 1718
rect 674 1708 718 1711
rect 1242 1708 1774 1711
rect 2122 1708 2942 1711
rect 3522 1708 3998 1711
rect 4410 1708 4614 1711
rect 4618 1708 4621 1711
rect 1054 1703 1057 1707
rect 1053 1702 1058 1703
rect 1063 1702 1064 1707
rect 2078 1703 2081 1707
rect 2077 1702 2082 1703
rect 2087 1702 2088 1707
rect 3102 1703 3105 1707
rect 3101 1702 3106 1703
rect 3111 1702 3112 1707
rect 4118 1703 4121 1707
rect 4117 1702 4122 1703
rect 4127 1702 4128 1707
rect 1186 1698 1270 1701
rect 1746 1698 1750 1701
rect 2194 1698 2397 1701
rect 3122 1698 3854 1701
rect 4450 1698 4461 1701
rect 4858 1698 4861 1701
rect 1282 1688 1854 1691
rect 1858 1688 2446 1691
rect 3306 1688 3414 1691
rect 3794 1688 3998 1691
rect 4082 1688 4230 1691
rect 782 1682 785 1687
rect 594 1678 782 1681
rect 954 1678 957 1681
rect 1162 1678 1542 1681
rect 2090 1678 2438 1681
rect 2442 1678 2758 1681
rect 2786 1678 3086 1681
rect 3098 1678 3822 1681
rect 3994 1678 3997 1681
rect 4450 1678 4582 1681
rect 4634 1678 4862 1681
rect 370 1668 574 1671
rect 770 1668 926 1671
rect 954 1668 1910 1671
rect 1914 1668 2361 1671
rect 2370 1668 2670 1671
rect 2674 1668 3382 1671
rect 3690 1668 3693 1671
rect 1450 1658 1822 1661
rect 1882 1658 2285 1661
rect 2358 1661 2361 1668
rect 4546 1668 4614 1671
rect 4618 1668 4670 1671
rect 2358 1658 2526 1661
rect 2578 1658 3278 1661
rect 3282 1658 3502 1661
rect 3842 1658 4374 1661
rect 4470 1661 4473 1668
rect 4402 1658 4473 1661
rect 674 1648 1246 1651
rect 1274 1648 1326 1651
rect 1330 1648 2830 1651
rect 2866 1648 3166 1651
rect 3170 1648 3198 1651
rect 3218 1648 4158 1651
rect 4338 1648 4502 1651
rect 674 1638 822 1641
rect 1754 1638 2134 1641
rect 1518 1632 1521 1638
rect 2210 1638 2221 1641
rect 2226 1638 2446 1641
rect 2450 1638 3134 1641
rect 3154 1638 3342 1641
rect 3570 1638 3774 1641
rect 4554 1638 4686 1641
rect 458 1628 1094 1631
rect 2178 1628 2326 1631
rect 2394 1628 2926 1631
rect 4078 1631 4081 1638
rect 2946 1628 4081 1631
rect 4190 1628 4718 1631
rect 4722 1628 4765 1631
rect 1806 1622 1809 1627
rect 410 1618 1670 1621
rect 1818 1618 1822 1621
rect 1826 1618 2286 1621
rect 2290 1618 2870 1621
rect 2898 1618 3318 1621
rect 4190 1621 4193 1628
rect 3602 1618 4193 1621
rect 2626 1608 3094 1611
rect 3330 1608 3334 1611
rect 3714 1608 3757 1611
rect 542 1603 545 1607
rect 541 1602 546 1603
rect 551 1602 552 1607
rect 1566 1603 1569 1607
rect 1565 1602 1570 1603
rect 1575 1602 1576 1607
rect 2590 1603 2593 1607
rect 2589 1602 2594 1603
rect 2599 1602 2600 1607
rect 3614 1603 3617 1607
rect 3613 1602 3618 1603
rect 3623 1602 3624 1607
rect 4638 1603 4641 1607
rect 4637 1602 4642 1603
rect 4647 1602 4648 1607
rect 1594 1598 1597 1601
rect 1938 1598 2166 1601
rect 2778 1598 3598 1601
rect 3762 1598 4038 1601
rect 4346 1598 4470 1601
rect 1026 1588 1086 1591
rect 1098 1588 1693 1591
rect 1890 1588 2262 1591
rect 2322 1588 2366 1591
rect 2370 1588 3470 1591
rect 3474 1588 4206 1591
rect 4610 1588 4710 1591
rect 850 1578 1374 1581
rect 1410 1578 1702 1581
rect 1706 1578 2486 1581
rect 2850 1578 3006 1581
rect 3650 1578 3670 1581
rect 3674 1578 4078 1581
rect 4106 1578 4350 1581
rect 1082 1568 1142 1571
rect 1178 1568 1886 1571
rect 1954 1568 2217 1571
rect 2282 1568 2701 1571
rect 1074 1558 1326 1561
rect 1578 1558 2094 1561
rect 2214 1561 2217 1568
rect 2738 1568 3622 1571
rect 3794 1568 3798 1571
rect 3858 1568 3878 1571
rect 4066 1568 4902 1571
rect 2214 1558 3630 1561
rect 4074 1558 5014 1561
rect 890 1548 958 1551
rect 962 1548 1486 1551
rect 1558 1551 1561 1558
rect 1558 1548 1598 1551
rect 1954 1548 1958 1551
rect 2206 1551 2209 1558
rect 2058 1548 2209 1551
rect 2306 1548 2462 1551
rect 3450 1548 3838 1551
rect 4282 1548 4398 1551
rect 730 1538 990 1541
rect 1218 1538 2237 1541
rect 2834 1538 2854 1541
rect 3218 1538 3549 1541
rect 3554 1538 3582 1541
rect 3586 1538 3894 1541
rect 418 1528 589 1531
rect 594 1528 1422 1531
rect 1722 1528 2278 1531
rect 2294 1528 2753 1531
rect 2762 1528 3038 1531
rect 3066 1528 3150 1531
rect 946 1518 1302 1521
rect 2294 1521 2297 1528
rect 1914 1518 2297 1521
rect 2750 1521 2753 1528
rect 3338 1528 3342 1531
rect 3354 1528 3590 1531
rect 3866 1528 4166 1531
rect 2750 1518 2894 1521
rect 2906 1518 3958 1521
rect 1770 1508 1942 1511
rect 2122 1508 2862 1511
rect 1054 1503 1057 1507
rect 1053 1502 1058 1503
rect 1063 1502 1064 1507
rect 1390 1501 1393 1508
rect 3778 1508 4062 1511
rect 2078 1503 2081 1507
rect 2077 1502 2082 1503
rect 2087 1502 2088 1507
rect 3102 1503 3105 1507
rect 3101 1502 3106 1503
rect 3111 1502 3112 1507
rect 4118 1503 4121 1507
rect 4117 1502 4122 1503
rect 4127 1502 4128 1507
rect 1390 1498 1678 1501
rect 1690 1498 1725 1501
rect 2778 1498 3054 1501
rect 3226 1498 3229 1501
rect 3242 1498 3805 1501
rect 3906 1498 3910 1501
rect 4186 1498 5054 1501
rect 5086 1492 5089 1497
rect 1362 1488 1373 1491
rect 1482 1488 1485 1491
rect 1506 1488 2158 1491
rect 2194 1488 2198 1491
rect 2202 1488 2621 1491
rect 2698 1488 3118 1491
rect 3186 1488 3214 1491
rect 4322 1488 4502 1491
rect 4658 1488 4742 1491
rect 1226 1478 1702 1481
rect 1978 1478 2061 1481
rect 766 1472 769 1478
rect 2290 1478 3293 1481
rect 3810 1478 4126 1481
rect 4362 1478 4430 1481
rect 4742 1481 4745 1488
rect 4738 1478 4745 1481
rect 226 1468 765 1471
rect 1178 1468 1181 1471
rect 1186 1468 1198 1471
rect 1346 1468 1422 1471
rect 1898 1468 1997 1471
rect 2002 1468 2190 1471
rect 2194 1468 2702 1471
rect 2810 1468 3005 1471
rect 3146 1468 3182 1471
rect 4258 1468 4366 1471
rect 1194 1458 2166 1461
rect 2194 1458 3078 1461
rect 3090 1458 3486 1461
rect 3490 1458 3878 1461
rect 386 1448 430 1451
rect 434 1448 486 1451
rect 490 1448 1230 1451
rect 1330 1448 1550 1451
rect 1570 1448 1782 1451
rect 3130 1448 3574 1451
rect 3578 1448 3677 1451
rect 3682 1448 3718 1451
rect 810 1438 813 1441
rect 826 1438 1166 1441
rect 1170 1438 1190 1441
rect 1202 1438 1470 1441
rect 1474 1438 1622 1441
rect 1634 1438 2125 1441
rect 2290 1438 3446 1441
rect 3818 1438 3821 1441
rect 386 1428 1214 1431
rect 1234 1428 2158 1431
rect 2250 1428 4726 1431
rect 298 1418 398 1421
rect 402 1418 598 1421
rect 602 1418 2302 1421
rect 2410 1418 3102 1421
rect 3114 1418 3469 1421
rect 3938 1418 4566 1421
rect 834 1408 845 1411
rect 954 1408 966 1411
rect 1138 1408 1422 1411
rect 1802 1408 2246 1411
rect 2922 1408 3430 1411
rect 542 1403 545 1407
rect 541 1402 546 1403
rect 551 1402 552 1407
rect 1566 1403 1569 1407
rect 1565 1402 1570 1403
rect 1575 1402 1576 1407
rect 2590 1403 2593 1407
rect 2589 1402 2594 1403
rect 2599 1402 2600 1407
rect 3614 1403 3617 1407
rect 3613 1402 3618 1403
rect 3623 1402 3624 1407
rect 4638 1403 4641 1407
rect 4637 1402 4642 1403
rect 4647 1402 4648 1407
rect 626 1398 1446 1401
rect 1642 1398 2086 1401
rect 2138 1398 2398 1401
rect 3090 1398 3454 1401
rect 506 1388 806 1391
rect 1650 1388 2574 1391
rect 3002 1388 3742 1391
rect 3746 1388 3949 1391
rect 1234 1378 1245 1381
rect 1394 1378 2558 1381
rect 2842 1378 3414 1381
rect 1154 1368 1198 1371
rect 1266 1368 1958 1371
rect 2954 1368 3565 1371
rect 4050 1368 4077 1371
rect 4138 1368 4141 1371
rect 642 1358 934 1361
rect 1138 1358 1230 1361
rect 1346 1358 1366 1361
rect 1370 1358 2022 1361
rect 2050 1358 3358 1361
rect 3362 1358 3597 1361
rect 3802 1358 3805 1361
rect 3874 1358 4390 1361
rect 578 1348 717 1351
rect 938 1348 1398 1351
rect 1562 1348 1613 1351
rect 1622 1348 1902 1351
rect 2314 1348 2393 1351
rect 3106 1348 3758 1351
rect 4290 1348 4550 1351
rect 634 1338 925 1341
rect 1622 1341 1625 1348
rect 930 1338 1625 1341
rect 2390 1342 2393 1348
rect 3330 1338 4518 1341
rect 882 1328 886 1331
rect 890 1328 1238 1331
rect 2026 1328 2542 1331
rect 2866 1328 2926 1331
rect 3626 1328 4054 1331
rect 362 1318 750 1321
rect 754 1318 1102 1321
rect 1250 1318 1342 1321
rect 1938 1318 3254 1321
rect 450 1308 1038 1311
rect 1234 1308 1350 1311
rect 2146 1308 2797 1311
rect 3170 1308 3814 1311
rect 3818 1308 3982 1311
rect 1054 1303 1057 1307
rect 1053 1302 1058 1303
rect 1063 1302 1064 1307
rect 2078 1303 2081 1307
rect 2077 1302 2082 1303
rect 2087 1302 2088 1307
rect 3102 1303 3105 1307
rect 3101 1302 3106 1303
rect 3111 1302 3112 1307
rect 4118 1303 4121 1307
rect 4117 1302 4122 1303
rect 4127 1302 4128 1307
rect 1386 1298 1942 1301
rect 3138 1298 3213 1301
rect 3218 1298 3246 1301
rect 3314 1298 3870 1301
rect 1170 1288 1198 1291
rect 1202 1288 2198 1291
rect 2274 1288 2697 1291
rect 1466 1278 2326 1281
rect 2586 1278 2637 1281
rect 2694 1281 2697 1288
rect 2706 1288 3998 1291
rect 2694 1278 3038 1281
rect 3058 1278 3950 1281
rect 4574 1272 4577 1277
rect 594 1268 598 1271
rect 1002 1268 1126 1271
rect 1882 1268 2070 1271
rect 2578 1268 3622 1271
rect 386 1258 782 1261
rect 1202 1258 1326 1261
rect 2086 1261 2089 1268
rect 2086 1258 2093 1261
rect 2162 1258 2638 1261
rect 2882 1258 3182 1261
rect 3258 1258 3518 1261
rect 3834 1258 4342 1261
rect 4678 1261 4681 1268
rect 4678 1258 5094 1261
rect 474 1248 590 1251
rect 594 1248 1406 1251
rect 1450 1248 1894 1251
rect 2946 1248 3286 1251
rect 3290 1248 3405 1251
rect 3530 1248 3878 1251
rect 5014 1248 5021 1251
rect 5014 1242 5017 1248
rect 1114 1238 1261 1241
rect 2514 1238 3110 1241
rect 3378 1238 3726 1241
rect 3730 1238 3838 1241
rect 842 1228 2473 1231
rect 2482 1228 3209 1231
rect 3218 1228 4598 1231
rect 1466 1218 2214 1221
rect 2470 1221 2473 1228
rect 2470 1218 3197 1221
rect 3206 1221 3209 1228
rect 3206 1218 3485 1221
rect 3490 1218 3558 1221
rect 4386 1218 4486 1221
rect 1198 1212 1201 1217
rect 2834 1208 2941 1211
rect 2946 1208 3294 1211
rect 3298 1208 3469 1211
rect 542 1203 545 1207
rect 541 1202 546 1203
rect 551 1202 552 1207
rect 1566 1203 1569 1207
rect 1565 1202 1570 1203
rect 1575 1202 1576 1207
rect 2590 1203 2593 1207
rect 2589 1202 2594 1203
rect 2599 1202 2600 1207
rect 3614 1203 3617 1207
rect 3613 1202 3618 1203
rect 3623 1202 3624 1207
rect 4638 1203 4641 1207
rect 4637 1202 4642 1203
rect 4647 1202 4648 1207
rect 1626 1198 2273 1201
rect 2770 1198 3374 1201
rect 4530 1198 4582 1201
rect 2270 1191 2273 1198
rect 1338 1188 2265 1191
rect 2270 1188 3302 1191
rect 3346 1188 3638 1191
rect 1026 1178 2253 1181
rect 2262 1181 2265 1188
rect 2262 1178 2622 1181
rect 2802 1178 3678 1181
rect 3714 1178 4358 1181
rect 4362 1178 4685 1181
rect 4690 1178 4702 1181
rect 1994 1168 2093 1171
rect 2154 1168 2654 1171
rect 2706 1168 3182 1171
rect 3386 1168 4054 1171
rect 4058 1168 4342 1171
rect 4530 1168 4534 1171
rect 138 1158 214 1161
rect 962 1158 1389 1161
rect 470 1151 473 1158
rect 3074 1158 3174 1161
rect 3298 1158 3366 1161
rect 3370 1158 3806 1161
rect 3810 1158 3846 1161
rect 4098 1158 4542 1161
rect 470 1148 477 1151
rect 482 1148 838 1151
rect 906 1148 941 1151
rect 1034 1148 1214 1151
rect 1218 1148 1478 1151
rect 1706 1148 2246 1151
rect 2938 1148 3750 1151
rect 3802 1148 3830 1151
rect 4694 1151 4697 1158
rect 4650 1148 4697 1151
rect 754 1138 894 1141
rect 898 1138 1238 1141
rect 1242 1138 1902 1141
rect 1954 1138 2054 1141
rect 2058 1138 2526 1141
rect 2682 1138 3133 1141
rect 3410 1138 4230 1141
rect 626 1128 998 1131
rect 1050 1128 1798 1131
rect 1842 1128 2046 1131
rect 2050 1128 2118 1131
rect 2130 1128 3518 1131
rect 4122 1128 4422 1131
rect 754 1118 870 1121
rect 1026 1118 1213 1121
rect 1562 1118 2062 1121
rect 2594 1118 3126 1121
rect 3138 1118 3405 1121
rect 1362 1108 1710 1111
rect 2138 1108 2845 1111
rect 3154 1108 4078 1111
rect 1054 1103 1057 1107
rect 1053 1102 1058 1103
rect 1063 1102 1064 1107
rect 2078 1103 2081 1107
rect 2077 1102 2082 1103
rect 2087 1102 2088 1107
rect 3102 1103 3105 1107
rect 3101 1102 3106 1103
rect 3111 1102 3112 1107
rect 4118 1103 4121 1107
rect 4117 1102 4122 1103
rect 4127 1102 4128 1107
rect 2258 1098 3078 1101
rect 3666 1098 3670 1101
rect 922 1088 2518 1091
rect 2822 1088 4678 1091
rect 426 1078 854 1081
rect 1650 1078 2590 1081
rect 2822 1081 2825 1088
rect 2610 1078 2825 1081
rect 2994 1078 3486 1081
rect 794 1068 1454 1071
rect 1458 1068 2726 1071
rect 2730 1068 3438 1071
rect 226 1058 862 1061
rect 970 1058 1094 1061
rect 1546 1058 2622 1061
rect 2658 1058 2718 1061
rect 3370 1058 3853 1061
rect 3858 1058 3862 1061
rect 2018 1048 3070 1051
rect 3206 1048 4758 1051
rect 4818 1048 4829 1051
rect 1530 1038 1806 1041
rect 1906 1038 2605 1041
rect 3206 1041 3209 1048
rect 2786 1038 3209 1041
rect 3346 1038 3934 1041
rect 1034 1028 1046 1031
rect 1050 1028 2118 1031
rect 2514 1028 4430 1031
rect 1778 1018 1878 1021
rect 1882 1018 2222 1021
rect 2226 1018 2734 1021
rect 3202 1018 4358 1021
rect 4626 1018 4694 1021
rect 1586 1008 2478 1011
rect 542 1003 545 1007
rect 541 1002 546 1003
rect 551 1002 552 1007
rect 1566 1003 1569 1007
rect 1565 1002 1570 1003
rect 1575 1002 1576 1007
rect 2590 1003 2593 1007
rect 2589 1002 2594 1003
rect 2599 1002 2600 1007
rect 3614 1003 3617 1007
rect 3613 1002 3618 1003
rect 3623 1002 3624 1007
rect 4638 1003 4641 1007
rect 4637 1002 4642 1003
rect 4647 1002 4648 1007
rect 1658 998 2349 1001
rect 2354 998 2374 1001
rect 2610 998 2793 1001
rect 698 988 814 991
rect 890 988 2742 991
rect 2790 991 2793 998
rect 2790 988 4846 991
rect 354 978 598 981
rect 602 978 814 981
rect 818 978 1598 981
rect 1618 978 1774 981
rect 1778 978 2606 981
rect 2666 978 3630 981
rect 1418 968 2558 971
rect 2570 968 4182 971
rect 4330 968 4902 971
rect 802 958 813 961
rect 818 958 1462 961
rect 1834 958 2086 961
rect 2842 958 3294 961
rect 3418 958 4014 961
rect 4674 958 4710 961
rect 1490 948 2654 951
rect 2682 948 3374 951
rect 3890 948 3918 951
rect 3994 948 4333 951
rect 4694 948 4782 951
rect 4694 942 4697 948
rect 714 938 990 941
rect 3314 938 4486 941
rect 4490 938 4678 941
rect 4714 938 4838 941
rect 2378 928 3142 931
rect 3146 928 3565 931
rect 4362 928 5149 931
rect 5154 928 5166 931
rect 1090 918 2205 921
rect 2642 918 2974 921
rect 3298 908 3806 911
rect 3810 908 3965 911
rect 1054 903 1057 907
rect 1053 902 1058 903
rect 1063 902 1064 907
rect 2078 903 2081 907
rect 2077 902 2082 903
rect 2087 902 2088 907
rect 3102 903 3105 907
rect 3101 902 3106 903
rect 3111 902 3112 907
rect 4118 903 4121 907
rect 4117 902 4122 903
rect 4127 902 4128 907
rect 1530 888 1822 891
rect 2050 888 2093 891
rect 2098 888 2102 891
rect 2258 888 2470 891
rect 2474 888 3238 891
rect 3434 888 3926 891
rect 4946 888 4973 891
rect 962 878 982 881
rect 2954 878 2957 881
rect 138 868 462 871
rect 786 868 1949 871
rect 2894 868 3278 871
rect 3354 868 4614 871
rect 2894 862 2897 868
rect 514 858 966 861
rect 1298 858 1630 861
rect 1730 858 2134 861
rect 2138 858 2301 861
rect 2306 858 2846 861
rect 3346 858 3350 861
rect 3386 858 4766 861
rect 5182 852 5185 858
rect 730 848 1086 851
rect 1650 848 1933 851
rect 2274 848 2333 851
rect 2338 848 3174 851
rect 3274 848 3782 851
rect 590 842 593 847
rect 890 838 1430 841
rect 2090 838 3438 841
rect 3442 838 3581 841
rect 3586 838 3934 841
rect 4242 838 4254 841
rect 994 828 1942 831
rect 3850 828 4326 831
rect 1242 818 1622 821
rect 1690 818 2966 821
rect 922 808 1414 811
rect 542 803 545 807
rect 541 802 546 803
rect 551 802 552 807
rect 1566 803 1569 807
rect 1565 802 1570 803
rect 1575 802 1576 807
rect 2590 803 2593 807
rect 2589 802 2594 803
rect 2599 802 2600 807
rect 3614 803 3617 807
rect 3613 802 3618 803
rect 3623 802 3624 807
rect 4638 803 4641 807
rect 4637 802 4642 803
rect 4647 802 4648 807
rect 1610 798 2573 801
rect 2610 798 2798 801
rect 2802 798 3214 801
rect 3282 798 3518 801
rect 1690 788 2766 791
rect 2834 788 3830 791
rect 1426 778 1934 781
rect 1986 778 2614 781
rect 2618 778 2653 781
rect 2658 778 4502 781
rect 306 768 726 771
rect 914 768 925 771
rect 1418 768 2605 771
rect 2802 768 2845 771
rect 1066 758 1590 761
rect 2578 758 2910 761
rect 3134 761 3137 768
rect 3570 768 4557 771
rect 4562 768 4630 771
rect 2914 758 3137 761
rect 3266 758 3309 761
rect 826 748 1678 751
rect 2530 748 3070 751
rect 3730 748 3741 751
rect 3746 748 4086 751
rect 4310 751 4313 758
rect 4306 748 4313 751
rect 4418 748 4510 751
rect 1050 738 1478 741
rect 1482 738 2454 741
rect 2458 738 3230 741
rect 3234 738 3358 741
rect 3722 738 3757 741
rect 4274 738 5062 741
rect 970 728 1094 731
rect 1538 728 2694 731
rect 3210 728 4029 731
rect 4954 728 4966 731
rect 706 718 742 721
rect 746 718 974 721
rect 1938 718 1998 721
rect 2418 718 3094 721
rect 3778 718 4534 721
rect 1054 703 1057 707
rect 1053 702 1058 703
rect 1063 702 1064 707
rect 2078 703 2081 707
rect 2077 702 2082 703
rect 2087 702 2088 707
rect 3102 703 3105 707
rect 3101 702 3106 703
rect 3111 702 3112 707
rect 4118 703 4121 707
rect 4117 702 4122 703
rect 4127 702 4128 707
rect 1714 688 2633 691
rect 3138 688 4854 691
rect 2630 682 2633 688
rect 1250 678 1286 681
rect 1290 678 2006 681
rect 2634 678 4062 681
rect 1682 658 2110 661
rect 2658 658 3062 661
rect 3198 661 3201 668
rect 4750 662 4753 668
rect 3162 658 3201 661
rect 3474 658 4054 661
rect 4754 658 4830 661
rect 1250 648 1758 651
rect 2106 648 2109 651
rect 2426 648 2926 651
rect 2930 648 5038 651
rect 1106 638 1757 641
rect 1762 638 2422 641
rect 3522 628 4621 631
rect 714 618 758 621
rect 762 618 1518 621
rect 1522 618 2142 621
rect 542 603 545 607
rect 541 602 546 603
rect 551 602 552 607
rect 1566 603 1569 607
rect 1565 602 1570 603
rect 1575 602 1576 607
rect 2590 603 2593 607
rect 2589 602 2594 603
rect 2599 602 2600 607
rect 3614 603 3617 607
rect 3613 602 3618 603
rect 3623 602 3624 607
rect 4638 603 4641 607
rect 4637 602 4642 603
rect 4647 602 4648 607
rect 874 588 1805 591
rect 1810 588 2398 591
rect 3018 588 3998 591
rect 2970 578 5006 581
rect 946 568 1070 571
rect 1546 568 2030 571
rect 594 558 902 561
rect 930 558 2062 561
rect 2306 558 3534 561
rect 3538 558 3558 561
rect 3562 558 4030 561
rect 202 548 862 551
rect 930 548 1686 551
rect 1938 548 2798 551
rect 2802 548 3501 551
rect 3578 548 4406 551
rect 4410 548 4494 551
rect 642 538 1254 541
rect 1450 538 2246 541
rect 3458 538 4054 541
rect 4478 532 4481 538
rect 642 528 934 531
rect 1194 528 1469 531
rect 1474 528 2998 531
rect 3426 528 4477 531
rect 570 518 686 521
rect 690 518 854 521
rect 858 518 1070 521
rect 1138 518 2342 521
rect 3422 521 3425 528
rect 2402 518 3425 521
rect 3650 518 4126 521
rect 1054 503 1057 507
rect 1053 502 1058 503
rect 1063 502 1064 507
rect 2078 503 2081 507
rect 2077 502 2082 503
rect 2087 502 2088 507
rect 3102 503 3105 507
rect 3101 502 3106 503
rect 3111 502 3112 507
rect 4118 503 4121 507
rect 4117 502 4122 503
rect 4127 502 4128 507
rect 1622 488 3302 491
rect 1622 481 1625 488
rect 1042 478 1625 481
rect 1778 478 2910 481
rect 354 468 422 471
rect 2650 468 4206 471
rect 4314 468 4382 471
rect 626 458 838 461
rect 958 461 961 468
rect 958 458 1398 461
rect 1518 452 1521 457
rect 4030 452 4033 458
rect 1930 448 2830 451
rect 542 403 545 407
rect 541 402 546 403
rect 551 402 552 407
rect 1566 403 1569 407
rect 1565 402 1570 403
rect 1575 402 1576 407
rect 2590 403 2593 407
rect 2589 402 2594 403
rect 2599 402 2600 407
rect 3614 403 3617 407
rect 3613 402 3618 403
rect 3623 402 3624 407
rect 4638 403 4641 407
rect 4637 402 4642 403
rect 4647 402 4648 407
rect 1402 388 2014 391
rect 1274 378 1750 381
rect 1330 368 1425 371
rect 1698 368 2670 371
rect 3650 368 3686 371
rect 1422 362 1425 368
rect 354 348 782 351
rect 2186 348 2686 351
rect 3874 348 3958 351
rect 4146 348 4198 351
rect 4490 348 4526 351
rect 874 338 1350 341
rect 2994 338 3254 341
rect 194 328 598 331
rect 1054 303 1057 307
rect 1053 302 1058 303
rect 1063 302 1064 307
rect 2078 303 2081 307
rect 2077 302 2082 303
rect 2087 302 2088 307
rect 3102 303 3105 307
rect 3101 302 3106 303
rect 3111 302 3112 307
rect 4118 303 4121 307
rect 4117 302 4122 303
rect 4127 302 4128 307
rect 450 288 862 291
rect 5122 288 5182 291
rect 1082 278 1325 281
rect 1330 278 1526 281
rect 1530 278 2438 281
rect 138 268 454 271
rect 2170 268 2238 271
rect 2786 268 4174 271
rect 4862 262 4865 267
rect 1890 258 2206 261
rect 2874 258 3805 261
rect 3810 258 4286 261
rect 4290 258 4366 261
rect 554 238 1062 241
rect 542 203 545 207
rect 541 202 546 203
rect 551 202 552 207
rect 1566 203 1569 207
rect 1565 202 1570 203
rect 1575 202 1576 207
rect 2590 203 2593 207
rect 2589 202 2594 203
rect 2599 202 2600 207
rect 3614 203 3617 207
rect 3613 202 3618 203
rect 3623 202 3624 207
rect 4638 203 4641 207
rect 4637 202 4642 203
rect 4647 202 4648 207
rect 5106 188 5110 191
rect 3486 152 3489 157
rect 226 148 534 151
rect 1458 148 1486 151
rect 2514 148 2518 151
rect 1770 138 1926 141
rect 2842 138 3406 141
rect 3410 138 4038 141
rect 4042 138 4214 141
rect 4234 138 4518 141
rect 4570 138 4669 141
rect 2594 128 2726 131
rect 2378 118 2750 121
rect 4602 108 4605 111
rect 1054 103 1057 107
rect 1053 102 1058 103
rect 1063 102 1064 107
rect 2078 103 2081 107
rect 2077 102 2082 103
rect 2087 102 2088 107
rect 3102 103 3105 107
rect 3101 102 3106 103
rect 3111 102 3112 107
rect 4118 103 4121 107
rect 4117 102 4122 103
rect 4127 102 4128 107
rect 5010 88 5014 91
rect 3674 78 4206 81
rect 4210 78 4398 81
rect 4954 78 4957 81
rect 354 68 974 71
rect 2378 68 2686 71
rect 3954 68 4086 71
rect 4090 68 4438 71
rect 4542 62 4545 68
rect 810 58 934 61
rect 2290 58 2750 61
rect 3418 58 3510 61
rect 4698 58 4717 61
rect 4762 58 5142 61
rect 2658 48 2822 51
rect 4050 48 4126 51
rect 4562 48 4589 51
rect 4818 48 4822 51
rect 542 3 545 7
rect 541 2 546 3
rect 551 2 552 7
rect 1566 3 1569 7
rect 1565 2 1570 3
rect 1575 2 1576 7
rect 2590 3 2593 7
rect 2589 2 2594 3
rect 2599 2 2600 7
rect 3614 3 3617 7
rect 3613 2 3618 3
rect 3623 2 3624 7
rect 4638 3 4641 7
rect 4637 2 4642 3
rect 4647 2 4648 7
<< m6contact >>
rect 1048 4903 1050 4907
rect 1050 4903 1053 4907
rect 1058 4903 1061 4907
rect 1061 4903 1063 4907
rect 1048 4902 1053 4903
rect 1058 4902 1063 4903
rect 2072 4903 2074 4907
rect 2074 4903 2077 4907
rect 2082 4903 2085 4907
rect 2085 4903 2087 4907
rect 2072 4902 2077 4903
rect 2082 4902 2087 4903
rect 3096 4903 3098 4907
rect 3098 4903 3101 4907
rect 3106 4903 3109 4907
rect 3109 4903 3111 4907
rect 3096 4902 3101 4903
rect 3106 4902 3111 4903
rect 4112 4903 4114 4907
rect 4114 4903 4117 4907
rect 4122 4903 4125 4907
rect 4125 4903 4127 4907
rect 4112 4902 4117 4903
rect 4122 4902 4127 4903
rect 2381 4857 2386 4862
rect 5101 4857 5106 4862
rect 4861 4847 4866 4852
rect 4925 4847 4930 4852
rect 536 4803 538 4807
rect 538 4803 541 4807
rect 546 4803 549 4807
rect 549 4803 551 4807
rect 536 4802 541 4803
rect 546 4802 551 4803
rect 1560 4803 1562 4807
rect 1562 4803 1565 4807
rect 1570 4803 1573 4807
rect 1573 4803 1575 4807
rect 1560 4802 1565 4803
rect 1570 4802 1575 4803
rect 2584 4803 2586 4807
rect 2586 4803 2589 4807
rect 2594 4803 2597 4807
rect 2597 4803 2599 4807
rect 2584 4802 2589 4803
rect 2594 4802 2599 4803
rect 3608 4803 3610 4807
rect 3610 4803 3613 4807
rect 3618 4803 3621 4807
rect 3621 4803 3623 4807
rect 3608 4802 3613 4803
rect 3618 4802 3623 4803
rect 4632 4803 4634 4807
rect 4634 4803 4637 4807
rect 4642 4803 4645 4807
rect 4645 4803 4647 4807
rect 4632 4802 4637 4803
rect 4642 4802 4647 4803
rect 1048 4703 1050 4707
rect 1050 4703 1053 4707
rect 1058 4703 1061 4707
rect 1061 4703 1063 4707
rect 1048 4702 1053 4703
rect 1058 4702 1063 4703
rect 2072 4703 2074 4707
rect 2074 4703 2077 4707
rect 2082 4703 2085 4707
rect 2085 4703 2087 4707
rect 2072 4702 2077 4703
rect 2082 4702 2087 4703
rect 3096 4703 3098 4707
rect 3098 4703 3101 4707
rect 3106 4703 3109 4707
rect 3109 4703 3111 4707
rect 3096 4702 3101 4703
rect 3106 4702 3111 4703
rect 4112 4703 4114 4707
rect 4114 4703 4117 4707
rect 4122 4703 4125 4707
rect 4125 4703 4127 4707
rect 4112 4702 4117 4703
rect 4122 4702 4127 4703
rect 1597 4637 1602 4642
rect 536 4603 538 4607
rect 538 4603 541 4607
rect 546 4603 549 4607
rect 549 4603 551 4607
rect 536 4602 541 4603
rect 546 4602 551 4603
rect 1560 4603 1562 4607
rect 1562 4603 1565 4607
rect 1570 4603 1573 4607
rect 1573 4603 1575 4607
rect 1560 4602 1565 4603
rect 1570 4602 1575 4603
rect 2584 4603 2586 4607
rect 2586 4603 2589 4607
rect 2594 4603 2597 4607
rect 2597 4603 2599 4607
rect 2584 4602 2589 4603
rect 2594 4602 2599 4603
rect 3608 4603 3610 4607
rect 3610 4603 3613 4607
rect 3618 4603 3621 4607
rect 3621 4603 3623 4607
rect 3608 4602 3613 4603
rect 3618 4602 3623 4603
rect 4632 4603 4634 4607
rect 4634 4603 4637 4607
rect 4642 4603 4645 4607
rect 4645 4603 4647 4607
rect 4632 4602 4637 4603
rect 4642 4602 4647 4603
rect 749 4537 754 4542
rect 1629 4527 1634 4532
rect 3549 4517 3554 4522
rect 1048 4503 1050 4507
rect 1050 4503 1053 4507
rect 1058 4503 1061 4507
rect 1061 4503 1063 4507
rect 1048 4502 1053 4503
rect 1058 4502 1063 4503
rect 2072 4503 2074 4507
rect 2074 4503 2077 4507
rect 2082 4503 2085 4507
rect 2085 4503 2087 4507
rect 2072 4502 2077 4503
rect 2082 4502 2087 4503
rect 3096 4503 3098 4507
rect 3098 4503 3101 4507
rect 3106 4503 3109 4507
rect 3109 4503 3111 4507
rect 3096 4502 3101 4503
rect 3106 4502 3111 4503
rect 4112 4503 4114 4507
rect 4114 4503 4117 4507
rect 4122 4503 4125 4507
rect 4125 4503 4127 4507
rect 4112 4502 4117 4503
rect 4122 4502 4127 4503
rect 4749 4457 4754 4462
rect 1661 4447 1666 4452
rect 2733 4437 2738 4442
rect 2333 4427 2338 4432
rect 4397 4407 4402 4412
rect 536 4403 538 4407
rect 538 4403 541 4407
rect 546 4403 549 4407
rect 549 4403 551 4407
rect 536 4402 541 4403
rect 546 4402 551 4403
rect 1560 4403 1562 4407
rect 1562 4403 1565 4407
rect 1570 4403 1573 4407
rect 1573 4403 1575 4407
rect 1560 4402 1565 4403
rect 1570 4402 1575 4403
rect 2584 4403 2586 4407
rect 2586 4403 2589 4407
rect 2594 4403 2597 4407
rect 2597 4403 2599 4407
rect 2584 4402 2589 4403
rect 2594 4402 2599 4403
rect 3608 4403 3610 4407
rect 3610 4403 3613 4407
rect 3618 4403 3621 4407
rect 3621 4403 3623 4407
rect 3608 4402 3613 4403
rect 3618 4402 3623 4403
rect 4632 4403 4634 4407
rect 4634 4403 4637 4407
rect 4642 4403 4645 4407
rect 4645 4403 4647 4407
rect 4632 4402 4637 4403
rect 4642 4402 4647 4403
rect 4541 4397 4546 4402
rect 1805 4387 1810 4392
rect 3549 4387 3554 4392
rect 2717 4367 2722 4372
rect 2733 4367 2738 4372
rect 5069 4367 5074 4372
rect 493 4347 498 4352
rect 4557 4337 4562 4342
rect 2717 4327 2722 4332
rect 781 4317 786 4322
rect 2189 4307 2194 4312
rect 3933 4307 3938 4312
rect 1048 4303 1050 4307
rect 1050 4303 1053 4307
rect 1058 4303 1061 4307
rect 1061 4303 1063 4307
rect 1048 4302 1053 4303
rect 1058 4302 1063 4303
rect 2072 4303 2074 4307
rect 2074 4303 2077 4307
rect 2082 4303 2085 4307
rect 2085 4303 2087 4307
rect 2072 4302 2077 4303
rect 2082 4302 2087 4303
rect 3096 4303 3098 4307
rect 3098 4303 3101 4307
rect 3106 4303 3109 4307
rect 3109 4303 3111 4307
rect 3096 4302 3101 4303
rect 3106 4302 3111 4303
rect 4112 4303 4114 4307
rect 4114 4303 4117 4307
rect 4122 4303 4125 4307
rect 4125 4303 4127 4307
rect 4112 4302 4117 4303
rect 4122 4302 4127 4303
rect 3533 4267 3538 4272
rect 2557 4257 2562 4262
rect 4269 4257 4274 4262
rect 2477 4247 2482 4252
rect 3533 4247 3538 4252
rect 4013 4247 4018 4252
rect 2477 4227 2482 4232
rect 4397 4227 4402 4232
rect 4045 4217 4050 4222
rect 536 4203 538 4207
rect 538 4203 541 4207
rect 546 4203 549 4207
rect 549 4203 551 4207
rect 536 4202 541 4203
rect 546 4202 551 4203
rect 1560 4203 1562 4207
rect 1562 4203 1565 4207
rect 1570 4203 1573 4207
rect 1573 4203 1575 4207
rect 1560 4202 1565 4203
rect 1570 4202 1575 4203
rect 2584 4203 2586 4207
rect 2586 4203 2589 4207
rect 2594 4203 2597 4207
rect 2597 4203 2599 4207
rect 2584 4202 2589 4203
rect 2594 4202 2599 4203
rect 3608 4203 3610 4207
rect 3610 4203 3613 4207
rect 3618 4203 3621 4207
rect 3621 4203 3623 4207
rect 3608 4202 3613 4203
rect 3618 4202 3623 4203
rect 4632 4203 4634 4207
rect 4634 4203 4637 4207
rect 4642 4203 4645 4207
rect 4645 4203 4647 4207
rect 4632 4202 4637 4203
rect 4642 4202 4647 4203
rect 3133 4197 3138 4202
rect 2941 4187 2946 4192
rect 3437 4187 3442 4192
rect 2173 4167 2178 4172
rect 3133 4177 3138 4182
rect 4621 4177 4626 4182
rect 2941 4157 2946 4162
rect 3981 4137 3986 4142
rect 4525 4137 4530 4142
rect 1261 4117 1266 4122
rect 1048 4103 1050 4107
rect 1050 4103 1053 4107
rect 1058 4103 1061 4107
rect 1061 4103 1063 4107
rect 1048 4102 1053 4103
rect 1058 4102 1063 4103
rect 2072 4103 2074 4107
rect 2074 4103 2077 4107
rect 2082 4103 2085 4107
rect 2085 4103 2087 4107
rect 2072 4102 2077 4103
rect 2082 4102 2087 4103
rect 3096 4103 3098 4107
rect 3098 4103 3101 4107
rect 3106 4103 3109 4107
rect 3109 4103 3111 4107
rect 3096 4102 3101 4103
rect 3106 4102 3111 4103
rect 4112 4103 4114 4107
rect 4114 4103 4117 4107
rect 4122 4103 4125 4107
rect 4125 4103 4127 4107
rect 4112 4102 4117 4103
rect 4122 4102 4127 4103
rect 2365 4057 2370 4062
rect 4061 4047 4066 4052
rect 4101 4047 4106 4052
rect 2829 4037 2834 4042
rect 2365 4027 2370 4032
rect 4973 4017 4978 4022
rect 536 4003 538 4007
rect 538 4003 541 4007
rect 546 4003 549 4007
rect 549 4003 551 4007
rect 536 4002 541 4003
rect 546 4002 551 4003
rect 1560 4003 1562 4007
rect 1562 4003 1565 4007
rect 1570 4003 1573 4007
rect 1573 4003 1575 4007
rect 1560 4002 1565 4003
rect 1570 4002 1575 4003
rect 2584 4003 2586 4007
rect 2586 4003 2589 4007
rect 2594 4003 2597 4007
rect 2597 4003 2599 4007
rect 2584 4002 2589 4003
rect 2594 4002 2599 4003
rect 3608 4003 3610 4007
rect 3610 4003 3613 4007
rect 3618 4003 3621 4007
rect 3621 4003 3623 4007
rect 3608 4002 3613 4003
rect 3618 4002 3623 4003
rect 4632 4003 4634 4007
rect 4634 4003 4637 4007
rect 4642 4003 4645 4007
rect 4645 4003 4647 4007
rect 4632 4002 4637 4003
rect 4642 4002 4647 4003
rect 2989 3997 2994 4002
rect 5149 3997 5154 4002
rect 3341 3977 3346 3982
rect 2493 3957 2498 3962
rect 3293 3947 3298 3952
rect 4765 3937 4770 3942
rect 4573 3927 4578 3932
rect 2061 3907 2066 3912
rect 3389 3907 3394 3912
rect 1048 3903 1050 3907
rect 1050 3903 1053 3907
rect 1058 3903 1061 3907
rect 1061 3903 1063 3907
rect 1048 3902 1053 3903
rect 1058 3902 1063 3903
rect 2072 3903 2074 3907
rect 2074 3903 2077 3907
rect 2082 3903 2085 3907
rect 2085 3903 2087 3907
rect 2072 3902 2077 3903
rect 2082 3902 2087 3903
rect 3096 3903 3098 3907
rect 3098 3903 3101 3907
rect 3106 3903 3109 3907
rect 3109 3903 3111 3907
rect 3096 3902 3101 3903
rect 3106 3902 3111 3903
rect 4112 3903 4114 3907
rect 4114 3903 4117 3907
rect 4122 3903 4125 3907
rect 4125 3903 4127 3907
rect 4112 3902 4117 3903
rect 4122 3902 4127 3903
rect 909 3887 914 3892
rect 2397 3887 2402 3892
rect 797 3867 802 3872
rect 4221 3857 4226 3862
rect 1549 3847 1554 3852
rect 3405 3837 3410 3842
rect 4285 3837 4290 3842
rect 2413 3817 2418 3822
rect 3597 3817 3602 3822
rect 3213 3807 3218 3812
rect 4509 3807 4514 3812
rect 536 3803 538 3807
rect 538 3803 541 3807
rect 546 3803 549 3807
rect 549 3803 551 3807
rect 536 3802 541 3803
rect 546 3802 551 3803
rect 1560 3803 1562 3807
rect 1562 3803 1565 3807
rect 1570 3803 1573 3807
rect 1573 3803 1575 3807
rect 1560 3802 1565 3803
rect 1570 3802 1575 3803
rect 2584 3803 2586 3807
rect 2586 3803 2589 3807
rect 2594 3803 2597 3807
rect 2597 3803 2599 3807
rect 2584 3802 2589 3803
rect 2594 3802 2599 3803
rect 3608 3803 3610 3807
rect 3610 3803 3613 3807
rect 3618 3803 3621 3807
rect 3621 3803 3623 3807
rect 3608 3802 3613 3803
rect 3618 3802 3623 3803
rect 4632 3803 4634 3807
rect 4634 3803 4637 3807
rect 4642 3803 4645 3807
rect 4645 3803 4647 3807
rect 4632 3802 4637 3803
rect 4642 3802 4647 3803
rect 2157 3787 2162 3792
rect 1725 3767 1730 3772
rect 3485 3757 3490 3762
rect 381 3747 386 3752
rect 1933 3737 1938 3742
rect 2029 3737 2034 3742
rect 1949 3727 1954 3732
rect 2397 3727 2402 3732
rect 3533 3727 3538 3732
rect 1405 3717 1410 3722
rect 2061 3717 2066 3722
rect 3725 3717 3730 3722
rect 2221 3707 2226 3712
rect 2989 3707 2994 3712
rect 1048 3703 1050 3707
rect 1050 3703 1053 3707
rect 1058 3703 1061 3707
rect 1061 3703 1063 3707
rect 1048 3702 1053 3703
rect 1058 3702 1063 3703
rect 2072 3703 2074 3707
rect 2074 3703 2077 3707
rect 2082 3703 2085 3707
rect 2085 3703 2087 3707
rect 2072 3702 2077 3703
rect 2082 3702 2087 3703
rect 3096 3703 3098 3707
rect 3098 3703 3101 3707
rect 3106 3703 3109 3707
rect 3109 3703 3111 3707
rect 3096 3702 3101 3703
rect 3106 3702 3111 3703
rect 4112 3703 4114 3707
rect 4114 3703 4117 3707
rect 4122 3703 4125 3707
rect 4125 3703 4127 3707
rect 4112 3702 4117 3703
rect 4122 3702 4127 3703
rect 1037 3697 1042 3702
rect 1597 3697 1602 3702
rect 1709 3697 1714 3702
rect 2317 3697 2322 3702
rect 669 3687 674 3692
rect 2317 3677 2322 3682
rect 2749 3677 2754 3682
rect 3485 3677 3490 3682
rect 3069 3657 3074 3662
rect 3949 3657 3954 3662
rect 4589 3657 4594 3662
rect 1821 3647 1826 3652
rect 4333 3647 4338 3652
rect 1085 3637 1090 3642
rect 3373 3637 3378 3642
rect 4077 3637 4082 3642
rect 1853 3627 1858 3632
rect 3757 3627 3762 3632
rect 3405 3617 3410 3622
rect 2285 3607 2290 3612
rect 2477 3607 2482 3612
rect 3517 3607 3522 3612
rect 4573 3607 4578 3612
rect 536 3603 538 3607
rect 538 3603 541 3607
rect 546 3603 549 3607
rect 549 3603 551 3607
rect 536 3602 541 3603
rect 546 3602 551 3603
rect 1560 3603 1562 3607
rect 1562 3603 1565 3607
rect 1570 3603 1573 3607
rect 1573 3603 1575 3607
rect 1560 3602 1565 3603
rect 1570 3602 1575 3603
rect 2584 3603 2586 3607
rect 2586 3603 2589 3607
rect 2594 3603 2597 3607
rect 2597 3603 2599 3607
rect 2584 3602 2589 3603
rect 2594 3602 2599 3603
rect 3608 3603 3610 3607
rect 3610 3603 3613 3607
rect 3618 3603 3621 3607
rect 3621 3603 3623 3607
rect 3608 3602 3613 3603
rect 3618 3602 3623 3603
rect 4632 3603 4634 3607
rect 4634 3603 4637 3607
rect 4642 3603 4645 3607
rect 4645 3603 4647 3607
rect 4632 3602 4637 3603
rect 4642 3602 4647 3603
rect 1309 3597 1314 3602
rect 2093 3597 2098 3602
rect 4269 3587 4274 3592
rect 1741 3577 1746 3582
rect 2093 3577 2098 3582
rect 3421 3567 3426 3572
rect 3645 3557 3650 3562
rect 3677 3557 3682 3562
rect 1661 3537 1666 3542
rect 1437 3517 1442 3522
rect 1453 3517 1458 3522
rect 3917 3507 3922 3512
rect 4269 3507 4274 3512
rect 1048 3503 1050 3507
rect 1050 3503 1053 3507
rect 1058 3503 1061 3507
rect 1061 3503 1063 3507
rect 1048 3502 1053 3503
rect 1058 3502 1063 3503
rect 2072 3503 2074 3507
rect 2074 3503 2077 3507
rect 2082 3503 2085 3507
rect 2085 3503 2087 3507
rect 2072 3502 2077 3503
rect 2082 3502 2087 3503
rect 3096 3503 3098 3507
rect 3098 3503 3101 3507
rect 3106 3503 3109 3507
rect 3109 3503 3111 3507
rect 3096 3502 3101 3503
rect 3106 3502 3111 3503
rect 4112 3503 4114 3507
rect 4114 3503 4117 3507
rect 4122 3503 4125 3507
rect 4125 3503 4127 3507
rect 4112 3502 4117 3503
rect 4122 3502 4127 3503
rect 477 3497 482 3502
rect 1469 3497 1474 3502
rect 2173 3497 2178 3502
rect 2541 3497 2546 3502
rect 3821 3497 3826 3502
rect 1821 3487 1826 3492
rect 765 3477 770 3482
rect 1453 3467 1458 3472
rect 1069 3457 1074 3462
rect 2541 3467 2546 3472
rect 3629 3467 3634 3472
rect 4373 3467 4378 3472
rect 4397 3467 4402 3472
rect 4685 3467 4690 3472
rect 2381 3457 2386 3462
rect 685 3447 690 3452
rect 1917 3437 1922 3442
rect 1277 3427 1282 3432
rect 3597 3427 3602 3432
rect 877 3417 882 3422
rect 1357 3417 1362 3422
rect 1581 3417 1586 3422
rect 1789 3417 1794 3422
rect 733 3407 738 3412
rect 1133 3407 1138 3412
rect 536 3403 538 3407
rect 538 3403 541 3407
rect 546 3403 549 3407
rect 549 3403 551 3407
rect 536 3402 541 3403
rect 546 3402 551 3403
rect 1560 3403 1562 3407
rect 1562 3403 1565 3407
rect 1570 3403 1573 3407
rect 1573 3403 1575 3407
rect 1560 3402 1565 3403
rect 1570 3402 1575 3403
rect 2584 3403 2586 3407
rect 2586 3403 2589 3407
rect 2594 3403 2597 3407
rect 2597 3403 2599 3407
rect 2584 3402 2589 3403
rect 2594 3402 2599 3403
rect 3608 3403 3610 3407
rect 3610 3403 3613 3407
rect 3618 3403 3621 3407
rect 3621 3403 3623 3407
rect 3608 3402 3613 3403
rect 3618 3402 3623 3403
rect 4632 3403 4634 3407
rect 4634 3403 4637 3407
rect 4642 3403 4645 3407
rect 4645 3403 4647 3407
rect 4632 3402 4637 3403
rect 4642 3402 4647 3403
rect 685 3397 690 3402
rect 3309 3397 3314 3402
rect 4557 3387 4562 3392
rect 3293 3367 3298 3372
rect 2029 3357 2034 3362
rect 1629 3347 1634 3352
rect 1197 3337 1202 3342
rect 4477 3337 4482 3342
rect 4541 3337 4546 3342
rect 1453 3327 1458 3332
rect 2029 3327 2034 3332
rect 2125 3327 2130 3332
rect 1645 3317 1650 3322
rect 1357 3307 1362 3312
rect 2557 3307 2562 3312
rect 4205 3307 4210 3312
rect 1048 3303 1050 3307
rect 1050 3303 1053 3307
rect 1058 3303 1061 3307
rect 1061 3303 1063 3307
rect 1048 3302 1053 3303
rect 1058 3302 1063 3303
rect 2072 3303 2074 3307
rect 2074 3303 2077 3307
rect 2082 3303 2085 3307
rect 2085 3303 2087 3307
rect 2072 3302 2077 3303
rect 2082 3302 2087 3303
rect 3096 3303 3098 3307
rect 3098 3303 3101 3307
rect 3106 3303 3109 3307
rect 3109 3303 3111 3307
rect 3096 3302 3101 3303
rect 3106 3302 3111 3303
rect 4112 3303 4114 3307
rect 4114 3303 4117 3307
rect 4122 3303 4125 3307
rect 4125 3303 4127 3307
rect 4112 3302 4117 3303
rect 4122 3302 4127 3303
rect 1757 3297 1762 3302
rect 4029 3297 4034 3302
rect 949 3287 954 3292
rect 1629 3277 1634 3282
rect 2125 3277 2130 3282
rect 3197 3277 3202 3282
rect 3981 3277 3986 3282
rect 3085 3267 3090 3272
rect 925 3257 930 3262
rect 2669 3257 2674 3262
rect 3037 3247 3042 3252
rect 3741 3247 3746 3252
rect 957 3237 962 3242
rect 2013 3237 2018 3242
rect 1341 3227 1346 3232
rect 1485 3227 1490 3232
rect 1629 3227 1634 3232
rect 2701 3227 2706 3232
rect 3373 3217 3378 3222
rect 1149 3207 1154 3212
rect 1325 3207 1330 3212
rect 1709 3207 1714 3212
rect 1933 3207 1938 3212
rect 536 3203 538 3207
rect 538 3203 541 3207
rect 546 3203 549 3207
rect 549 3203 551 3207
rect 536 3202 541 3203
rect 546 3202 551 3203
rect 1560 3203 1562 3207
rect 1562 3203 1565 3207
rect 1570 3203 1573 3207
rect 1573 3203 1575 3207
rect 1560 3202 1565 3203
rect 1570 3202 1575 3203
rect 2584 3203 2586 3207
rect 2586 3203 2589 3207
rect 2594 3203 2597 3207
rect 2597 3203 2599 3207
rect 2584 3202 2589 3203
rect 2594 3202 2599 3203
rect 3608 3203 3610 3207
rect 3610 3203 3613 3207
rect 3618 3203 3621 3207
rect 3621 3203 3623 3207
rect 3608 3202 3613 3203
rect 3618 3202 3623 3203
rect 4632 3203 4634 3207
rect 4634 3203 4637 3207
rect 4642 3203 4645 3207
rect 4645 3203 4647 3207
rect 4632 3202 4637 3203
rect 4642 3202 4647 3203
rect 2397 3197 2402 3202
rect 829 3177 834 3182
rect 1069 3177 1074 3182
rect 2733 3177 2738 3182
rect 4525 3177 4530 3182
rect 1389 3167 1394 3172
rect 1293 3157 1298 3162
rect 1773 3157 1778 3162
rect 2141 3157 2146 3162
rect 717 3147 722 3152
rect 1533 3147 1538 3152
rect 3469 3157 3474 3162
rect 4013 3157 4018 3162
rect 1165 3137 1170 3142
rect 2061 3137 2066 3142
rect 2109 3137 2114 3142
rect 3581 3137 3586 3142
rect 4525 3147 4530 3152
rect 4733 3137 4738 3142
rect 1421 3127 1426 3132
rect 3197 3127 3202 3132
rect 1837 3117 1842 3122
rect 2285 3117 2290 3122
rect 2685 3117 2690 3122
rect 3133 3117 3138 3122
rect 2621 3107 2626 3112
rect 2941 3107 2946 3112
rect 1048 3103 1050 3107
rect 1050 3103 1053 3107
rect 1058 3103 1061 3107
rect 1061 3103 1063 3107
rect 1048 3102 1053 3103
rect 1058 3102 1063 3103
rect 2072 3103 2074 3107
rect 2074 3103 2077 3107
rect 2082 3103 2085 3107
rect 2085 3103 2087 3107
rect 2072 3102 2077 3103
rect 2082 3102 2087 3103
rect 3096 3103 3098 3107
rect 3098 3103 3101 3107
rect 3106 3103 3109 3107
rect 3109 3103 3111 3107
rect 3096 3102 3101 3103
rect 3106 3102 3111 3103
rect 4112 3103 4114 3107
rect 4114 3103 4117 3107
rect 4122 3103 4125 3107
rect 4125 3103 4127 3107
rect 4112 3102 4117 3103
rect 4122 3102 4127 3103
rect 2301 3097 2306 3102
rect 1485 3087 1490 3092
rect 2269 3087 2274 3092
rect 3181 3067 3186 3072
rect 3325 3067 3330 3072
rect 3917 3067 3922 3072
rect 1597 3057 1602 3062
rect 2301 3057 2306 3062
rect 5165 3047 5170 3052
rect 1213 3037 1218 3042
rect 1261 3037 1266 3042
rect 1725 3037 1730 3042
rect 941 3027 946 3032
rect 1357 3027 1362 3032
rect 4157 3027 4162 3032
rect 1037 3017 1042 3022
rect 1213 3017 1218 3022
rect 1981 3017 1986 3022
rect 2045 3017 2050 3022
rect 4093 3017 4098 3022
rect 2221 3007 2226 3012
rect 2749 3007 2754 3012
rect 4189 3007 4194 3012
rect 536 3003 538 3007
rect 538 3003 541 3007
rect 546 3003 549 3007
rect 549 3003 551 3007
rect 536 3002 541 3003
rect 546 3002 551 3003
rect 1560 3003 1562 3007
rect 1562 3003 1565 3007
rect 1570 3003 1573 3007
rect 1573 3003 1575 3007
rect 1560 3002 1565 3003
rect 1570 3002 1575 3003
rect 2584 3003 2586 3007
rect 2586 3003 2589 3007
rect 2594 3003 2597 3007
rect 2597 3003 2599 3007
rect 2584 3002 2589 3003
rect 2594 3002 2599 3003
rect 3608 3003 3610 3007
rect 3610 3003 3613 3007
rect 3618 3003 3621 3007
rect 3621 3003 3623 3007
rect 3608 3002 3613 3003
rect 3618 3002 3623 3003
rect 4632 3003 4634 3007
rect 4634 3003 4637 3007
rect 4642 3003 4645 3007
rect 4645 3003 4647 3007
rect 4632 3002 4637 3003
rect 4642 3002 4647 3003
rect 1965 2997 1970 3002
rect 2573 2997 2578 3002
rect 4045 2997 4050 3002
rect 1213 2987 1218 2992
rect 3933 2987 3938 2992
rect 4253 2987 4258 2992
rect 941 2977 946 2982
rect 1709 2977 1714 2982
rect 2573 2977 2578 2982
rect 3645 2977 3650 2982
rect 3869 2977 3874 2982
rect 4461 2967 4466 2972
rect 797 2947 802 2952
rect 861 2947 866 2952
rect 1901 2947 1906 2952
rect 3549 2947 3554 2952
rect 3629 2947 3634 2952
rect 5117 2947 5122 2952
rect 1037 2937 1042 2942
rect 2653 2937 2658 2942
rect 1309 2927 1314 2932
rect 1501 2927 1506 2932
rect 1885 2927 1890 2932
rect 1901 2917 1906 2922
rect 4173 2927 4178 2932
rect 4093 2917 4098 2922
rect 1181 2907 1186 2912
rect 2125 2907 2130 2912
rect 3165 2907 3170 2912
rect 1048 2903 1050 2907
rect 1050 2903 1053 2907
rect 1058 2903 1061 2907
rect 1061 2903 1063 2907
rect 1048 2902 1053 2903
rect 1058 2902 1063 2903
rect 2072 2903 2074 2907
rect 2074 2903 2077 2907
rect 2082 2903 2085 2907
rect 2085 2903 2087 2907
rect 2072 2902 2077 2903
rect 2082 2902 2087 2903
rect 3096 2903 3098 2907
rect 3098 2903 3101 2907
rect 3106 2903 3109 2907
rect 3109 2903 3111 2907
rect 3096 2902 3101 2903
rect 3106 2902 3111 2903
rect 5021 2907 5026 2912
rect 4112 2903 4114 2907
rect 4114 2903 4117 2907
rect 4122 2903 4125 2907
rect 4125 2903 4127 2907
rect 4112 2902 4117 2903
rect 4122 2902 4127 2903
rect 1645 2897 1650 2902
rect 2317 2887 2322 2892
rect 3965 2897 3970 2902
rect 3405 2887 3410 2892
rect 3773 2887 3778 2892
rect 3997 2887 4002 2892
rect 4301 2887 4306 2892
rect 5069 2887 5074 2892
rect 1373 2877 1378 2882
rect 2157 2877 2162 2882
rect 2541 2877 2546 2882
rect 3837 2878 3838 2882
rect 3838 2878 3842 2882
rect 3837 2877 3842 2878
rect 4621 2877 4626 2882
rect 1021 2867 1026 2872
rect 3405 2867 3410 2872
rect 3933 2867 3938 2872
rect 2621 2857 2626 2862
rect 2125 2847 2130 2852
rect 1437 2837 1442 2842
rect 3661 2837 3666 2842
rect 1629 2807 1634 2812
rect 2509 2807 2514 2812
rect 4381 2807 4386 2812
rect 536 2803 538 2807
rect 538 2803 541 2807
rect 546 2803 549 2807
rect 549 2803 551 2807
rect 536 2802 541 2803
rect 546 2802 551 2803
rect 1560 2803 1562 2807
rect 1562 2803 1565 2807
rect 1570 2803 1573 2807
rect 1573 2803 1575 2807
rect 1560 2802 1565 2803
rect 1570 2802 1575 2803
rect 2584 2803 2586 2807
rect 2586 2803 2589 2807
rect 2594 2803 2597 2807
rect 2597 2803 2599 2807
rect 2584 2802 2589 2803
rect 2594 2802 2599 2803
rect 3608 2803 3610 2807
rect 3610 2803 3613 2807
rect 3618 2803 3621 2807
rect 3621 2803 3623 2807
rect 3608 2802 3613 2803
rect 3618 2802 3623 2803
rect 4632 2803 4634 2807
rect 4634 2803 4637 2807
rect 4642 2803 4645 2807
rect 4645 2803 4647 2807
rect 4632 2802 4637 2803
rect 4642 2802 4647 2803
rect 1725 2797 1730 2802
rect 2365 2797 2370 2802
rect 3629 2797 3634 2802
rect 4525 2787 4530 2792
rect 5085 2787 5090 2792
rect 653 2777 658 2782
rect 2189 2777 2194 2782
rect 3933 2777 3938 2782
rect 4141 2767 4146 2772
rect 3005 2757 3010 2762
rect 3901 2757 3906 2762
rect 4525 2757 4530 2762
rect 701 2747 706 2752
rect 1629 2747 1634 2752
rect 1741 2747 1746 2752
rect 2381 2747 2386 2752
rect 3885 2747 3890 2752
rect 1981 2737 1986 2742
rect 3693 2737 3698 2742
rect 2749 2717 2754 2722
rect 3629 2717 3634 2722
rect 1533 2707 1538 2712
rect 1645 2707 1650 2712
rect 1805 2707 1810 2712
rect 2093 2707 2098 2712
rect 1048 2703 1050 2707
rect 1050 2703 1053 2707
rect 1058 2703 1061 2707
rect 1061 2703 1063 2707
rect 1048 2702 1053 2703
rect 1058 2702 1063 2703
rect 2072 2703 2074 2707
rect 2074 2703 2077 2707
rect 2082 2703 2085 2707
rect 2085 2703 2087 2707
rect 2072 2702 2077 2703
rect 2082 2702 2087 2703
rect 3096 2703 3098 2707
rect 3098 2703 3101 2707
rect 3106 2703 3109 2707
rect 3109 2703 3111 2707
rect 3096 2702 3101 2703
rect 3106 2702 3111 2703
rect 4112 2703 4114 2707
rect 4114 2703 4117 2707
rect 4122 2703 4125 2707
rect 4125 2703 4127 2707
rect 4112 2702 4117 2703
rect 4122 2702 4127 2703
rect 2157 2697 2162 2702
rect 2637 2687 2642 2692
rect 4397 2687 4402 2692
rect 845 2677 850 2682
rect 1293 2677 1298 2682
rect 1901 2677 1906 2682
rect 2381 2677 2386 2682
rect 2493 2677 2498 2682
rect 2205 2667 2210 2672
rect 1533 2657 1538 2662
rect 1581 2657 1586 2662
rect 1997 2657 2002 2662
rect 2397 2657 2402 2662
rect 5181 2657 5186 2662
rect 3981 2647 3986 2652
rect 1485 2637 1490 2642
rect 1661 2637 1666 2642
rect 3085 2637 3090 2642
rect 1741 2627 1746 2632
rect 2301 2627 2306 2632
rect 5101 2627 5106 2632
rect 1661 2617 1666 2622
rect 1949 2617 1954 2622
rect 2253 2617 2258 2622
rect 3133 2617 3138 2622
rect 1677 2607 1682 2612
rect 3373 2607 3378 2612
rect 536 2603 538 2607
rect 538 2603 541 2607
rect 546 2603 549 2607
rect 549 2603 551 2607
rect 536 2602 541 2603
rect 546 2602 551 2603
rect 1560 2603 1562 2607
rect 1562 2603 1565 2607
rect 1570 2603 1573 2607
rect 1573 2603 1575 2607
rect 1560 2602 1565 2603
rect 1570 2602 1575 2603
rect 2584 2603 2586 2607
rect 2586 2603 2589 2607
rect 2594 2603 2597 2607
rect 2597 2603 2599 2607
rect 2584 2602 2589 2603
rect 2594 2602 2599 2603
rect 3608 2603 3610 2607
rect 3610 2603 3613 2607
rect 3618 2603 3621 2607
rect 3621 2603 3623 2607
rect 3608 2602 3613 2603
rect 3618 2602 3623 2603
rect 4632 2603 4634 2607
rect 4634 2603 4637 2607
rect 4642 2603 4645 2607
rect 4645 2603 4647 2607
rect 4632 2602 4637 2603
rect 4642 2602 4647 2603
rect 493 2577 498 2582
rect 1981 2577 1986 2582
rect 2045 2577 2050 2582
rect 3837 2587 3842 2592
rect 4445 2587 4450 2592
rect 3133 2567 3138 2572
rect 3469 2567 3474 2572
rect 1149 2547 1154 2552
rect 1949 2557 1954 2562
rect 5101 2567 5106 2572
rect 5133 2557 5138 2562
rect 1213 2547 1218 2552
rect 1821 2537 1826 2542
rect 2397 2537 2402 2542
rect 5005 2537 5010 2542
rect 925 2527 930 2532
rect 3453 2527 3458 2532
rect 1693 2507 1698 2512
rect 1709 2507 1714 2512
rect 2109 2517 2114 2522
rect 2141 2517 2146 2522
rect 2349 2517 2354 2522
rect 1805 2507 1810 2512
rect 1048 2503 1050 2507
rect 1050 2503 1053 2507
rect 1058 2503 1061 2507
rect 1061 2503 1063 2507
rect 1048 2502 1053 2503
rect 1058 2502 1063 2503
rect 2072 2503 2074 2507
rect 2074 2503 2077 2507
rect 2082 2503 2085 2507
rect 2085 2503 2087 2507
rect 2072 2502 2077 2503
rect 2082 2502 2087 2503
rect 1069 2497 1074 2502
rect 1357 2497 1362 2502
rect 2045 2497 2050 2502
rect 2189 2497 2194 2502
rect 2333 2497 2338 2502
rect 3096 2503 3098 2507
rect 3098 2503 3101 2507
rect 3106 2503 3109 2507
rect 3109 2503 3111 2507
rect 3096 2502 3101 2503
rect 3106 2502 3111 2503
rect 2701 2487 2706 2492
rect 3117 2497 3122 2502
rect 4077 2497 4082 2502
rect 4112 2503 4114 2507
rect 4114 2503 4117 2507
rect 4122 2503 4125 2507
rect 4125 2503 4127 2507
rect 4112 2502 4117 2503
rect 4122 2502 4127 2503
rect 4077 2487 4082 2492
rect 1485 2477 1490 2482
rect 1549 2477 1554 2482
rect 2173 2477 2178 2482
rect 4205 2477 4210 2482
rect 1933 2467 1938 2472
rect 1997 2467 2002 2472
rect 2669 2467 2674 2472
rect 3117 2467 3122 2472
rect 589 2447 594 2452
rect 1533 2447 1538 2452
rect 1549 2447 1554 2452
rect 1597 2447 1602 2452
rect 1981 2457 1986 2462
rect 3005 2447 3010 2452
rect 3629 2447 3634 2452
rect 3933 2447 3938 2452
rect 1597 2437 1602 2442
rect 1613 2437 1618 2442
rect 1901 2437 1906 2442
rect 2045 2437 2050 2442
rect 2765 2437 2770 2442
rect 3117 2437 3122 2442
rect 3357 2437 3362 2442
rect 4365 2437 4370 2442
rect 1517 2427 1522 2432
rect 1533 2427 1538 2432
rect 1997 2427 2002 2432
rect 3469 2427 3474 2432
rect 3565 2427 3570 2432
rect 5149 2427 5154 2432
rect 1901 2417 1906 2422
rect 5149 2417 5154 2422
rect 1229 2407 1234 2412
rect 1309 2407 1314 2412
rect 2333 2407 2338 2412
rect 3565 2407 3570 2412
rect 536 2403 538 2407
rect 538 2403 541 2407
rect 546 2403 549 2407
rect 549 2403 551 2407
rect 536 2402 541 2403
rect 546 2402 551 2403
rect 1560 2403 1562 2407
rect 1562 2403 1565 2407
rect 1570 2403 1573 2407
rect 1573 2403 1575 2407
rect 1560 2402 1565 2403
rect 1570 2402 1575 2403
rect 2584 2403 2586 2407
rect 2586 2403 2589 2407
rect 2594 2403 2597 2407
rect 2597 2403 2599 2407
rect 2584 2402 2589 2403
rect 2594 2402 2599 2403
rect 3608 2403 3610 2407
rect 3610 2403 3613 2407
rect 3618 2403 3621 2407
rect 3621 2403 3623 2407
rect 3608 2402 3613 2403
rect 3618 2402 3623 2403
rect 4632 2403 4634 2407
rect 4634 2403 4637 2407
rect 4642 2403 4645 2407
rect 4645 2403 4647 2407
rect 4632 2402 4637 2403
rect 4642 2402 4647 2403
rect 1533 2397 1538 2402
rect 1597 2397 1602 2402
rect 1421 2387 1426 2392
rect 1725 2387 1730 2392
rect 2909 2397 2914 2402
rect 4429 2397 4434 2402
rect 2381 2387 2386 2392
rect 2941 2387 2946 2392
rect 3485 2387 3490 2392
rect 4573 2387 4578 2392
rect 1373 2377 1378 2382
rect 2093 2377 2098 2382
rect 2125 2377 2130 2382
rect 2141 2377 2146 2382
rect 2941 2377 2946 2382
rect 3117 2377 3122 2382
rect 4605 2377 4610 2382
rect 1597 2367 1602 2372
rect 2493 2367 2498 2372
rect 3597 2367 3602 2372
rect 3773 2367 3778 2372
rect 4349 2357 4354 2362
rect 1437 2347 1442 2352
rect 1517 2347 1522 2352
rect 2045 2347 2050 2352
rect 2509 2347 2514 2352
rect 3165 2347 3170 2352
rect 3341 2347 3346 2352
rect 3565 2347 3570 2352
rect 1357 2337 1362 2342
rect 1261 2327 1266 2332
rect 1453 2327 1458 2332
rect 1725 2327 1730 2332
rect 2205 2327 2210 2332
rect 2669 2327 2674 2332
rect 1389 2307 1394 2312
rect 2093 2307 2098 2312
rect 3293 2307 3298 2312
rect 3437 2307 3442 2312
rect 3581 2307 3586 2312
rect 1048 2303 1050 2307
rect 1050 2303 1053 2307
rect 1058 2303 1061 2307
rect 1061 2303 1063 2307
rect 1048 2302 1053 2303
rect 1058 2302 1063 2303
rect 2072 2303 2074 2307
rect 2074 2303 2077 2307
rect 2082 2303 2085 2307
rect 2085 2303 2087 2307
rect 2072 2302 2077 2303
rect 2082 2302 2087 2303
rect 3096 2303 3098 2307
rect 3098 2303 3101 2307
rect 3106 2303 3109 2307
rect 3109 2303 3111 2307
rect 3096 2302 3101 2303
rect 3106 2302 3111 2303
rect 4112 2303 4114 2307
rect 4114 2303 4117 2307
rect 4122 2303 4125 2307
rect 4125 2303 4127 2307
rect 4112 2302 4117 2303
rect 4122 2302 4127 2303
rect 4957 2307 4962 2312
rect 1197 2297 1202 2302
rect 1885 2297 1890 2302
rect 2157 2297 2162 2302
rect 2957 2297 2962 2302
rect 3229 2297 3234 2302
rect 2333 2287 2338 2292
rect 4413 2287 4418 2292
rect 2157 2277 2162 2282
rect 2189 2277 2194 2282
rect 5133 2277 5138 2282
rect 2093 2267 2098 2272
rect 2109 2267 2114 2272
rect 4541 2267 4546 2272
rect 4829 2267 4834 2272
rect 1645 2257 1650 2262
rect 1693 2257 1698 2262
rect 2813 2257 2818 2262
rect 4253 2257 4258 2262
rect 5085 2257 5090 2262
rect 1405 2247 1410 2252
rect 1821 2247 1826 2252
rect 1373 2237 1378 2242
rect 1917 2247 1922 2252
rect 1981 2247 1986 2252
rect 2125 2247 2130 2252
rect 2909 2247 2914 2252
rect 4285 2247 4290 2252
rect 4573 2247 4578 2252
rect 2029 2237 2034 2242
rect 2557 2237 2562 2242
rect 3773 2237 3778 2242
rect 3805 2237 3810 2242
rect 4237 2237 4242 2242
rect 909 2227 914 2232
rect 1773 2227 1778 2232
rect 2125 2227 2130 2232
rect 2317 2227 2322 2232
rect 3437 2227 3442 2232
rect 957 2207 962 2212
rect 1581 2207 1586 2212
rect 536 2203 538 2207
rect 538 2203 541 2207
rect 546 2203 549 2207
rect 549 2203 551 2207
rect 536 2202 541 2203
rect 546 2202 551 2203
rect 1560 2203 1562 2207
rect 1562 2203 1565 2207
rect 1570 2203 1573 2207
rect 1573 2203 1575 2207
rect 1560 2202 1565 2203
rect 1570 2202 1575 2203
rect 2584 2203 2586 2207
rect 2586 2203 2589 2207
rect 2594 2203 2597 2207
rect 2597 2203 2599 2207
rect 2584 2202 2589 2203
rect 2594 2202 2599 2203
rect 1837 2197 1842 2202
rect 2237 2197 2242 2202
rect 3309 2207 3314 2212
rect 3608 2203 3610 2207
rect 3610 2203 3613 2207
rect 3618 2203 3621 2207
rect 3621 2203 3623 2207
rect 3608 2202 3613 2203
rect 3618 2202 3623 2203
rect 4632 2203 4634 2207
rect 4634 2203 4637 2207
rect 4642 2203 4645 2207
rect 4645 2203 4647 2207
rect 4632 2202 4637 2203
rect 4642 2202 4647 2203
rect 829 2187 834 2192
rect 1581 2187 1586 2192
rect 2253 2187 2258 2192
rect 1629 2177 1634 2182
rect 2477 2177 2482 2182
rect 3037 2177 3042 2182
rect 3981 2178 3982 2182
rect 3982 2178 3986 2182
rect 3981 2177 3986 2178
rect 1901 2167 1906 2172
rect 1645 2157 1650 2162
rect 1789 2157 1794 2162
rect 2269 2157 2274 2162
rect 2813 2157 2818 2162
rect 3149 2157 3154 2162
rect 733 2137 738 2142
rect 2541 2147 2546 2152
rect 4749 2157 4754 2162
rect 4525 2147 4530 2152
rect 1213 2137 1218 2142
rect 2317 2137 2322 2142
rect 2429 2137 2434 2142
rect 2765 2137 2770 2142
rect 2845 2137 2850 2142
rect 3805 2137 3810 2142
rect 4589 2137 4594 2142
rect 4093 2127 4098 2132
rect 1709 2117 1714 2122
rect 1773 2117 1778 2122
rect 3405 2117 3410 2122
rect 4557 2117 4562 2122
rect 685 2107 690 2112
rect 2045 2107 2050 2112
rect 1048 2103 1050 2107
rect 1050 2103 1053 2107
rect 1058 2103 1061 2107
rect 1061 2103 1063 2107
rect 1048 2102 1053 2103
rect 1058 2102 1063 2103
rect 2072 2103 2074 2107
rect 2074 2103 2077 2107
rect 2082 2103 2085 2107
rect 2085 2103 2087 2107
rect 2072 2102 2077 2103
rect 2082 2102 2087 2103
rect 3096 2103 3098 2107
rect 3098 2103 3101 2107
rect 3106 2103 3109 2107
rect 3109 2103 3111 2107
rect 3096 2102 3101 2103
rect 3106 2102 3111 2103
rect 1709 2097 1714 2102
rect 4112 2103 4114 2107
rect 4114 2103 4117 2107
rect 4122 2103 4125 2107
rect 4125 2103 4127 2107
rect 4112 2102 4117 2103
rect 4122 2102 4127 2103
rect 1341 2087 1346 2092
rect 1805 2087 1810 2092
rect 1965 2087 1970 2092
rect 1037 2077 1042 2082
rect 1645 2077 1650 2082
rect 2797 2087 2802 2092
rect 4717 2087 4722 2092
rect 1581 2067 1586 2072
rect 3629 2077 3634 2082
rect 4093 2077 4098 2082
rect 4477 2077 4482 2082
rect 4509 2077 4514 2082
rect 4589 2077 4594 2082
rect 5085 2077 5090 2082
rect 2333 2067 2338 2072
rect 2797 2057 2802 2062
rect 3437 2067 3442 2072
rect 4669 2067 4674 2072
rect 4157 2057 4162 2062
rect 4189 2047 4194 2052
rect 653 2037 658 2042
rect 1853 2037 1858 2042
rect 2045 2037 2050 2042
rect 1069 2027 1074 2032
rect 1629 2027 1634 2032
rect 2109 2037 2114 2042
rect 3709 2037 3714 2042
rect 3933 2037 3938 2042
rect 5165 2037 5170 2042
rect 3181 2027 3186 2032
rect 1693 2017 1698 2022
rect 2509 2017 2514 2022
rect 2045 2007 2050 2012
rect 3533 2007 3538 2012
rect 3549 2007 3554 2012
rect 3581 2007 3586 2012
rect 3725 2007 3730 2012
rect 536 2003 538 2007
rect 538 2003 541 2007
rect 546 2003 549 2007
rect 549 2003 551 2007
rect 536 2002 541 2003
rect 546 2002 551 2003
rect 1560 2003 1562 2007
rect 1562 2003 1565 2007
rect 1570 2003 1573 2007
rect 1573 2003 1575 2007
rect 1560 2002 1565 2003
rect 1570 2002 1575 2003
rect 2584 2003 2586 2007
rect 2586 2003 2589 2007
rect 2594 2003 2597 2007
rect 2597 2003 2599 2007
rect 2584 2002 2589 2003
rect 2594 2002 2599 2003
rect 3608 2003 3610 2007
rect 3610 2003 3613 2007
rect 3618 2003 3621 2007
rect 3621 2003 3623 2007
rect 3608 2002 3613 2003
rect 3618 2002 3623 2003
rect 4632 2003 4634 2007
rect 4634 2003 4637 2007
rect 4642 2003 4645 2007
rect 4645 2003 4647 2007
rect 4632 2002 4637 2003
rect 4642 2002 4647 2003
rect 2141 1997 2146 2002
rect 2669 1997 2674 2002
rect 1341 1987 1346 1992
rect 4861 1987 4866 1992
rect 1149 1977 1154 1982
rect 1469 1977 1474 1982
rect 4221 1977 4226 1982
rect 1437 1967 1442 1972
rect 2109 1967 2114 1972
rect 1165 1947 1170 1952
rect 3421 1947 3426 1952
rect 3501 1947 3506 1952
rect 3869 1947 3874 1952
rect 861 1937 866 1942
rect 1501 1937 1506 1942
rect 2333 1937 2338 1942
rect 2493 1937 2498 1942
rect 4173 1937 4178 1942
rect 1405 1917 1410 1922
rect 2749 1917 2754 1922
rect 3309 1917 3314 1922
rect 4925 1917 4930 1922
rect 3053 1907 3058 1912
rect 3357 1907 3362 1912
rect 3517 1907 3522 1912
rect 3597 1907 3602 1912
rect 4061 1907 4066 1912
rect 1048 1903 1050 1907
rect 1050 1903 1053 1907
rect 1058 1903 1061 1907
rect 1061 1903 1063 1907
rect 1048 1902 1053 1903
rect 1058 1902 1063 1903
rect 2072 1903 2074 1907
rect 2074 1903 2077 1907
rect 2082 1903 2085 1907
rect 2085 1903 2087 1907
rect 2072 1902 2077 1903
rect 2082 1902 2087 1903
rect 3096 1903 3098 1907
rect 3098 1903 3101 1907
rect 3106 1903 3109 1907
rect 3109 1903 3111 1907
rect 3096 1902 3101 1903
rect 3106 1902 3111 1903
rect 4112 1903 4114 1907
rect 4114 1903 4117 1907
rect 4122 1903 4125 1907
rect 4125 1903 4127 1907
rect 4112 1902 4117 1903
rect 4122 1902 4127 1903
rect 1405 1897 1410 1902
rect 1981 1897 1986 1902
rect 2413 1897 2418 1902
rect 4349 1897 4354 1902
rect 3933 1887 3938 1892
rect 4301 1887 4306 1892
rect 1165 1867 1170 1872
rect 2685 1877 2690 1882
rect 3485 1877 3490 1882
rect 3757 1877 3762 1882
rect 1309 1867 1314 1872
rect 1613 1867 1618 1872
rect 1661 1867 1666 1872
rect 2189 1867 2194 1872
rect 1293 1857 1298 1862
rect 1613 1857 1618 1862
rect 3469 1857 3474 1862
rect 4301 1867 4306 1872
rect 5021 1867 5026 1872
rect 4477 1857 4482 1862
rect 1549 1847 1554 1852
rect 4557 1847 4562 1852
rect 1389 1837 1394 1842
rect 2013 1837 2018 1842
rect 3933 1837 3938 1842
rect 4749 1827 4754 1832
rect 1677 1817 1682 1822
rect 3453 1817 3458 1822
rect 1581 1807 1586 1812
rect 2429 1807 2434 1812
rect 536 1803 538 1807
rect 538 1803 541 1807
rect 546 1803 549 1807
rect 549 1803 551 1807
rect 536 1802 541 1803
rect 546 1802 551 1803
rect 1560 1803 1562 1807
rect 1562 1803 1565 1807
rect 1570 1803 1573 1807
rect 1573 1803 1575 1807
rect 1560 1802 1565 1803
rect 1570 1802 1575 1803
rect 2584 1803 2586 1807
rect 2586 1803 2589 1807
rect 2594 1803 2597 1807
rect 2597 1803 2599 1807
rect 2584 1802 2589 1803
rect 2594 1802 2599 1803
rect 3608 1803 3610 1807
rect 3610 1803 3613 1807
rect 3618 1803 3621 1807
rect 3621 1803 3623 1807
rect 3608 1802 3613 1803
rect 3618 1802 3623 1803
rect 4632 1803 4634 1807
rect 4634 1803 4637 1807
rect 4642 1803 4645 1807
rect 4645 1803 4647 1807
rect 4632 1802 4637 1803
rect 4642 1802 4647 1803
rect 1469 1797 1474 1802
rect 3389 1777 3394 1782
rect 3789 1777 3794 1782
rect 3117 1767 3122 1772
rect 3469 1767 3474 1772
rect 4813 1767 4818 1772
rect 3085 1757 3090 1762
rect 1197 1747 1202 1752
rect 2093 1747 2098 1752
rect 2541 1747 2546 1752
rect 4333 1747 4338 1752
rect 4429 1747 4434 1752
rect 1085 1737 1090 1742
rect 701 1727 706 1732
rect 3277 1727 3282 1732
rect 2157 1717 2162 1722
rect 2765 1717 2770 1722
rect 4621 1707 4626 1712
rect 5021 1707 5026 1712
rect 1048 1703 1050 1707
rect 1050 1703 1053 1707
rect 1058 1703 1061 1707
rect 1061 1703 1063 1707
rect 1048 1702 1053 1703
rect 1058 1702 1063 1703
rect 2072 1703 2074 1707
rect 2074 1703 2077 1707
rect 2082 1703 2085 1707
rect 2085 1703 2087 1707
rect 2072 1702 2077 1703
rect 2082 1702 2087 1703
rect 3096 1703 3098 1707
rect 3098 1703 3101 1707
rect 3106 1703 3109 1707
rect 3109 1703 3111 1707
rect 3096 1702 3101 1703
rect 3106 1702 3111 1703
rect 4112 1703 4114 1707
rect 4114 1703 4117 1707
rect 4122 1703 4125 1707
rect 4125 1703 4127 1707
rect 4112 1702 4117 1703
rect 4122 1702 4127 1703
rect 1741 1697 1746 1702
rect 2397 1697 2402 1702
rect 3117 1697 3122 1702
rect 4461 1697 4466 1702
rect 4861 1697 4866 1702
rect 781 1687 786 1692
rect 1277 1687 1282 1692
rect 957 1677 962 1682
rect 3997 1677 4002 1682
rect 4445 1677 4450 1682
rect 2285 1657 2290 1662
rect 3693 1667 3698 1672
rect 4397 1657 4402 1662
rect 669 1637 674 1642
rect 2205 1637 2210 1642
rect 2221 1637 2226 1642
rect 3149 1637 3154 1642
rect 1517 1627 1522 1632
rect 1805 1627 1810 1632
rect 2173 1627 2178 1632
rect 4765 1627 4770 1632
rect 2621 1607 2626 1612
rect 3325 1607 3330 1612
rect 3757 1607 3762 1612
rect 536 1603 538 1607
rect 538 1603 541 1607
rect 546 1603 549 1607
rect 549 1603 551 1607
rect 536 1602 541 1603
rect 546 1602 551 1603
rect 1560 1603 1562 1607
rect 1562 1603 1565 1607
rect 1570 1603 1573 1607
rect 1573 1603 1575 1607
rect 1560 1602 1565 1603
rect 1570 1602 1575 1603
rect 2584 1603 2586 1607
rect 2586 1603 2589 1607
rect 2594 1603 2597 1607
rect 2597 1603 2599 1607
rect 2584 1602 2589 1603
rect 2594 1602 2599 1603
rect 3608 1603 3610 1607
rect 3610 1603 3613 1607
rect 3618 1603 3621 1607
rect 3621 1603 3623 1607
rect 3608 1602 3613 1603
rect 3618 1602 3623 1603
rect 4632 1603 4634 1607
rect 4634 1603 4637 1607
rect 4642 1603 4645 1607
rect 4645 1603 4647 1607
rect 4632 1602 4637 1603
rect 4642 1602 4647 1603
rect 1597 1597 1602 1602
rect 1021 1587 1026 1592
rect 1693 1587 1698 1592
rect 2317 1587 2322 1592
rect 1069 1557 1074 1562
rect 2701 1567 2706 1572
rect 3789 1567 3794 1572
rect 3853 1567 3858 1572
rect 1949 1547 1954 1552
rect 2237 1537 2242 1542
rect 2829 1537 2834 1542
rect 3549 1537 3554 1542
rect 589 1527 594 1532
rect 3333 1527 3338 1532
rect 1048 1503 1050 1507
rect 1050 1503 1053 1507
rect 1058 1503 1061 1507
rect 1061 1503 1063 1507
rect 1048 1502 1053 1503
rect 1058 1502 1063 1503
rect 3773 1507 3778 1512
rect 2072 1503 2074 1507
rect 2074 1503 2077 1507
rect 2082 1503 2085 1507
rect 2085 1503 2087 1507
rect 2072 1502 2077 1503
rect 2082 1502 2087 1503
rect 3096 1503 3098 1507
rect 3098 1503 3101 1507
rect 3106 1503 3109 1507
rect 3109 1503 3111 1507
rect 3096 1502 3101 1503
rect 3106 1502 3111 1503
rect 4112 1503 4114 1507
rect 4114 1503 4117 1507
rect 4122 1503 4125 1507
rect 4125 1503 4127 1507
rect 4112 1502 4117 1503
rect 4122 1502 4127 1503
rect 1725 1497 1730 1502
rect 3229 1497 3234 1502
rect 3805 1497 3810 1502
rect 3901 1497 3906 1502
rect 5085 1497 5090 1502
rect 1373 1487 1378 1492
rect 1485 1487 1490 1492
rect 2189 1487 2194 1492
rect 2621 1487 2626 1492
rect 2061 1477 2066 1482
rect 3293 1477 3298 1482
rect 3805 1477 3810 1482
rect 4733 1477 4738 1482
rect 765 1467 770 1472
rect 1181 1467 1186 1472
rect 1997 1467 2002 1472
rect 3005 1467 3010 1472
rect 3085 1457 3090 1462
rect 381 1447 386 1452
rect 3677 1447 3682 1452
rect 813 1437 818 1442
rect 2125 1437 2130 1442
rect 2285 1437 2290 1442
rect 3821 1437 3826 1442
rect 3469 1417 3474 1422
rect 845 1407 850 1412
rect 536 1403 538 1407
rect 538 1403 541 1407
rect 546 1403 549 1407
rect 549 1403 551 1407
rect 536 1402 541 1403
rect 546 1402 551 1403
rect 1560 1403 1562 1407
rect 1562 1403 1565 1407
rect 1570 1403 1573 1407
rect 1573 1403 1575 1407
rect 1560 1402 1565 1403
rect 1570 1402 1575 1403
rect 2584 1403 2586 1407
rect 2586 1403 2589 1407
rect 2594 1403 2597 1407
rect 2597 1403 2599 1407
rect 2584 1402 2589 1403
rect 2594 1402 2599 1403
rect 3608 1403 3610 1407
rect 3610 1403 3613 1407
rect 3618 1403 3621 1407
rect 3621 1403 3623 1407
rect 3608 1402 3613 1403
rect 3618 1402 3623 1403
rect 4632 1403 4634 1407
rect 4634 1403 4637 1407
rect 4642 1403 4645 1407
rect 4645 1403 4647 1407
rect 4632 1402 4637 1403
rect 4642 1402 4647 1403
rect 3949 1387 3954 1392
rect 1229 1377 1234 1382
rect 1245 1377 1250 1382
rect 1149 1367 1154 1372
rect 3565 1367 3570 1372
rect 4077 1367 4082 1372
rect 4141 1367 4146 1372
rect 1133 1357 1138 1362
rect 1341 1357 1346 1362
rect 3597 1357 3602 1362
rect 3805 1357 3810 1362
rect 3869 1357 3874 1362
rect 717 1348 718 1352
rect 718 1348 722 1352
rect 717 1347 722 1348
rect 1613 1347 1618 1352
rect 925 1337 930 1342
rect 877 1327 882 1332
rect 1933 1317 1938 1322
rect 2797 1307 2802 1312
rect 1048 1303 1050 1307
rect 1050 1303 1053 1307
rect 1058 1303 1061 1307
rect 1061 1303 1063 1307
rect 1048 1302 1053 1303
rect 1058 1302 1063 1303
rect 2072 1303 2074 1307
rect 2074 1303 2077 1307
rect 2082 1303 2085 1307
rect 2085 1303 2087 1307
rect 2072 1302 2077 1303
rect 2082 1302 2087 1303
rect 3096 1303 3098 1307
rect 3098 1303 3101 1307
rect 3106 1303 3109 1307
rect 3109 1303 3111 1307
rect 3096 1302 3101 1303
rect 3106 1302 3111 1303
rect 4112 1303 4114 1307
rect 4114 1303 4117 1307
rect 4122 1303 4125 1307
rect 4125 1303 4127 1307
rect 4112 1302 4117 1303
rect 4122 1302 4127 1303
rect 3213 1297 3218 1302
rect 1165 1287 1170 1292
rect 2637 1277 2642 1282
rect 2701 1287 2706 1292
rect 3053 1277 3058 1282
rect 4573 1277 4578 1282
rect 589 1267 594 1272
rect 2093 1257 2098 1262
rect 3405 1247 3410 1252
rect 5021 1247 5026 1252
rect 1261 1237 1266 1242
rect 1197 1217 1202 1222
rect 3197 1217 3202 1222
rect 3485 1217 3490 1222
rect 4381 1217 4386 1222
rect 2941 1207 2946 1212
rect 3469 1207 3474 1212
rect 536 1203 538 1207
rect 538 1203 541 1207
rect 546 1203 549 1207
rect 549 1203 551 1207
rect 536 1202 541 1203
rect 546 1202 551 1203
rect 1560 1203 1562 1207
rect 1562 1203 1565 1207
rect 1570 1203 1573 1207
rect 1573 1203 1575 1207
rect 1560 1202 1565 1203
rect 1570 1202 1575 1203
rect 2584 1203 2586 1207
rect 2586 1203 2589 1207
rect 2594 1203 2597 1207
rect 2597 1203 2599 1207
rect 2584 1202 2589 1203
rect 2594 1202 2599 1203
rect 3608 1203 3610 1207
rect 3610 1203 3613 1207
rect 3618 1203 3621 1207
rect 3621 1203 3623 1207
rect 3608 1202 3613 1203
rect 3618 1202 3623 1203
rect 4632 1203 4634 1207
rect 4634 1203 4637 1207
rect 4642 1203 4645 1207
rect 4645 1203 4647 1207
rect 4632 1202 4637 1203
rect 4642 1202 4647 1203
rect 2253 1177 2258 1182
rect 2797 1177 2802 1182
rect 3709 1177 3714 1182
rect 4685 1177 4690 1182
rect 2093 1167 2098 1172
rect 4525 1167 4530 1172
rect 1389 1157 1394 1162
rect 3069 1157 3074 1162
rect 4093 1157 4098 1162
rect 477 1147 482 1152
rect 941 1147 946 1152
rect 749 1137 754 1142
rect 1949 1137 1954 1142
rect 3133 1137 3138 1142
rect 3405 1137 3410 1142
rect 2125 1127 2130 1132
rect 1213 1117 1218 1122
rect 3133 1117 3138 1122
rect 3405 1117 3410 1122
rect 1357 1107 1362 1112
rect 2845 1107 2850 1112
rect 1048 1103 1050 1107
rect 1050 1103 1053 1107
rect 1058 1103 1061 1107
rect 1061 1103 1063 1107
rect 1048 1102 1053 1103
rect 1058 1102 1063 1103
rect 2072 1103 2074 1107
rect 2074 1103 2077 1107
rect 2082 1103 2085 1107
rect 2085 1103 2087 1107
rect 2072 1102 2077 1103
rect 2082 1102 2087 1103
rect 3096 1103 3098 1107
rect 3098 1103 3101 1107
rect 3106 1103 3109 1107
rect 3109 1103 3111 1107
rect 3096 1102 3101 1103
rect 3106 1102 3111 1103
rect 4112 1103 4114 1107
rect 4114 1103 4117 1107
rect 4122 1103 4125 1107
rect 4125 1103 4127 1107
rect 4112 1102 4117 1103
rect 4122 1102 4127 1103
rect 2253 1097 2258 1102
rect 3661 1097 3666 1102
rect 3853 1057 3858 1062
rect 2605 1037 2610 1042
rect 4829 1047 4834 1052
rect 1773 1017 1778 1022
rect 3197 1017 3202 1022
rect 4621 1017 4626 1022
rect 536 1003 538 1007
rect 538 1003 541 1007
rect 546 1003 549 1007
rect 549 1003 551 1007
rect 536 1002 541 1003
rect 546 1002 551 1003
rect 1560 1003 1562 1007
rect 1562 1003 1565 1007
rect 1570 1003 1573 1007
rect 1573 1003 1575 1007
rect 1560 1002 1565 1003
rect 1570 1002 1575 1003
rect 2584 1003 2586 1007
rect 2586 1003 2589 1007
rect 2594 1003 2597 1007
rect 2597 1003 2599 1007
rect 2584 1002 2589 1003
rect 2594 1002 2599 1003
rect 3608 1003 3610 1007
rect 3610 1003 3613 1007
rect 3618 1003 3621 1007
rect 3621 1003 3623 1007
rect 3608 1002 3613 1003
rect 3618 1002 3623 1003
rect 4632 1003 4634 1007
rect 4634 1003 4637 1007
rect 4642 1003 4645 1007
rect 4645 1003 4647 1007
rect 4632 1002 4637 1003
rect 4642 1002 4647 1003
rect 2349 997 2354 1002
rect 2605 997 2610 1002
rect 813 957 818 962
rect 3885 947 3890 952
rect 4333 947 4338 952
rect 3309 937 3314 942
rect 3565 927 3570 932
rect 5149 927 5154 932
rect 2205 917 2210 922
rect 3965 907 3970 912
rect 1048 903 1050 907
rect 1050 903 1053 907
rect 1058 903 1061 907
rect 1061 903 1063 907
rect 1048 902 1053 903
rect 1058 902 1063 903
rect 2072 903 2074 907
rect 2074 903 2077 907
rect 2082 903 2085 907
rect 2085 903 2087 907
rect 2072 902 2077 903
rect 2082 902 2087 903
rect 3096 903 3098 907
rect 3098 903 3101 907
rect 3106 903 3109 907
rect 3109 903 3111 907
rect 3096 902 3101 903
rect 3106 902 3111 903
rect 4112 903 4114 907
rect 4114 903 4117 907
rect 4122 903 4125 907
rect 4125 903 4127 907
rect 4112 902 4117 903
rect 4122 902 4127 903
rect 2093 887 2098 892
rect 4973 887 4978 892
rect 957 877 962 882
rect 2957 877 2962 882
rect 1949 867 1954 872
rect 1293 857 1298 862
rect 2301 857 2306 862
rect 3341 857 3346 862
rect 589 847 594 852
rect 1933 847 1938 852
rect 2333 847 2338 852
rect 5181 847 5186 852
rect 3581 837 3586 842
rect 4237 837 4242 842
rect 536 803 538 807
rect 538 803 541 807
rect 546 803 549 807
rect 549 803 551 807
rect 536 802 541 803
rect 546 802 551 803
rect 1560 803 1562 807
rect 1562 803 1565 807
rect 1570 803 1573 807
rect 1573 803 1575 807
rect 1560 802 1565 803
rect 1570 802 1575 803
rect 2584 803 2586 807
rect 2586 803 2589 807
rect 2594 803 2597 807
rect 2597 803 2599 807
rect 2584 802 2589 803
rect 2594 802 2599 803
rect 3608 803 3610 807
rect 3610 803 3613 807
rect 3618 803 3621 807
rect 3621 803 3623 807
rect 3608 802 3613 803
rect 3618 802 3623 803
rect 4632 803 4634 807
rect 4634 803 4637 807
rect 4642 803 4645 807
rect 4645 803 4647 807
rect 4632 802 4637 803
rect 4642 802 4647 803
rect 2573 797 2578 802
rect 2605 797 2610 802
rect 3277 797 3282 802
rect 2829 787 2834 792
rect 2653 777 2658 782
rect 925 767 930 772
rect 2605 767 2610 772
rect 2845 767 2850 772
rect 2573 757 2578 762
rect 3565 767 3570 772
rect 4557 767 4562 772
rect 3309 757 3314 762
rect 3741 747 3746 752
rect 4301 747 4306 752
rect 4413 747 4418 752
rect 3757 737 3762 742
rect 4029 727 4034 732
rect 1048 703 1050 707
rect 1050 703 1053 707
rect 1058 703 1061 707
rect 1061 703 1063 707
rect 1048 702 1053 703
rect 1058 702 1063 703
rect 2072 703 2074 707
rect 2074 703 2077 707
rect 2082 703 2085 707
rect 2085 703 2087 707
rect 2072 702 2077 703
rect 2082 702 2087 703
rect 3096 703 3098 707
rect 3098 703 3101 707
rect 3106 703 3109 707
rect 3109 703 3111 707
rect 3096 702 3101 703
rect 3106 702 3111 703
rect 4112 703 4114 707
rect 4114 703 4117 707
rect 4122 703 4125 707
rect 4125 703 4127 707
rect 4112 702 4117 703
rect 4122 702 4127 703
rect 1245 677 1250 682
rect 3469 657 3474 662
rect 4749 657 4754 662
rect 2109 647 2114 652
rect 1757 637 1762 642
rect 4621 627 4626 632
rect 536 603 538 607
rect 538 603 541 607
rect 546 603 549 607
rect 549 603 551 607
rect 536 602 541 603
rect 546 602 551 603
rect 1560 603 1562 607
rect 1562 603 1565 607
rect 1570 603 1573 607
rect 1573 603 1575 607
rect 1560 602 1565 603
rect 1570 602 1575 603
rect 2584 603 2586 607
rect 2586 603 2589 607
rect 2594 603 2597 607
rect 2597 603 2599 607
rect 2584 602 2589 603
rect 2594 602 2599 603
rect 3608 603 3610 607
rect 3610 603 3613 607
rect 3618 603 3621 607
rect 3621 603 3623 607
rect 3608 602 3613 603
rect 3618 602 3623 603
rect 4632 603 4634 607
rect 4634 603 4637 607
rect 4642 603 4645 607
rect 4645 603 4647 607
rect 4632 602 4637 603
rect 4642 602 4647 603
rect 1805 587 1810 592
rect 941 567 946 572
rect 3501 547 3506 552
rect 1469 527 1474 532
rect 4477 527 4482 532
rect 1048 503 1050 507
rect 1050 503 1053 507
rect 1058 503 1061 507
rect 1061 503 1063 507
rect 1048 502 1053 503
rect 1058 502 1063 503
rect 2072 503 2074 507
rect 2074 503 2077 507
rect 2082 503 2085 507
rect 2085 503 2087 507
rect 2072 502 2077 503
rect 2082 502 2087 503
rect 3096 503 3098 507
rect 3098 503 3101 507
rect 3106 503 3109 507
rect 3109 503 3111 507
rect 3096 502 3101 503
rect 3106 502 3111 503
rect 4112 503 4114 507
rect 4114 503 4117 507
rect 4122 503 4125 507
rect 4125 503 4127 507
rect 4112 502 4117 503
rect 4122 502 4127 503
rect 1517 457 1522 462
rect 4029 447 4034 452
rect 536 403 538 407
rect 538 403 541 407
rect 546 403 549 407
rect 549 403 551 407
rect 536 402 541 403
rect 546 402 551 403
rect 1560 403 1562 407
rect 1562 403 1565 407
rect 1570 403 1573 407
rect 1573 403 1575 407
rect 1560 402 1565 403
rect 1570 402 1575 403
rect 2584 403 2586 407
rect 2586 403 2589 407
rect 2594 403 2597 407
rect 2597 403 2599 407
rect 2584 402 2589 403
rect 2594 402 2599 403
rect 3608 403 3610 407
rect 3610 403 3613 407
rect 3618 403 3621 407
rect 3621 403 3623 407
rect 3608 402 3613 403
rect 3618 402 3623 403
rect 4632 403 4634 407
rect 4634 403 4637 407
rect 4642 403 4645 407
rect 4645 403 4647 407
rect 4632 402 4637 403
rect 4642 402 4647 403
rect 1048 303 1050 307
rect 1050 303 1053 307
rect 1058 303 1061 307
rect 1061 303 1063 307
rect 1048 302 1053 303
rect 1058 302 1063 303
rect 2072 303 2074 307
rect 2074 303 2077 307
rect 2082 303 2085 307
rect 2085 303 2087 307
rect 2072 302 2077 303
rect 2082 302 2087 303
rect 3096 303 3098 307
rect 3098 303 3101 307
rect 3106 303 3109 307
rect 3109 303 3111 307
rect 3096 302 3101 303
rect 3106 302 3111 303
rect 4112 303 4114 307
rect 4114 303 4117 307
rect 4122 303 4125 307
rect 4125 303 4127 307
rect 4112 302 4117 303
rect 4122 302 4127 303
rect 5117 287 5122 292
rect 1325 277 1330 282
rect 4861 267 4866 272
rect 3805 257 3810 262
rect 536 203 538 207
rect 538 203 541 207
rect 546 203 549 207
rect 549 203 551 207
rect 536 202 541 203
rect 546 202 551 203
rect 1560 203 1562 207
rect 1562 203 1565 207
rect 1570 203 1573 207
rect 1573 203 1575 207
rect 1560 202 1565 203
rect 1570 202 1575 203
rect 2584 203 2586 207
rect 2586 203 2589 207
rect 2594 203 2597 207
rect 2597 203 2599 207
rect 2584 202 2589 203
rect 2594 202 2599 203
rect 3608 203 3610 207
rect 3610 203 3613 207
rect 3618 203 3621 207
rect 3621 203 3623 207
rect 3608 202 3613 203
rect 3618 202 3623 203
rect 4632 203 4634 207
rect 4634 203 4637 207
rect 4642 203 4645 207
rect 4645 203 4647 207
rect 4632 202 4637 203
rect 4642 202 4647 203
rect 5101 187 5106 192
rect 3485 157 3490 162
rect 2509 147 2514 152
rect 4669 137 4674 142
rect 4605 107 4610 112
rect 1048 103 1050 107
rect 1050 103 1053 107
rect 1058 103 1061 107
rect 1061 103 1063 107
rect 1048 102 1053 103
rect 1058 102 1063 103
rect 2072 103 2074 107
rect 2074 103 2077 107
rect 2082 103 2085 107
rect 2085 103 2087 107
rect 2072 102 2077 103
rect 2082 102 2087 103
rect 3096 103 3098 107
rect 3098 103 3101 107
rect 3106 103 3109 107
rect 3109 103 3111 107
rect 3096 102 3101 103
rect 3106 102 3111 103
rect 4112 103 4114 107
rect 4114 103 4117 107
rect 4122 103 4125 107
rect 4125 103 4127 107
rect 4112 102 4117 103
rect 4122 102 4127 103
rect 5005 87 5010 92
rect 4957 77 4962 82
rect 4541 57 4546 62
rect 4717 57 4722 62
rect 4589 47 4594 52
rect 4813 47 4818 52
rect 536 3 538 7
rect 538 3 541 7
rect 546 3 549 7
rect 549 3 551 7
rect 536 2 541 3
rect 546 2 551 3
rect 1560 3 1562 7
rect 1562 3 1565 7
rect 1570 3 1573 7
rect 1573 3 1575 7
rect 1560 2 1565 3
rect 1570 2 1575 3
rect 2584 3 2586 7
rect 2586 3 2589 7
rect 2594 3 2597 7
rect 2597 3 2599 7
rect 2584 2 2589 3
rect 2594 2 2599 3
rect 3608 3 3610 7
rect 3610 3 3613 7
rect 3618 3 3621 7
rect 3621 3 3623 7
rect 3608 2 3613 3
rect 3618 2 3623 3
rect 4632 3 4634 7
rect 4634 3 4637 7
rect 4642 3 4645 7
rect 4645 3 4647 7
rect 4632 2 4637 3
rect 4642 2 4647 3
<< metal6 >>
rect 536 4807 552 4930
rect 541 4802 546 4807
rect 551 4802 552 4807
rect 536 4607 552 4802
rect 541 4602 546 4607
rect 551 4602 552 4607
rect 536 4407 552 4602
rect 1048 4907 1064 4930
rect 1053 4902 1058 4907
rect 1063 4902 1064 4907
rect 1048 4707 1064 4902
rect 1053 4702 1058 4707
rect 1063 4702 1064 4707
rect 541 4402 546 4407
rect 551 4402 552 4407
rect 381 1452 386 3747
rect 477 1152 482 3497
rect 493 2582 498 4347
rect 536 4207 552 4402
rect 541 4202 546 4207
rect 551 4202 552 4207
rect 536 4007 552 4202
rect 541 4002 546 4007
rect 551 4002 552 4007
rect 536 3807 552 4002
rect 541 3802 546 3807
rect 551 3802 552 3807
rect 536 3607 552 3802
rect 541 3602 546 3607
rect 551 3602 552 3607
rect 536 3407 552 3602
rect 541 3402 546 3407
rect 551 3402 552 3407
rect 536 3207 552 3402
rect 541 3202 546 3207
rect 551 3202 552 3207
rect 536 3007 552 3202
rect 541 3002 546 3007
rect 551 3002 552 3007
rect 536 2807 552 3002
rect 541 2802 546 2807
rect 551 2802 552 2807
rect 536 2607 552 2802
rect 541 2602 546 2607
rect 551 2602 552 2607
rect 536 2407 552 2602
rect 541 2402 546 2407
rect 551 2402 552 2407
rect 536 2207 552 2402
rect 541 2202 546 2207
rect 551 2202 552 2207
rect 536 2007 552 2202
rect 541 2002 546 2007
rect 551 2002 552 2007
rect 536 1807 552 2002
rect 541 1802 546 1807
rect 551 1802 552 1807
rect 536 1607 552 1802
rect 541 1602 546 1607
rect 551 1602 552 1607
rect 536 1407 552 1602
rect 589 1532 594 2447
rect 653 2042 658 2777
rect 669 1642 674 3687
rect 685 3402 690 3447
rect 685 2112 690 3397
rect 701 1732 706 2747
rect 541 1402 546 1407
rect 551 1402 552 1407
rect 536 1207 552 1402
rect 717 1352 722 3147
rect 733 2142 738 3407
rect 541 1202 546 1207
rect 551 1202 552 1207
rect 536 1007 552 1202
rect 541 1002 546 1007
rect 551 1002 552 1007
rect 536 807 552 1002
rect 589 852 594 1267
rect 749 1142 754 4537
rect 1048 4507 1064 4702
rect 1053 4502 1058 4507
rect 1063 4502 1064 4507
rect 765 1472 770 3477
rect 781 1692 786 4317
rect 1048 4307 1064 4502
rect 1053 4302 1058 4307
rect 1063 4302 1064 4307
rect 1048 4107 1064 4302
rect 1560 4807 1576 4930
rect 1565 4802 1570 4807
rect 1575 4802 1576 4807
rect 1560 4607 1576 4802
rect 2072 4907 2088 4930
rect 2077 4902 2082 4907
rect 2087 4902 2088 4907
rect 2072 4707 2088 4902
rect 2077 4702 2082 4707
rect 2087 4702 2088 4707
rect 1565 4602 1570 4607
rect 1575 4602 1576 4607
rect 1560 4407 1576 4602
rect 1565 4402 1570 4407
rect 1575 4402 1576 4407
rect 1560 4207 1576 4402
rect 1565 4202 1570 4207
rect 1575 4202 1576 4207
rect 1053 4102 1058 4107
rect 1063 4102 1064 4107
rect 1048 3907 1064 4102
rect 1053 3902 1058 3907
rect 1063 3902 1064 3907
rect 797 2952 802 3867
rect 829 2192 834 3177
rect 813 962 818 1437
rect 845 1412 850 2677
rect 861 1942 866 2947
rect 877 1332 882 3417
rect 909 2232 914 3887
rect 1048 3707 1064 3902
rect 1053 3702 1058 3707
rect 1063 3702 1064 3707
rect 941 3287 949 3292
rect 925 2532 930 3257
rect 941 3032 946 3287
rect 541 802 546 807
rect 551 802 552 807
rect 536 607 552 802
rect 925 772 930 1337
rect 941 1152 946 2977
rect 957 2212 962 3237
rect 1037 3022 1042 3697
rect 1048 3507 1064 3702
rect 1053 3502 1058 3507
rect 1063 3502 1064 3507
rect 1048 3307 1064 3502
rect 1053 3302 1058 3307
rect 1063 3302 1064 3307
rect 1048 3107 1064 3302
rect 1053 3102 1058 3107
rect 1063 3102 1064 3107
rect 541 602 546 607
rect 551 602 552 607
rect 536 407 552 602
rect 941 572 946 1147
rect 957 882 962 1677
rect 1021 1592 1026 2867
rect 1037 2082 1042 2937
rect 1048 2907 1064 3102
rect 1053 2902 1058 2907
rect 1063 2902 1064 2907
rect 1048 2707 1064 2902
rect 1053 2702 1058 2707
rect 1063 2702 1064 2707
rect 1048 2507 1064 2702
rect 1053 2502 1058 2507
rect 1063 2502 1064 2507
rect 1048 2307 1064 2502
rect 1069 3182 1074 3457
rect 1069 2502 1074 3177
rect 1053 2302 1058 2307
rect 1063 2302 1064 2307
rect 1048 2107 1064 2302
rect 1053 2102 1058 2107
rect 1063 2102 1064 2107
rect 1048 1907 1064 2102
rect 1053 1902 1058 1907
rect 1063 1902 1064 1907
rect 1048 1707 1064 1902
rect 1053 1702 1058 1707
rect 1063 1702 1064 1707
rect 1048 1507 1064 1702
rect 1069 1562 1074 2027
rect 1085 1742 1090 3637
rect 1053 1502 1058 1507
rect 1063 1502 1064 1507
rect 1048 1307 1064 1502
rect 1133 1362 1138 3407
rect 1149 2552 1154 3207
rect 1149 1372 1154 1977
rect 1165 1952 1170 3137
rect 1053 1302 1058 1307
rect 1063 1302 1064 1307
rect 1048 1107 1064 1302
rect 1165 1292 1170 1867
rect 1181 1472 1186 2907
rect 1197 2302 1202 3337
rect 1261 3042 1266 4117
rect 1560 4007 1576 4202
rect 1565 4002 1570 4007
rect 1575 4002 1576 4007
rect 1213 3022 1218 3037
rect 1213 2552 1218 2987
rect 1197 1222 1202 1747
rect 1213 1122 1218 2137
rect 1229 1382 1234 2407
rect 1053 1102 1058 1107
rect 1063 1102 1064 1107
rect 1048 907 1064 1102
rect 1053 902 1058 907
rect 1063 902 1064 907
rect 1048 707 1064 902
rect 1053 702 1058 707
rect 1063 702 1064 707
rect 541 402 546 407
rect 551 402 552 407
rect 536 207 552 402
rect 541 202 546 207
rect 551 202 552 207
rect 536 7 552 202
rect 541 2 546 7
rect 551 2 552 7
rect 536 -30 552 2
rect 1048 507 1064 702
rect 1245 682 1250 1377
rect 1261 1242 1266 2327
rect 1277 1692 1282 3427
rect 1293 2682 1298 3157
rect 1309 2932 1314 3597
rect 1357 3312 1362 3417
rect 1309 1872 1314 2407
rect 1293 862 1298 1857
rect 1053 502 1058 507
rect 1063 502 1064 507
rect 1048 307 1064 502
rect 1053 302 1058 307
rect 1063 302 1064 307
rect 1048 107 1064 302
rect 1325 282 1330 3207
rect 1341 2092 1346 3227
rect 1357 2502 1362 3027
rect 1373 2382 1378 2877
rect 1341 1362 1346 1987
rect 1357 1112 1362 2337
rect 1389 2312 1394 3167
rect 1405 2252 1410 3717
rect 1421 2392 1426 3127
rect 1437 2842 1442 3517
rect 1453 3472 1458 3517
rect 1373 1492 1378 2237
rect 1437 1972 1442 2347
rect 1453 2332 1458 3327
rect 1469 1982 1474 3497
rect 1485 3092 1490 3227
rect 1485 2642 1490 3087
rect 1405 1902 1410 1917
rect 1389 1162 1394 1837
rect 1469 532 1474 1797
rect 1485 1492 1490 2477
rect 1501 1942 1506 2927
rect 1533 2712 1538 3147
rect 1533 2452 1538 2657
rect 1549 2482 1554 3847
rect 1560 3807 1576 4002
rect 1565 3802 1570 3807
rect 1575 3802 1576 3807
rect 1560 3607 1576 3802
rect 1597 3702 1602 4637
rect 1565 3602 1570 3607
rect 1575 3602 1576 3607
rect 1560 3407 1576 3602
rect 1565 3402 1570 3407
rect 1575 3402 1576 3407
rect 1560 3207 1576 3402
rect 1565 3202 1570 3207
rect 1575 3202 1576 3207
rect 1560 3007 1576 3202
rect 1565 3002 1570 3007
rect 1575 3002 1576 3007
rect 1560 2807 1576 3002
rect 1565 2802 1570 2807
rect 1575 2802 1576 2807
rect 1560 2607 1576 2802
rect 1581 2662 1586 3417
rect 1629 3352 1634 4527
rect 2072 4507 2088 4702
rect 2077 4502 2082 4507
rect 2087 4502 2088 4507
rect 1661 3542 1666 4447
rect 1629 3232 1634 3277
rect 1565 2602 1570 2607
rect 1575 2602 1576 2607
rect 1517 2352 1522 2427
rect 1533 2402 1538 2427
rect 1549 1852 1554 2447
rect 1560 2407 1576 2602
rect 1597 2452 1602 3057
rect 1645 2902 1650 3317
rect 1629 2752 1634 2807
rect 1565 2402 1570 2407
rect 1575 2402 1576 2407
rect 1560 2207 1576 2402
rect 1597 2402 1602 2437
rect 1565 2202 1570 2207
rect 1575 2202 1576 2207
rect 1560 2007 1576 2202
rect 1581 2192 1586 2207
rect 1565 2002 1570 2007
rect 1575 2002 1576 2007
rect 1560 1807 1576 2002
rect 1581 1812 1586 2067
rect 1565 1802 1570 1807
rect 1575 1802 1576 1807
rect 1517 462 1522 1627
rect 1560 1607 1576 1802
rect 1565 1602 1570 1607
rect 1575 1602 1576 1607
rect 1560 1407 1576 1602
rect 1597 1602 1602 2367
rect 1613 1872 1618 2437
rect 1645 2262 1650 2707
rect 1661 2642 1666 3537
rect 1709 3212 1714 3697
rect 1725 3042 1730 3767
rect 1629 2032 1634 2177
rect 1645 2082 1650 2157
rect 1661 1872 1666 2617
rect 1565 1402 1570 1407
rect 1575 1402 1576 1407
rect 1560 1207 1576 1402
rect 1613 1352 1618 1857
rect 1677 1822 1682 2607
rect 1709 2512 1714 2977
rect 1693 2262 1698 2507
rect 1725 2392 1730 2797
rect 1741 2752 1746 3577
rect 1709 2102 1714 2117
rect 1693 1592 1698 2017
rect 1725 1502 1730 2327
rect 1741 1702 1746 2627
rect 1565 1202 1570 1207
rect 1575 1202 1576 1207
rect 1560 1007 1576 1202
rect 1565 1002 1570 1007
rect 1575 1002 1576 1007
rect 1560 807 1576 1002
rect 1565 802 1570 807
rect 1575 802 1576 807
rect 1560 607 1576 802
rect 1757 642 1762 3297
rect 1773 2232 1778 3157
rect 1789 2162 1794 3417
rect 1805 2712 1810 4387
rect 2072 4307 2088 4502
rect 2077 4302 2082 4307
rect 2087 4302 2088 4307
rect 2072 4107 2088 4302
rect 2077 4102 2082 4107
rect 2087 4102 2088 4107
rect 1821 3492 1826 3647
rect 1773 1022 1778 2117
rect 1805 2092 1810 2507
rect 1821 2252 1826 2537
rect 1837 2202 1842 3117
rect 1853 2042 1858 3627
rect 1885 2302 1890 2927
rect 1901 2922 1906 2947
rect 1901 2442 1906 2677
rect 1901 2172 1906 2417
rect 1917 2252 1922 3437
rect 1933 3212 1938 3737
rect 1949 2622 1954 3727
rect 2029 3362 2034 3737
rect 2061 3722 2066 3907
rect 2072 3907 2088 4102
rect 2077 3902 2082 3907
rect 2087 3902 2088 3907
rect 2072 3707 2088 3902
rect 2077 3702 2082 3707
rect 2087 3702 2088 3707
rect 2072 3507 2088 3702
rect 2093 3582 2098 3597
rect 2077 3502 2082 3507
rect 2087 3502 2088 3507
rect 1565 602 1570 607
rect 1575 602 1576 607
rect 1560 407 1576 602
rect 1805 592 1810 1627
rect 1933 1322 1938 2467
rect 1949 1552 1954 2557
rect 1965 2092 1970 2997
rect 1981 2742 1986 3017
rect 1981 2462 1986 2577
rect 1997 2472 2002 2657
rect 1981 1902 1986 2247
rect 1997 1472 2002 2427
rect 2013 1842 2018 3237
rect 2029 2242 2034 3327
rect 2072 3307 2088 3502
rect 2077 3302 2082 3307
rect 2087 3302 2088 3307
rect 2045 2582 2050 3017
rect 2045 2442 2050 2497
rect 2045 2112 2050 2347
rect 2045 2012 2050 2037
rect 2061 1482 2066 3137
rect 2072 3107 2088 3302
rect 2125 3282 2130 3327
rect 2077 3102 2082 3107
rect 2087 3102 2088 3107
rect 2072 2907 2088 3102
rect 2077 2902 2082 2907
rect 2087 2902 2088 2907
rect 2072 2707 2088 2902
rect 2077 2702 2082 2707
rect 2087 2702 2088 2707
rect 2072 2507 2088 2702
rect 2077 2502 2082 2507
rect 2087 2502 2088 2507
rect 2072 2307 2088 2502
rect 2093 2382 2098 2707
rect 2109 2522 2114 3137
rect 2125 2852 2130 2907
rect 2125 2382 2130 2847
rect 2141 2522 2146 3157
rect 2157 2882 2162 3787
rect 2173 3502 2178 4167
rect 2189 2782 2194 4307
rect 2221 3012 2226 3707
rect 2317 3682 2322 3697
rect 2285 3122 2290 3607
rect 2077 2302 2082 2307
rect 2087 2302 2088 2307
rect 2072 2107 2088 2302
rect 2093 2272 2098 2307
rect 2077 2102 2082 2107
rect 2087 2102 2088 2107
rect 2072 1907 2088 2102
rect 2109 2042 2114 2267
rect 2125 2232 2130 2247
rect 2141 2002 2146 2377
rect 2157 2302 2162 2697
rect 2077 1902 2082 1907
rect 2087 1902 2088 1907
rect 2072 1707 2088 1902
rect 2077 1702 2082 1707
rect 2087 1702 2088 1707
rect 2072 1507 2088 1702
rect 2077 1502 2082 1507
rect 2087 1502 2088 1507
rect 1933 852 1938 1317
rect 2072 1307 2088 1502
rect 2077 1302 2082 1307
rect 2087 1302 2088 1307
rect 1949 872 1954 1137
rect 2072 1107 2088 1302
rect 2093 1262 2098 1747
rect 2077 1102 2082 1107
rect 2087 1102 2088 1107
rect 2072 907 2088 1102
rect 2077 902 2082 907
rect 2087 902 2088 907
rect 2072 707 2088 902
rect 2093 892 2098 1167
rect 2077 702 2082 707
rect 2087 702 2088 707
rect 1565 402 1570 407
rect 1575 402 1576 407
rect 1053 102 1058 107
rect 1063 102 1064 107
rect 1048 -30 1064 102
rect 1560 207 1576 402
rect 1565 202 1570 207
rect 1575 202 1576 207
rect 1560 7 1576 202
rect 1565 2 1570 7
rect 1575 2 1576 7
rect 1560 -30 1576 2
rect 2072 507 2088 702
rect 2109 652 2114 1967
rect 2157 1722 2162 2277
rect 2173 1632 2178 2477
rect 2189 2282 2194 2497
rect 2205 2332 2210 2667
rect 2189 1492 2194 1867
rect 2221 1642 2226 3007
rect 2125 1132 2130 1437
rect 2205 922 2210 1637
rect 2237 1542 2242 2197
rect 2253 2192 2258 2617
rect 2269 2162 2274 3087
rect 2301 3062 2306 3097
rect 2285 1442 2290 1657
rect 2253 1102 2258 1177
rect 2301 862 2306 2627
rect 2317 2232 2322 2887
rect 2333 2502 2338 4427
rect 2365 4032 2370 4057
rect 2365 2802 2370 4027
rect 2381 3462 2386 4857
rect 2584 4807 2600 4930
rect 2589 4802 2594 4807
rect 2599 4802 2600 4807
rect 2584 4607 2600 4802
rect 2589 4602 2594 4607
rect 2599 4602 2600 4607
rect 2584 4407 2600 4602
rect 3096 4907 3112 4930
rect 3101 4902 3106 4907
rect 3111 4902 3112 4907
rect 3096 4707 3112 4902
rect 3101 4702 3106 4707
rect 3111 4702 3112 4707
rect 3096 4507 3112 4702
rect 3608 4807 3624 4930
rect 3613 4802 3618 4807
rect 3623 4802 3624 4807
rect 3608 4607 3624 4802
rect 3613 4602 3618 4607
rect 3623 4602 3624 4607
rect 3101 4502 3106 4507
rect 3111 4502 3112 4507
rect 2589 4402 2594 4407
rect 2599 4402 2600 4407
rect 2477 4232 2482 4247
rect 2397 3732 2402 3887
rect 2381 2682 2386 2747
rect 2333 2292 2338 2407
rect 2317 1592 2322 2137
rect 2333 2072 2338 2287
rect 2333 852 2338 1937
rect 2349 1002 2354 2517
rect 2381 2392 2386 2677
rect 2397 2662 2402 3197
rect 2397 1702 2402 2537
rect 2413 1902 2418 3817
rect 2477 2182 2482 3607
rect 2493 2682 2498 3957
rect 2541 3472 2546 3497
rect 2541 2882 2546 3467
rect 2557 3312 2562 4257
rect 2429 1812 2434 2137
rect 2493 1942 2498 2367
rect 2509 2352 2514 2807
rect 2557 2242 2562 3307
rect 2584 4207 2600 4402
rect 2733 4372 2738 4437
rect 2717 4332 2722 4367
rect 2589 4202 2594 4207
rect 2599 4202 2600 4207
rect 2584 4007 2600 4202
rect 2589 4002 2594 4007
rect 2599 4002 2600 4007
rect 2584 3807 2600 4002
rect 2589 3802 2594 3807
rect 2599 3802 2600 3807
rect 2584 3607 2600 3802
rect 2589 3602 2594 3607
rect 2599 3602 2600 3607
rect 2584 3407 2600 3602
rect 2589 3402 2594 3407
rect 2599 3402 2600 3407
rect 2584 3207 2600 3402
rect 2589 3202 2594 3207
rect 2599 3202 2600 3207
rect 2584 3007 2600 3202
rect 2589 3002 2594 3007
rect 2599 3002 2600 3007
rect 2573 2982 2578 2997
rect 2584 2807 2600 3002
rect 2621 2862 2626 3107
rect 2589 2802 2594 2807
rect 2599 2802 2600 2807
rect 2584 2607 2600 2802
rect 2589 2602 2594 2607
rect 2599 2602 2600 2607
rect 2584 2407 2600 2602
rect 2589 2402 2594 2407
rect 2599 2402 2600 2407
rect 2584 2207 2600 2402
rect 2589 2202 2594 2207
rect 2599 2202 2600 2207
rect 2077 502 2082 507
rect 2087 502 2088 507
rect 2072 307 2088 502
rect 2077 302 2082 307
rect 2087 302 2088 307
rect 2072 107 2088 302
rect 2509 152 2514 2017
rect 2541 1752 2546 2147
rect 2584 2007 2600 2202
rect 2589 2002 2594 2007
rect 2599 2002 2600 2007
rect 2584 1807 2600 2002
rect 2589 1802 2594 1807
rect 2599 1802 2600 1807
rect 2584 1607 2600 1802
rect 2589 1602 2594 1607
rect 2599 1602 2600 1607
rect 2584 1407 2600 1602
rect 2621 1492 2626 1607
rect 2589 1402 2594 1407
rect 2599 1402 2600 1407
rect 2584 1207 2600 1402
rect 2637 1282 2642 2687
rect 2589 1202 2594 1207
rect 2599 1202 2600 1207
rect 2584 1007 2600 1202
rect 2589 1002 2594 1007
rect 2599 1002 2600 1007
rect 2584 807 2600 1002
rect 2605 1002 2610 1037
rect 2589 802 2594 807
rect 2599 802 2600 807
rect 2573 762 2578 797
rect 2584 607 2600 802
rect 2605 772 2610 797
rect 2653 782 2658 2937
rect 2669 2472 2674 3257
rect 2669 2002 2674 2327
rect 2685 1882 2690 3117
rect 2701 2492 2706 3227
rect 2733 3182 2738 4367
rect 3096 4307 3112 4502
rect 3101 4302 3106 4307
rect 3111 4302 3112 4307
rect 2941 4162 2946 4187
rect 3096 4107 3112 4302
rect 3549 4392 3554 4517
rect 3533 4252 3538 4267
rect 3101 4102 3106 4107
rect 3111 4102 3112 4107
rect 2749 3012 2754 3677
rect 2749 1922 2754 2717
rect 2765 2142 2770 2437
rect 2813 2162 2818 2257
rect 2765 1722 2770 2137
rect 2797 2062 2802 2087
rect 2701 1292 2706 1567
rect 2829 1542 2834 4037
rect 2989 3712 2994 3997
rect 3096 3907 3112 4102
rect 3101 3902 3106 3907
rect 3111 3902 3112 3907
rect 3096 3707 3112 3902
rect 3101 3702 3106 3707
rect 3111 3702 3112 3707
rect 2909 2252 2914 2397
rect 2941 2392 2946 3107
rect 3005 2452 3010 2757
rect 2797 1182 2802 1307
rect 2829 792 2834 1537
rect 2845 1112 2850 2137
rect 2941 1212 2946 2377
rect 2845 772 2850 1107
rect 2957 882 2962 2297
rect 3005 1472 3010 2447
rect 3037 2182 3042 3247
rect 3053 1282 3058 1907
rect 3069 1162 3074 3657
rect 3096 3507 3112 3702
rect 3101 3502 3106 3507
rect 3111 3502 3112 3507
rect 3096 3307 3112 3502
rect 3101 3302 3106 3307
rect 3111 3302 3112 3307
rect 3085 2642 3090 3267
rect 3096 3107 3112 3302
rect 3133 4182 3138 4197
rect 3133 3122 3138 4177
rect 3197 3132 3202 3277
rect 3101 3102 3106 3107
rect 3111 3102 3112 3107
rect 3096 2907 3112 3102
rect 3101 2902 3106 2907
rect 3111 2902 3112 2907
rect 3096 2707 3112 2902
rect 3101 2702 3106 2707
rect 3111 2702 3112 2707
rect 3096 2507 3112 2702
rect 3133 2572 3138 2617
rect 3101 2502 3106 2507
rect 3111 2502 3112 2507
rect 3096 2307 3112 2502
rect 3117 2472 3122 2497
rect 3117 2382 3122 2437
rect 3165 2352 3170 2907
rect 3101 2302 3106 2307
rect 3111 2302 3112 2307
rect 3096 2107 3112 2302
rect 3101 2102 3106 2107
rect 3111 2102 3112 2107
rect 3096 1907 3112 2102
rect 3101 1902 3106 1907
rect 3111 1902 3112 1907
rect 3085 1462 3090 1757
rect 3096 1707 3112 1902
rect 3101 1702 3106 1707
rect 3111 1702 3112 1707
rect 3096 1507 3112 1702
rect 3117 1702 3122 1767
rect 3149 1642 3154 2157
rect 3181 2032 3186 3067
rect 3101 1502 3106 1507
rect 3111 1502 3112 1507
rect 3096 1307 3112 1502
rect 3101 1302 3106 1307
rect 3111 1302 3112 1307
rect 3096 1107 3112 1302
rect 3213 1302 3218 3807
rect 3293 3372 3298 3947
rect 3229 1502 3234 2297
rect 3133 1122 3138 1137
rect 3101 1102 3106 1107
rect 3111 1102 3112 1107
rect 3096 907 3112 1102
rect 3197 1022 3202 1217
rect 3101 902 3106 907
rect 3111 902 3112 907
rect 2589 602 2594 607
rect 2599 602 2600 607
rect 2584 407 2600 602
rect 2589 402 2594 407
rect 2599 402 2600 407
rect 2584 207 2600 402
rect 2589 202 2594 207
rect 2599 202 2600 207
rect 2077 102 2082 107
rect 2087 102 2088 107
rect 2072 -30 2088 102
rect 2584 7 2600 202
rect 2589 2 2594 7
rect 2599 2 2600 7
rect 2584 -30 2600 2
rect 3096 707 3112 902
rect 3277 802 3282 1727
rect 3293 1482 3298 2307
rect 3309 2212 3314 3397
rect 3309 942 3314 1917
rect 3325 1612 3330 3067
rect 3341 2352 3346 3977
rect 3373 3222 3378 3637
rect 3373 2612 3378 3217
rect 3357 1912 3362 2437
rect 3389 1782 3394 3907
rect 3405 3622 3410 3837
rect 3405 2872 3410 2887
rect 3338 1527 3346 1532
rect 3309 762 3314 937
rect 3341 862 3346 1527
rect 3405 1252 3410 2117
rect 3421 1952 3426 3567
rect 3437 2312 3442 4187
rect 3485 3682 3490 3757
rect 3533 3732 3538 4247
rect 3469 2572 3474 3157
rect 3437 2072 3442 2227
rect 3453 1822 3458 2527
rect 3469 1862 3474 2427
rect 3485 1882 3490 2387
rect 3469 1422 3474 1767
rect 3405 1122 3410 1137
rect 3101 702 3106 707
rect 3111 702 3112 707
rect 3096 507 3112 702
rect 3469 662 3474 1207
rect 3101 502 3106 507
rect 3111 502 3112 507
rect 3096 307 3112 502
rect 3101 302 3106 307
rect 3111 302 3112 307
rect 3096 107 3112 302
rect 3485 162 3490 1217
rect 3501 552 3506 1947
rect 3517 1912 3522 3607
rect 3533 2012 3538 3727
rect 3549 2952 3554 4387
rect 3608 4407 3624 4602
rect 3613 4402 3618 4407
rect 3623 4402 3624 4407
rect 3608 4207 3624 4402
rect 4112 4907 4128 4930
rect 4117 4902 4122 4907
rect 4127 4902 4128 4907
rect 4112 4707 4128 4902
rect 4117 4702 4122 4707
rect 4127 4702 4128 4707
rect 4112 4507 4128 4702
rect 4117 4502 4122 4507
rect 4127 4502 4128 4507
rect 3613 4202 3618 4207
rect 3623 4202 3624 4207
rect 3608 4007 3624 4202
rect 3613 4002 3618 4007
rect 3623 4002 3624 4007
rect 3597 3432 3602 3817
rect 3565 2412 3570 2427
rect 3549 1542 3554 2007
rect 3565 1372 3570 2347
rect 3581 2312 3586 3137
rect 3597 2372 3602 3427
rect 3608 3807 3624 4002
rect 3613 3802 3618 3807
rect 3623 3802 3624 3807
rect 3608 3607 3624 3802
rect 3613 3602 3618 3607
rect 3623 3602 3624 3607
rect 3608 3407 3624 3602
rect 3613 3402 3618 3407
rect 3623 3402 3624 3407
rect 3608 3207 3624 3402
rect 3613 3202 3618 3207
rect 3623 3202 3624 3207
rect 3608 3007 3624 3202
rect 3613 3002 3618 3007
rect 3623 3002 3624 3007
rect 3608 2807 3624 3002
rect 3629 2952 3634 3467
rect 3645 2982 3650 3557
rect 3613 2802 3618 2807
rect 3623 2802 3624 2807
rect 3608 2607 3624 2802
rect 3629 2722 3634 2797
rect 3613 2602 3618 2607
rect 3623 2602 3624 2607
rect 3608 2407 3624 2602
rect 3613 2402 3618 2407
rect 3623 2402 3624 2407
rect 3608 2207 3624 2402
rect 3613 2202 3618 2207
rect 3623 2202 3624 2207
rect 3565 772 3570 927
rect 3581 842 3586 2007
rect 3608 2007 3624 2202
rect 3629 2082 3634 2447
rect 3613 2002 3618 2007
rect 3623 2002 3624 2007
rect 3597 1362 3602 1907
rect 3608 1807 3624 2002
rect 3613 1802 3618 1807
rect 3623 1802 3624 1807
rect 3608 1607 3624 1802
rect 3613 1602 3618 1607
rect 3623 1602 3624 1607
rect 3608 1407 3624 1602
rect 3613 1402 3618 1407
rect 3623 1402 3624 1407
rect 3608 1207 3624 1402
rect 3613 1202 3618 1207
rect 3623 1202 3624 1207
rect 3608 1007 3624 1202
rect 3661 1102 3666 2837
rect 3677 1452 3682 3557
rect 3693 1672 3698 2737
rect 3709 1182 3714 2037
rect 3725 2012 3730 3717
rect 3613 1002 3618 1007
rect 3623 1002 3624 1007
rect 3608 807 3624 1002
rect 3613 802 3618 807
rect 3623 802 3624 807
rect 3608 607 3624 802
rect 3741 752 3746 3247
rect 3757 1882 3762 3627
rect 3773 2372 3778 2887
rect 3757 742 3762 1607
rect 3773 1512 3778 2237
rect 3805 2142 3810 2237
rect 3789 1572 3794 1777
rect 3805 1482 3810 1497
rect 3821 1442 3826 3497
rect 3917 3072 3922 3507
rect 3933 2992 3938 4307
rect 4112 4307 4128 4502
rect 4632 4807 4648 4930
rect 4637 4802 4642 4807
rect 4647 4802 4648 4807
rect 4632 4607 4648 4802
rect 4637 4602 4642 4607
rect 4647 4602 4648 4607
rect 4117 4302 4122 4307
rect 4127 4302 4128 4307
rect 3837 2592 3842 2877
rect 3869 1952 3874 2977
rect 3933 2782 3938 2867
rect 3613 602 3618 607
rect 3623 602 3624 607
rect 3608 407 3624 602
rect 3613 402 3618 407
rect 3623 402 3624 407
rect 3608 207 3624 402
rect 3805 262 3810 1357
rect 3853 1062 3858 1567
rect 3869 1362 3874 1947
rect 3885 952 3890 2747
rect 3901 1502 3906 2757
rect 3933 2042 3938 2447
rect 3933 1842 3938 1887
rect 3949 1392 3954 3657
rect 3981 3282 3986 4137
rect 4013 3162 4018 4247
rect 3965 912 3970 2897
rect 3981 2182 3986 2647
rect 3997 1682 4002 2887
rect 4029 732 4034 3297
rect 4045 3002 4050 4217
rect 4112 4107 4128 4302
rect 4117 4102 4122 4107
rect 4127 4102 4128 4107
rect 4061 1912 4066 4047
rect 4093 4047 4101 4052
rect 4077 2502 4082 3637
rect 4093 3022 4098 4047
rect 4112 3907 4128 4102
rect 4117 3902 4122 3907
rect 4127 3902 4128 3907
rect 4112 3707 4128 3902
rect 4117 3702 4122 3707
rect 4127 3702 4128 3707
rect 4112 3507 4128 3702
rect 4117 3502 4122 3507
rect 4127 3502 4128 3507
rect 4112 3307 4128 3502
rect 4117 3302 4122 3307
rect 4127 3302 4128 3307
rect 4112 3107 4128 3302
rect 4117 3102 4122 3107
rect 4127 3102 4128 3107
rect 4077 1372 4082 2487
rect 4093 2132 4098 2917
rect 4112 2907 4128 3102
rect 4117 2902 4122 2907
rect 4127 2902 4128 2907
rect 4112 2707 4128 2902
rect 4117 2702 4122 2707
rect 4127 2702 4128 2707
rect 4112 2507 4128 2702
rect 4117 2502 4122 2507
rect 4127 2502 4128 2507
rect 4112 2307 4128 2502
rect 4117 2302 4122 2307
rect 4127 2302 4128 2307
rect 4112 2107 4128 2302
rect 4117 2102 4122 2107
rect 4127 2102 4128 2107
rect 4093 1162 4098 2077
rect 4112 1907 4128 2102
rect 4117 1902 4122 1907
rect 4127 1902 4128 1907
rect 4112 1707 4128 1902
rect 4117 1702 4122 1707
rect 4127 1702 4128 1707
rect 4112 1507 4128 1702
rect 4117 1502 4122 1507
rect 4127 1502 4128 1507
rect 4112 1307 4128 1502
rect 4141 1372 4146 2767
rect 4157 2062 4162 3027
rect 4173 1942 4178 2927
rect 4189 2052 4194 3007
rect 4205 2482 4210 3307
rect 4221 1982 4226 3857
rect 4269 3592 4274 4257
rect 4397 4232 4402 4407
rect 4632 4407 4648 4602
rect 4637 4402 4642 4407
rect 4647 4402 4648 4407
rect 4269 3512 4274 3587
rect 4253 2262 4258 2987
rect 4285 2252 4290 3837
rect 4117 1302 4122 1307
rect 4127 1302 4128 1307
rect 4029 452 4034 727
rect 4112 1107 4128 1302
rect 4117 1102 4122 1107
rect 4127 1102 4128 1107
rect 4112 907 4128 1102
rect 4117 902 4122 907
rect 4127 902 4128 907
rect 4112 707 4128 902
rect 4237 842 4242 2237
rect 4301 1892 4306 2887
rect 4301 752 4306 1867
rect 4333 1752 4338 3647
rect 4397 3472 4402 4227
rect 4365 3467 4373 3472
rect 4365 2442 4370 3467
rect 4349 1902 4354 2357
rect 4333 952 4338 1747
rect 4381 1222 4386 2807
rect 4397 1662 4402 2687
rect 4413 752 4418 2287
rect 4429 1752 4434 2397
rect 4445 1682 4450 2587
rect 4461 1702 4466 2967
rect 4477 2082 4482 3337
rect 4509 2082 4514 3807
rect 4525 3182 4530 4137
rect 4541 3342 4546 4397
rect 4557 3392 4562 4337
rect 4632 4207 4648 4402
rect 4637 4202 4642 4207
rect 4647 4202 4648 4207
rect 4525 3152 4530 3177
rect 4525 2762 4530 2787
rect 4117 702 4122 707
rect 4127 702 4128 707
rect 4112 507 4128 702
rect 4477 532 4482 1857
rect 4525 1172 4530 2147
rect 4117 502 4122 507
rect 4127 502 4128 507
rect 4112 307 4128 502
rect 4117 302 4122 307
rect 4127 302 4128 307
rect 3613 202 3618 207
rect 3623 202 3624 207
rect 3101 102 3106 107
rect 3111 102 3112 107
rect 3096 -30 3112 102
rect 3608 7 3624 202
rect 3613 2 3618 7
rect 3623 2 3624 7
rect 3608 -30 3624 2
rect 4112 107 4128 302
rect 4117 102 4122 107
rect 4127 102 4128 107
rect 4112 -30 4128 102
rect 4541 62 4546 2267
rect 4557 2122 4562 3387
rect 4573 3612 4578 3927
rect 4573 2392 4578 3607
rect 4557 772 4562 1847
rect 4573 1282 4578 2247
rect 4589 2142 4594 3657
rect 4621 2882 4626 4177
rect 4632 4007 4648 4202
rect 4637 4002 4642 4007
rect 4647 4002 4648 4007
rect 4632 3807 4648 4002
rect 4637 3802 4642 3807
rect 4647 3802 4648 3807
rect 4632 3607 4648 3802
rect 4637 3602 4642 3607
rect 4647 3602 4648 3607
rect 4632 3407 4648 3602
rect 4637 3402 4642 3407
rect 4647 3402 4648 3407
rect 4632 3207 4648 3402
rect 4637 3202 4642 3207
rect 4647 3202 4648 3207
rect 4632 3007 4648 3202
rect 4637 3002 4642 3007
rect 4647 3002 4648 3007
rect 4632 2807 4648 3002
rect 4637 2802 4642 2807
rect 4647 2802 4648 2807
rect 4632 2607 4648 2802
rect 4637 2602 4642 2607
rect 4647 2602 4648 2607
rect 4632 2407 4648 2602
rect 4637 2402 4642 2407
rect 4647 2402 4648 2407
rect 4589 52 4594 2077
rect 4605 112 4610 2377
rect 4632 2207 4648 2402
rect 4637 2202 4642 2207
rect 4647 2202 4648 2207
rect 4632 2007 4648 2202
rect 4637 2002 4642 2007
rect 4647 2002 4648 2007
rect 4632 1807 4648 2002
rect 4637 1802 4642 1807
rect 4647 1802 4648 1807
rect 4621 1022 4626 1707
rect 4621 632 4626 1017
rect 4632 1607 4648 1802
rect 4637 1602 4642 1607
rect 4647 1602 4648 1607
rect 4632 1407 4648 1602
rect 4637 1402 4642 1407
rect 4647 1402 4648 1407
rect 4632 1207 4648 1402
rect 4637 1202 4642 1207
rect 4647 1202 4648 1207
rect 4632 1007 4648 1202
rect 4637 1002 4642 1007
rect 4647 1002 4648 1007
rect 4632 807 4648 1002
rect 4637 802 4642 807
rect 4647 802 4648 807
rect 4632 607 4648 802
rect 4637 602 4642 607
rect 4647 602 4648 607
rect 4632 407 4648 602
rect 4637 402 4642 407
rect 4647 402 4648 407
rect 4632 207 4648 402
rect 4637 202 4642 207
rect 4647 202 4648 207
rect 4632 7 4648 202
rect 4669 142 4674 2067
rect 4685 1182 4690 3467
rect 4717 62 4722 2087
rect 4733 1482 4738 3137
rect 4749 2162 4754 4457
rect 4749 662 4754 1827
rect 4765 1632 4770 3937
rect 4813 52 4818 1767
rect 4829 1052 4834 2267
rect 4861 1992 4866 4847
rect 4925 1922 4930 4847
rect 4861 272 4866 1697
rect 4957 82 4962 2307
rect 4973 892 4978 4017
rect 5005 92 5010 2537
rect 5021 1872 5026 2907
rect 5069 2892 5074 4367
rect 5085 2262 5090 2787
rect 5101 2632 5106 4857
rect 5021 1252 5026 1707
rect 5085 1502 5090 2077
rect 5101 192 5106 2567
rect 5117 292 5122 2947
rect 5133 2282 5138 2557
rect 5149 2432 5154 3997
rect 5149 932 5154 2417
rect 5165 2042 5170 3047
rect 5181 852 5186 2657
rect 4637 2 4642 7
rect 4647 2 4648 7
rect 4632 -30 4648 2
use CLKBUF1  CLKBUF1_99
timestamp 1607319584
transform -1 0 76 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_45
timestamp 1607319584
transform 1 0 76 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_682
timestamp 1607319584
transform 1 0 4 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_677
timestamp 1607319584
transform 1 0 100 0 1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_16
timestamp 1607319584
transform 1 0 148 0 -1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_468
timestamp 1607319584
transform -1 0 228 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_826
timestamp 1607319584
transform 1 0 220 0 -1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_109
timestamp 1607319584
transform 1 0 228 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_137
timestamp 1607319584
transform -1 0 284 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_458
timestamp 1607319584
transform -1 0 316 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_341
timestamp 1607319584
transform 1 0 316 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_295
timestamp 1607319584
transform 1 0 316 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_338
timestamp 1607319584
transform 1 0 332 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_1683
timestamp 1607319584
transform 1 0 412 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_339
timestamp 1607319584
transform 1 0 444 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_1677
timestamp 1607319584
transform 1 0 428 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1676
timestamp 1607319584
transform -1 0 492 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1682
timestamp 1607319584
transform -1 0 524 0 1 105
box -2 -3 34 103
use FILL  FILL_0_0_0
timestamp 1607319584
transform 1 0 540 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1607319584
transform 1 0 548 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_685
timestamp 1607319584
transform 1 0 556 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_0_0
timestamp 1607319584
transform 1 0 524 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1607319584
transform 1 0 532 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_1679
timestamp 1607319584
transform 1 0 540 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_474
timestamp 1607319584
transform 1 0 572 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_694
timestamp 1607319584
transform 1 0 604 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_342
timestamp 1607319584
transform -1 0 748 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_473
timestamp 1607319584
transform -1 0 732 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1685
timestamp 1607319584
transform 1 0 748 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1684
timestamp 1607319584
transform -1 0 812 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_471
timestamp 1607319584
transform 1 0 732 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_472
timestamp 1607319584
transform -1 0 796 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_470
timestamp 1607319584
transform 1 0 796 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_344
timestamp 1607319584
transform 1 0 812 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_1689
timestamp 1607319584
transform 1 0 908 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_469
timestamp 1607319584
transform 1 0 828 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_683
timestamp 1607319584
transform 1 0 860 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_1688
timestamp 1607319584
transform 1 0 940 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_365
timestamp 1607319584
transform 1 0 972 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_355
timestamp 1607319584
transform 1 0 956 0 1 105
box -2 -3 98 103
use FILL  FILL_0_1_0
timestamp 1607319584
transform -1 0 1076 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1607319584
transform -1 0 1084 0 -1 105
box -2 -3 10 103
use BUFX4  BUFX4_315
timestamp 1607319584
transform -1 0 1116 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1607319584
transform 1 0 1052 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1607319584
transform 1 0 1060 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_6
timestamp 1607319584
transform 1 0 1068 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_363
timestamp 1607319584
transform 1 0 1100 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_357
timestamp 1607319584
transform 1 0 1116 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_590
timestamp 1607319584
transform 1 0 1212 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_21
timestamp 1607319584
transform 1 0 1196 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_54
timestamp 1607319584
transform 1 0 1308 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_22
timestamp 1607319584
transform -1 0 1260 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1607319584
transform 1 0 1260 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_25
timestamp 1607319584
transform -1 0 1324 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1607319584
transform -1 0 1364 0 -1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_34
timestamp 1607319584
transform 1 0 1364 0 -1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_10
timestamp 1607319584
transform 1 0 1324 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_9
timestamp 1607319584
transform -1 0 1388 0 1 105
box -2 -3 34 103
use INVX1  INVX1_466
timestamp 1607319584
transform 1 0 1388 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_23
timestamp 1607319584
transform 1 0 1404 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_619
timestamp 1607319584
transform 1 0 1436 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_24
timestamp 1607319584
transform -1 0 1468 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_364
timestamp 1607319584
transform 1 0 1468 0 1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_52
timestamp 1607319584
transform 1 0 1532 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_2_0
timestamp 1607319584
transform -1 0 1572 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1607319584
transform -1 0 1580 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_66
timestamp 1607319584
transform -1 0 1604 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_588
timestamp 1607319584
transform 1 0 1604 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_2_0
timestamp 1607319584
transform 1 0 1564 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1607319584
transform 1 0 1572 0 1 105
box -2 -3 10 103
use BUFX4  BUFX4_318
timestamp 1607319584
transform 1 0 1580 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_372
timestamp 1607319584
transform 1 0 1612 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_368
timestamp 1607319584
transform -1 0 1796 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_40
timestamp 1607319584
transform 1 0 1708 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_365
timestamp 1607319584
transform -1 0 1828 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_39
timestamp 1607319584
transform 1 0 1740 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_366
timestamp 1607319584
transform -1 0 1804 0 1 105
box -2 -3 34 103
use INVX1  INVX1_212
timestamp 1607319584
transform 1 0 1804 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_1000
timestamp 1607319584
transform 1 0 1820 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_8
timestamp 1607319584
transform -1 0 1900 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_362
timestamp 1607319584
transform 1 0 1900 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_350
timestamp 1607319584
transform 1 0 1852 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_349
timestamp 1607319584
transform -1 0 1916 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_611
timestamp 1607319584
transform -1 0 2012 0 1 105
box -2 -3 98 103
use BUFX4  BUFX4_317
timestamp 1607319584
transform 1 0 1996 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_376
timestamp 1607319584
transform 1 0 2012 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_20
timestamp 1607319584
transform -1 0 2060 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_3
timestamp 1607319584
transform 1 0 2060 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_3_0
timestamp 1607319584
transform 1 0 2084 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1607319584
transform 1 0 2092 0 -1 105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_52
timestamp 1607319584
transform 1 0 2100 0 -1 105
box -2 -3 74 103
use FILL  FILL_1_3_0
timestamp 1607319584
transform 1 0 2108 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1607319584
transform 1 0 2116 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_48
timestamp 1607319584
transform 1 0 2124 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_64
timestamp 1607319584
transform 1 0 2172 0 -1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_47
timestamp 1607319584
transform -1 0 2188 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_32
timestamp 1607319584
transform -1 0 2220 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_31
timestamp 1607319584
transform -1 0 2252 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_252
timestamp 1607319584
transform 1 0 2244 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_19
timestamp 1607319584
transform -1 0 2284 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1607319584
transform 1 0 2284 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_29
timestamp 1607319584
transform 1 0 2316 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_246
timestamp 1607319584
transform 1 0 2340 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_367
timestamp 1607319584
transform 1 0 2348 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_254
timestamp 1607319584
transform 1 0 2436 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1027
timestamp 1607319584
transform -1 0 2540 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_250
timestamp 1607319584
transform -1 0 2628 0 -1 105
box -2 -3 98 103
use FILL  FILL_0_4_0
timestamp 1607319584
transform -1 0 2636 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_4_0
timestamp 1607319584
transform 1 0 2540 0 1 105
box -2 -3 10 103
use FILL  FILL_1_4_1
timestamp 1607319584
transform 1 0 2548 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_244
timestamp 1607319584
transform 1 0 2556 0 1 105
box -2 -3 98 103
use FILL  FILL_0_4_1
timestamp 1607319584
transform -1 0 2644 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_1581
timestamp 1607319584
transform -1 0 2676 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1573
timestamp 1607319584
transform 1 0 2676 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_89
timestamp 1607319584
transform -1 0 2740 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1561
timestamp 1607319584
transform -1 0 2684 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1560
timestamp 1607319584
transform -1 0 2716 0 1 105
box -2 -3 34 103
use INVX1  INVX1_204
timestamp 1607319584
transform 1 0 2716 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_276
timestamp 1607319584
transform 1 0 2740 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_347
timestamp 1607319584
transform -1 0 2796 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_222
timestamp 1607319584
transform 1 0 2796 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_1565
timestamp 1607319584
transform 1 0 2732 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1564
timestamp 1607319584
transform -1 0 2796 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1576
timestamp 1607319584
transform -1 0 2828 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1577
timestamp 1607319584
transform -1 0 2860 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_208
timestamp 1607319584
transform 1 0 2892 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_1580
timestamp 1607319584
transform -1 0 2892 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1572
timestamp 1607319584
transform 1 0 2892 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_230
timestamp 1607319584
transform -1 0 3020 0 1 105
box -2 -3 98 103
use BUFX4  BUFX4_94
timestamp 1607319584
transform -1 0 3020 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1519
timestamp 1607319584
transform -1 0 3052 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_35
timestamp 1607319584
transform 1 0 3020 0 1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_1520
timestamp 1607319584
transform -1 0 3084 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_5_0
timestamp 1607319584
transform -1 0 3092 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_5_1
timestamp 1607319584
transform -1 0 3100 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_224
timestamp 1607319584
transform -1 0 3196 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_5_0
timestamp 1607319584
transform -1 0 3100 0 1 105
box -2 -3 10 103
use FILL  FILL_1_5_1
timestamp 1607319584
transform -1 0 3108 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_225
timestamp 1607319584
transform -1 0 3204 0 1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_278
timestamp 1607319584
transform 1 0 3196 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_349
timestamp 1607319584
transform 1 0 3228 0 -1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_340
timestamp 1607319584
transform 1 0 3204 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_196
timestamp 1607319584
transform -1 0 3348 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_216
timestamp 1607319584
transform 1 0 3252 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_195
timestamp 1607319584
transform 1 0 3348 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_458
timestamp 1607319584
transform 1 0 3348 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_1246
timestamp 1607319584
transform 1 0 3364 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_699
timestamp 1607319584
transform -1 0 3420 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_1495
timestamp 1607319584
transform -1 0 3452 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1496
timestamp 1607319584
transform -1 0 3476 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1494
timestamp 1607319584
transform -1 0 3508 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1493
timestamp 1607319584
transform -1 0 3540 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_698
timestamp 1607319584
transform -1 0 3476 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_1245
timestamp 1607319584
transform -1 0 3508 0 1 105
box -2 -3 34 103
use INVX1  INVX1_457
timestamp 1607319584
transform -1 0 3524 0 1 105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_36
timestamp 1607319584
transform -1 0 3596 0 1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_900
timestamp 1607319584
transform 1 0 3540 0 -1 105
box -2 -3 98 103
use FILL  FILL_0_6_0
timestamp 1607319584
transform 1 0 3636 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_6_0
timestamp 1607319584
transform 1 0 3596 0 1 105
box -2 -3 10 103
use FILL  FILL_1_6_1
timestamp 1607319584
transform 1 0 3604 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_1503
timestamp 1607319584
transform 1 0 3612 0 1 105
box -2 -3 34 103
use FILL  FILL_0_6_1
timestamp 1607319584
transform 1 0 3644 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_682
timestamp 1607319584
transform 1 0 3652 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_681
timestamp 1607319584
transform -1 0 3716 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_51
timestamp 1607319584
transform -1 0 3788 0 -1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_1504
timestamp 1607319584
transform -1 0 3676 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_200
timestamp 1607319584
transform -1 0 3772 0 1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_9
timestamp 1607319584
transform 1 0 3788 0 -1 105
box -2 -3 74 103
use INVX1  INVX1_137
timestamp 1607319584
transform 1 0 3772 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_1510
timestamp 1607319584
transform 1 0 3788 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_1509
timestamp 1607319584
transform 1 0 3820 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_912
timestamp 1607319584
transform 1 0 3860 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_203
timestamp 1607319584
transform -1 0 3948 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_706
timestamp 1607319584
transform -1 0 3988 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_705
timestamp 1607319584
transform -1 0 4020 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_692
timestamp 1607319584
transform 1 0 4020 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_245
timestamp 1607319584
transform 1 0 3948 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_910
timestamp 1607319584
transform 1 0 3964 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_691
timestamp 1607319584
transform 1 0 4052 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_7_0
timestamp 1607319584
transform 1 0 4084 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_7_1
timestamp 1607319584
transform 1 0 4092 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_905
timestamp 1607319584
transform 1 0 4100 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_702
timestamp 1607319584
transform 1 0 4060 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_701
timestamp 1607319584
transform -1 0 4124 0 1 105
box -2 -3 34 103
use FILL  FILL_1_7_0
timestamp 1607319584
transform 1 0 4124 0 1 105
box -2 -3 10 103
use FILL  FILL_1_7_1
timestamp 1607319584
transform 1 0 4132 0 1 105
box -2 -3 10 103
use BUFX4  BUFX4_67
timestamp 1607319584
transform 1 0 4140 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_690
timestamp 1607319584
transform 1 0 4196 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_689
timestamp 1607319584
transform 1 0 4228 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_538
timestamp 1607319584
transform 1 0 4172 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_1097
timestamp 1607319584
transform -1 0 4228 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_699
timestamp 1607319584
transform 1 0 4228 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_904
timestamp 1607319584
transform -1 0 4356 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_909
timestamp 1607319584
transform -1 0 4356 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_675
timestamp 1607319584
transform 1 0 4356 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_676
timestamp 1607319584
transform -1 0 4420 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_897
timestamp 1607319584
transform 1 0 4420 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_700
timestamp 1607319584
transform -1 0 4388 0 1 105
box -2 -3 34 103
use INVX1  INVX1_501
timestamp 1607319584
transform 1 0 4388 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_907
timestamp 1607319584
transform -1 0 4500 0 1 105
box -2 -3 98 103
use BUFX4  BUFX4_137
timestamp 1607319584
transform -1 0 4548 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_218
timestamp 1607319584
transform -1 0 4580 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_66
timestamp 1607319584
transform 1 0 4500 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_21
timestamp 1607319584
transform -1 0 4604 0 1 105
box -2 -3 74 103
use NOR2X1  NOR2X1_286
timestamp 1607319584
transform -1 0 4604 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_8_0
timestamp 1607319584
transform -1 0 4612 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_8_1
timestamp 1607319584
transform -1 0 4620 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_169
timestamp 1607319584
transform -1 0 4716 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_309
timestamp 1607319584
transform -1 0 4620 0 1 105
box -2 -3 18 103
use FILL  FILL_1_8_0
timestamp 1607319584
transform -1 0 4628 0 1 105
box -2 -3 10 103
use FILL  FILL_1_8_1
timestamp 1607319584
transform -1 0 4636 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_901
timestamp 1607319584
transform -1 0 4732 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1607319584
transform 1 0 4716 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_684
timestamp 1607319584
transform 1 0 4732 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_880
timestamp 1607319584
transform -1 0 4844 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_98
timestamp 1607319584
transform -1 0 4916 0 -1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_683
timestamp 1607319584
transform -1 0 4796 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_15
timestamp 1607319584
transform -1 0 4844 0 1 105
box -2 -3 50 103
use OAI21X1  OAI21X1_679
timestamp 1607319584
transform 1 0 4844 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_154
timestamp 1607319584
transform 1 0 4916 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_680
timestamp 1607319584
transform -1 0 4908 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_903
timestamp 1607319584
transform -1 0 5004 0 1 105
box -2 -3 98 103
use BUFX4  BUFX4_447
timestamp 1607319584
transform -1 0 5044 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_37
timestamp 1607319584
transform -1 0 5116 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_899
timestamp 1607319584
transform -1 0 5100 0 1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_24
timestamp 1607319584
transform 1 0 5116 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_151
timestamp 1607319584
transform -1 0 5196 0 1 105
box -2 -3 98 103
use FILL  FILL_1_1
timestamp 1607319584
transform -1 0 5196 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_678
timestamp 1607319584
transform 1 0 4 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_460
timestamp 1607319584
transform 1 0 100 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_459
timestamp 1607319584
transform -1 0 164 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_467
timestamp 1607319584
transform -1 0 196 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_681
timestamp 1607319584
transform 1 0 196 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_457
timestamp 1607319584
transform -1 0 324 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_697
timestamp 1607319584
transform 1 0 324 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_497
timestamp 1607319584
transform -1 0 452 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_359
timestamp 1607319584
transform 1 0 452 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_686
timestamp 1607319584
transform 1 0 468 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_0_0
timestamp 1607319584
transform 1 0 564 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1607319584
transform 1 0 572 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_475
timestamp 1607319584
transform 1 0 580 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_476
timestamp 1607319584
transform -1 0 644 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_592
timestamp 1607319584
transform -1 0 668 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_1678
timestamp 1607319584
transform -1 0 700 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_523
timestamp 1607319584
transform -1 0 724 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_492
timestamp 1607319584
transform 1 0 724 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_491
timestamp 1607319584
transform -1 0 788 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_684
timestamp 1607319584
transform 1 0 788 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_702
timestamp 1607319584
transform 1 0 884 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1701
timestamp 1607319584
transform 1 0 980 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1700
timestamp 1607319584
transform -1 0 1044 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1607319584
transform -1 0 1052 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1607319584
transform -1 0 1060 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_266
timestamp 1607319584
transform -1 0 1084 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_5
timestamp 1607319584
transform -1 0 1116 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_352
timestamp 1607319584
transform 1 0 1116 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1705
timestamp 1607319584
transform 1 0 1212 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_364
timestamp 1607319584
transform -1 0 1268 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_1704
timestamp 1607319584
transform 1 0 1268 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_319
timestamp 1607319584
transform -1 0 1332 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_275
timestamp 1607319584
transform 1 0 1332 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_53
timestamp 1607319584
transform 1 0 1348 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_379
timestamp 1607319584
transform -1 0 1476 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_54
timestamp 1607319584
transform -1 0 1508 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_586
timestamp 1607319584
transform -1 0 1532 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_433
timestamp 1607319584
transform 1 0 1532 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_2_0
timestamp 1607319584
transform 1 0 1556 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1607319584
transform 1 0 1564 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_44
timestamp 1607319584
transform 1 0 1572 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1607319584
transform 1 0 1604 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_374
timestamp 1607319584
transform 1 0 1636 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_211
timestamp 1607319584
transform -1 0 1748 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_7
timestamp 1607319584
transform 1 0 1748 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_8
timestamp 1607319584
transform -1 0 1812 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_356
timestamp 1607319584
transform -1 0 1908 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_381
timestamp 1607319584
transform -1 0 1932 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_434
timestamp 1607319584
transform 1 0 1932 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_56
timestamp 1607319584
transform 1 0 1956 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_55
timestamp 1607319584
transform -1 0 2020 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_380
timestamp 1607319584
transform -1 0 2116 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_3_0
timestamp 1607319584
transform 1 0 2116 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1607319584
transform 1 0 2124 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_360
timestamp 1607319584
transform 1 0 2132 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_16
timestamp 1607319584
transform 1 0 2228 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1607319584
transform -1 0 2292 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_378
timestamp 1607319584
transform 1 0 2292 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_35
timestamp 1607319584
transform 1 0 2388 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1607319584
transform -1 0 2452 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_370
timestamp 1607319584
transform -1 0 2548 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_4_0
timestamp 1607319584
transform 1 0 2548 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_4_1
timestamp 1607319584
transform 1 0 2556 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_232
timestamp 1607319584
transform 1 0 2564 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1551
timestamp 1607319584
transform -1 0 2692 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1552
timestamp 1607319584
transform -1 0 2724 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_992
timestamp 1607319584
transform 1 0 2724 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_425
timestamp 1607319584
transform -1 0 2780 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_228
timestamp 1607319584
transform 1 0 2780 0 -1 305
box -2 -3 98 103
use BUFX4  BUFX4_95
timestamp 1607319584
transform 1 0 2876 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1547
timestamp 1607319584
transform 1 0 2908 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1548
timestamp 1607319584
transform -1 0 2972 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1550
timestamp 1607319584
transform 1 0 2972 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1549
timestamp 1607319584
transform 1 0 3004 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_231
timestamp 1607319584
transform 1 0 3036 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_5_0
timestamp 1607319584
transform 1 0 3132 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_5_1
timestamp 1607319584
transform 1 0 3140 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_1537
timestamp 1607319584
transform 1 0 3148 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1538
timestamp 1607319584
transform -1 0 3212 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_223
timestamp 1607319584
transform 1 0 3212 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_277
timestamp 1607319584
transform 1 0 3308 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_348
timestamp 1607319584
transform -1 0 3364 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_1536
timestamp 1607319584
transform 1 0 3364 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1535
timestamp 1607319584
transform -1 0 3428 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_630
timestamp 1607319584
transform -1 0 3452 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_194
timestamp 1607319584
transform -1 0 3548 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1499
timestamp 1607319584
transform 1 0 3548 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_6_0
timestamp 1607319584
transform -1 0 3588 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_6_1
timestamp 1607319584
transform -1 0 3596 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_198
timestamp 1607319584
transform -1 0 3692 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1500
timestamp 1607319584
transform -1 0 3724 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1501
timestamp 1607319584
transform 1 0 3724 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1502
timestamp 1607319584
transform 1 0 3756 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_199
timestamp 1607319584
transform -1 0 3884 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_271
timestamp 1607319584
transform 1 0 3884 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_217
timestamp 1607319584
transform -1 0 4012 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_149
timestamp 1607319584
transform 1 0 4012 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_185
timestamp 1607319584
transform -1 0 4068 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_926
timestamp 1607319584
transform -1 0 4164 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_7_0
timestamp 1607319584
transform -1 0 4172 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_7_1
timestamp 1607319584
transform -1 0 4180 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_745
timestamp 1607319584
transform -1 0 4204 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_697
timestamp 1607319584
transform 1 0 4204 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_698
timestamp 1607319584
transform -1 0 4268 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_928
timestamp 1607319584
transform 1 0 4268 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1289
timestamp 1607319584
transform -1 0 4396 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_695
timestamp 1607319584
transform 1 0 4396 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_696
timestamp 1607319584
transform -1 0 4460 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_925
timestamp 1607319584
transform -1 0 4556 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_941
timestamp 1607319584
transform 1 0 4556 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_8_0
timestamp 1607319584
transform 1 0 4652 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_8_1
timestamp 1607319584
transform 1 0 4660 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_157
timestamp 1607319584
transform 1 0 4668 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_195
timestamp 1607319584
transform 1 0 4700 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_687
timestamp 1607319584
transform 1 0 4724 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_688
timestamp 1607319584
transform -1 0 4788 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_191
timestamp 1607319584
transform -1 0 4812 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_937
timestamp 1607319584
transform -1 0 4908 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_921
timestamp 1607319584
transform -1 0 5004 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_939
timestamp 1607319584
transform 1 0 5004 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1029
timestamp 1607319584
transform 1 0 5100 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_662
timestamp 1607319584
transform 1 0 4 0 1 305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_38
timestamp 1607319584
transform 1 0 100 0 1 305
box -2 -3 74 103
use OAI21X1  OAI21X1_465
timestamp 1607319584
transform 1 0 172 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_466
timestamp 1607319584
transform -1 0 236 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_679
timestamp 1607319584
transform 1 0 236 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_462
timestamp 1607319584
transform 1 0 332 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_461
timestamp 1607319584
transform 1 0 364 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_498
timestamp 1607319584
transform -1 0 428 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_482
timestamp 1607319584
transform 1 0 428 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_481
timestamp 1607319584
transform 1 0 460 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1607319584
transform 1 0 492 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1607319584
transform 1 0 500 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_689
timestamp 1607319584
transform 1 0 508 0 1 305
box -2 -3 98 103
use INVX1  INVX1_423
timestamp 1607319584
transform 1 0 604 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_1147
timestamp 1607319584
transform 1 0 620 0 1 305
box -2 -3 34 103
use INVX1  INVX1_146
timestamp 1607319584
transform 1 0 652 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_1083
timestamp 1607319584
transform 1 0 668 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_687
timestamp 1607319584
transform 1 0 700 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_478
timestamp 1607319584
transform 1 0 796 0 1 305
box -2 -3 34 103
use INVX1  INVX1_360
timestamp 1607319584
transform 1 0 828 0 1 305
box -2 -3 18 103
use INVX1  INVX1_82
timestamp 1607319584
transform 1 0 844 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_507
timestamp 1607319584
transform 1 0 860 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_508
timestamp 1607319584
transform -1 0 924 0 1 305
box -2 -3 34 103
use INVX1  INVX1_338
timestamp 1607319584
transform 1 0 924 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_350
timestamp 1607319584
transform 1 0 940 0 1 305
box -2 -3 98 103
use INVX1  INVX1_147
timestamp 1607319584
transform 1 0 1036 0 1 305
box -2 -3 18 103
use FILL  FILL_3_1_0
timestamp 1607319584
transform 1 0 1052 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1607319584
transform 1 0 1060 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_1693
timestamp 1607319584
transform 1 0 1068 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1692
timestamp 1607319584
transform 1 0 1100 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_616
timestamp 1607319584
transform 1 0 1132 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_360
timestamp 1607319584
transform -1 0 1260 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_101
timestamp 1607319584
transform -1 0 1292 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_371
timestamp 1607319584
transform 1 0 1292 0 1 305
box -2 -3 98 103
use INVX1  INVX1_148
timestamp 1607319584
transform 1 0 1388 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_37
timestamp 1607319584
transform -1 0 1436 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_38
timestamp 1607319584
transform -1 0 1468 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_314
timestamp 1607319584
transform 1 0 1468 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_42
timestamp 1607319584
transform 1 0 1500 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_41
timestamp 1607319584
transform 1 0 1532 0 1 305
box -2 -3 34 103
use FILL  FILL_3_2_0
timestamp 1607319584
transform 1 0 1564 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1607319584
transform 1 0 1572 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_373
timestamp 1607319584
transform 1 0 1580 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_999
timestamp 1607319584
transform -1 0 1708 0 1 305
box -2 -3 34 103
use INVX1  INVX1_340
timestamp 1607319584
transform 1 0 1708 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_12
timestamp 1607319584
transform 1 0 1724 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1607319584
transform 1 0 1756 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_358
timestamp 1607319584
transform -1 0 1884 0 1 305
box -2 -3 98 103
use INVX1  INVX1_163
timestamp 1607319584
transform 1 0 1884 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_951
timestamp 1607319584
transform 1 0 1900 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_361
timestamp 1607319584
transform 1 0 1932 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_17
timestamp 1607319584
transform 1 0 2028 0 1 305
box -2 -3 34 103
use FILL  FILL_3_3_0
timestamp 1607319584
transform -1 0 2068 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1607319584
transform -1 0 2076 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_18
timestamp 1607319584
transform -1 0 2108 0 1 305
box -2 -3 34 103
use INVX1  INVX1_468
timestamp 1607319584
transform -1 0 2124 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_61
timestamp 1607319584
transform 1 0 2124 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_62
timestamp 1607319584
transform -1 0 2188 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_383
timestamp 1607319584
transform 1 0 2188 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_52
timestamp 1607319584
transform -1 0 2316 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_51
timestamp 1607319584
transform 1 0 2316 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_14
timestamp 1607319584
transform 1 0 2348 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1607319584
transform 1 0 2380 0 1 305
box -2 -3 34 103
use INVX1  INVX1_84
timestamp 1607319584
transform 1 0 2412 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_359
timestamp 1607319584
transform 1 0 2428 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_248
timestamp 1607319584
transform 1 0 2524 0 1 305
box -2 -3 98 103
use FILL  FILL_3_4_0
timestamp 1607319584
transform 1 0 2620 0 1 305
box -2 -3 10 103
use FILL  FILL_3_4_1
timestamp 1607319584
transform 1 0 2628 0 1 305
box -2 -3 10 103
use INVX1  INVX1_459
timestamp 1607319584
transform 1 0 2636 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_1247
timestamp 1607319584
transform 1 0 2652 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1569
timestamp 1607319584
transform 1 0 2684 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1568
timestamp 1607319584
transform -1 0 2748 0 1 305
box -2 -3 34 103
use INVX1  INVX1_332
timestamp 1607319584
transform 1 0 2748 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_1544
timestamp 1607319584
transform 1 0 2764 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1543
timestamp 1607319584
transform 1 0 2796 0 1 305
box -2 -3 34 103
use INVX1  INVX1_203
timestamp 1607319584
transform 1 0 2828 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_210
timestamp 1607319584
transform 1 0 2844 0 1 305
box -2 -3 98 103
use INVX1  INVX1_331
timestamp 1607319584
transform 1 0 2940 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_1524
timestamp 1607319584
transform -1 0 2988 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1570
timestamp 1607319584
transform 1 0 2988 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1571
timestamp 1607319584
transform -1 0 3052 0 1 305
box -2 -3 34 103
use FILL  FILL_3_5_0
timestamp 1607319584
transform 1 0 3052 0 1 305
box -2 -3 10 103
use FILL  FILL_3_5_1
timestamp 1607319584
transform 1 0 3060 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_249
timestamp 1607319584
transform 1 0 3068 0 1 305
box -2 -3 98 103
use INVX1  INVX1_395
timestamp 1607319584
transform 1 0 3164 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_215
timestamp 1607319584
transform 1 0 3180 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1534
timestamp 1607319584
transform 1 0 3276 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1533
timestamp 1607319584
transform -1 0 3340 0 1 305
box -2 -3 34 103
use INVX1  INVX1_201
timestamp 1607319584
transform -1 0 3356 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_202
timestamp 1607319584
transform 1 0 3356 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1508
timestamp 1607319584
transform -1 0 3484 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1491
timestamp 1607319584
transform -1 0 3516 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1492
timestamp 1607319584
transform -1 0 3548 0 1 305
box -2 -3 34 103
use INVX1  INVX1_394
timestamp 1607319584
transform 1 0 3548 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_1182
timestamp 1607319584
transform 1 0 3564 0 1 305
box -2 -3 34 103
use INVX1  INVX1_329
timestamp 1607319584
transform 1 0 3596 0 1 305
box -2 -3 18 103
use FILL  FILL_3_6_0
timestamp 1607319584
transform 1 0 3612 0 1 305
box -2 -3 10 103
use FILL  FILL_3_6_1
timestamp 1607319584
transform 1 0 3620 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_1497
timestamp 1607319584
transform 1 0 3628 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1498
timestamp 1607319584
transform 1 0 3660 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_197
timestamp 1607319584
transform -1 0 3788 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_1506
timestamp 1607319584
transform 1 0 3788 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1505
timestamp 1607319584
transform 1 0 3820 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1489
timestamp 1607319584
transform 1 0 3852 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_98
timestamp 1607319584
transform 1 0 3884 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_342
timestamp 1607319584
transform 1 0 3916 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_201
timestamp 1607319584
transform 1 0 3940 0 1 305
box -2 -3 98 103
use BUFX4  BUFX4_462
timestamp 1607319584
transform 1 0 4036 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_898
timestamp 1607319584
transform -1 0 4164 0 1 305
box -2 -3 98 103
use FILL  FILL_3_7_0
timestamp 1607319584
transform -1 0 4172 0 1 305
box -2 -3 10 103
use FILL  FILL_3_7_1
timestamp 1607319584
transform -1 0 4180 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_677
timestamp 1607319584
transform -1 0 4212 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_678
timestamp 1607319584
transform -1 0 4244 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_908
timestamp 1607319584
transform -1 0 4340 0 1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_151
timestamp 1607319584
transform 1 0 4340 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_187
timestamp 1607319584
transform 1 0 4372 0 1 305
box -2 -3 26 103
use INVX1  INVX1_373
timestamp 1607319584
transform 1 0 4396 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_902
timestamp 1607319584
transform -1 0 4508 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_685
timestamp 1607319584
transform -1 0 4540 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_686
timestamp 1607319584
transform -1 0 4572 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_184
timestamp 1607319584
transform 1 0 4572 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_148
timestamp 1607319584
transform -1 0 4628 0 1 305
box -2 -3 34 103
use FILL  FILL_3_8_0
timestamp 1607319584
transform -1 0 4636 0 1 305
box -2 -3 10 103
use FILL  FILL_3_8_1
timestamp 1607319584
transform -1 0 4644 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_944
timestamp 1607319584
transform -1 0 4740 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_178
timestamp 1607319584
transform -1 0 4764 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_143
timestamp 1607319584
transform -1 0 4796 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_17
timestamp 1607319584
transform 1 0 4796 0 1 305
box -2 -3 50 103
use INVX1  INVX1_181
timestamp 1607319584
transform -1 0 4860 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_16
timestamp 1607319584
transform 1 0 4860 0 1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_913
timestamp 1607319584
transform -1 0 5004 0 1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_144
timestamp 1607319584
transform 1 0 5004 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_180
timestamp 1607319584
transform 1 0 5036 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_155
timestamp 1607319584
transform 1 0 5060 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_193
timestamp 1607319584
transform -1 0 5116 0 1 305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_101
timestamp 1607319584
transform -1 0 5188 0 1 305
box -2 -3 74 103
use FILL  FILL_4_1
timestamp 1607319584
transform 1 0 5188 0 1 305
box -2 -3 10 103
use BUFX4  BUFX4_341
timestamp 1607319584
transform -1 0 36 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_428
timestamp 1607319584
transform -1 0 68 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_427
timestamp 1607319584
transform -1 0 100 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_336
timestamp 1607319584
transform 1 0 100 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_450
timestamp 1607319584
transform 1 0 132 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_449
timestamp 1607319584
transform 1 0 164 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_673
timestamp 1607319584
transform 1 0 196 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_55
timestamp 1607319584
transform 1 0 292 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_695
timestamp 1607319584
transform 1 0 308 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_494
timestamp 1607319584
transform 1 0 404 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_493
timestamp 1607319584
transform -1 0 468 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_265
timestamp 1607319584
transform -1 0 492 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1607319584
transform 1 0 492 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1607319584
transform 1 0 500 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_349
timestamp 1607319584
transform 1 0 508 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1699
timestamp 1607319584
transform 1 0 604 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_326
timestamp 1607319584
transform -1 0 660 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_675
timestamp 1607319584
transform 1 0 660 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_454
timestamp 1607319584
transform 1 0 756 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_453
timestamp 1607319584
transform -1 0 820 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_477
timestamp 1607319584
transform -1 0 852 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_340
timestamp 1607319584
transform -1 0 884 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_454
timestamp 1607319584
transform -1 0 908 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_661
timestamp 1607319584
transform -1 0 932 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_56
timestamp 1607319584
transform 1 0 932 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_1148
timestamp 1607319584
transform 1 0 948 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_593
timestamp 1607319584
transform -1 0 1004 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_210
timestamp 1607319584
transform -1 0 1020 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_570
timestamp 1607319584
transform -1 0 1044 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_1_0
timestamp 1607319584
transform -1 0 1052 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1607319584
transform -1 0 1060 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_844
timestamp 1607319584
transform -1 0 1092 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_346
timestamp 1607319584
transform 1 0 1092 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_294
timestamp 1607319584
transform -1 0 1212 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_359
timestamp 1607319584
transform 1 0 1212 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_935
timestamp 1607319584
transform -1 0 1276 0 -1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_28
timestamp 1607319584
transform 1 0 1276 0 -1 505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_340
timestamp 1607319584
transform -1 0 1444 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_365
timestamp 1607319584
transform -1 0 1468 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_1680
timestamp 1607319584
transform -1 0 1500 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1681
timestamp 1607319584
transform -1 0 1532 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_368
timestamp 1607319584
transform -1 0 1564 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_2_0
timestamp 1607319584
transform -1 0 1572 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1607319584
transform -1 0 1580 0 -1 505
box -2 -3 10 103
use BUFX4  BUFX4_370
timestamp 1607319584
transform -1 0 1612 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_381
timestamp 1607319584
transform -1 0 1708 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_57
timestamp 1607319584
transform -1 0 1740 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_58
timestamp 1607319584
transform -1 0 1772 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_155
timestamp 1607319584
transform 1 0 1772 0 -1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_27
timestamp 1607319584
transform 1 0 1820 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1607319584
transform -1 0 1884 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_366
timestamp 1607319584
transform -1 0 1980 0 -1 505
box -2 -3 98 103
use BUFX4  BUFX4_367
timestamp 1607319584
transform -1 0 2012 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_351
timestamp 1607319584
transform 1 0 2012 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_352
timestamp 1607319584
transform -1 0 2076 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_3_0
timestamp 1607319584
transform 1 0 2076 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1607319584
transform 1 0 2084 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_612
timestamp 1607319584
transform 1 0 2092 0 -1 505
box -2 -3 98 103
use BUFX4  BUFX4_313
timestamp 1607319584
transform 1 0 2188 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_354
timestamp 1607319584
transform 1 0 2220 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_4
timestamp 1607319584
transform 1 0 2316 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_3
timestamp 1607319584
transform -1 0 2380 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_295
timestamp 1607319584
transform -1 0 2404 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_296
timestamp 1607319584
transform -1 0 2428 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_872
timestamp 1607319584
transform 1 0 2428 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1607319584
transform 1 0 2460 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_640
timestamp 1607319584
transform -1 0 2516 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_375
timestamp 1607319584
transform 1 0 2516 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_4_0
timestamp 1607319584
transform -1 0 2620 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_4_1
timestamp 1607319584
transform -1 0 2628 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_45
timestamp 1607319584
transform -1 0 2660 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_700
timestamp 1607319584
transform 1 0 2660 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_256
timestamp 1607319584
transform 1 0 2684 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1585
timestamp 1607319584
transform 1 0 2780 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_701
timestamp 1607319584
transform -1 0 2836 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_1584
timestamp 1607319584
transform -1 0 2868 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_238
timestamp 1607319584
transform -1 0 2964 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1523
timestamp 1607319584
transform 1 0 2964 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_563
timestamp 1607319584
transform -1 0 3020 0 -1 505
box -2 -3 26 103
use BUFX4  BUFX4_93
timestamp 1607319584
transform 1 0 3020 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_96
timestamp 1607319584
transform 1 0 3052 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_5_0
timestamp 1607319584
transform 1 0 3084 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_5_1
timestamp 1607319584
transform 1 0 3092 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_1578
timestamp 1607319584
transform 1 0 3100 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1579
timestamp 1607319584
transform -1 0 3164 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_253
timestamp 1607319584
transform 1 0 3164 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_214
timestamp 1607319584
transform 1 0 3260 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_330
timestamp 1607319584
transform 1 0 3356 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_561
timestamp 1607319584
transform -1 0 3396 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_1183
timestamp 1607319584
transform 1 0 3396 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_631
timestamp 1607319584
transform 1 0 3428 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_356
timestamp 1607319584
transform -1 0 3476 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_284
timestamp 1607319584
transform -1 0 3508 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_239
timestamp 1607319584
transform -1 0 3604 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_6_0
timestamp 1607319584
transform 1 0 3604 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_6_1
timestamp 1607319584
transform 1 0 3612 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_560
timestamp 1607319584
transform 1 0 3620 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_1515
timestamp 1607319584
transform 1 0 3644 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_206
timestamp 1607319584
transform -1 0 3772 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1516
timestamp 1607319584
transform -1 0 3804 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1490
timestamp 1607319584
transform 1 0 3804 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_193
timestamp 1607319584
transform 1 0 3836 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_181
timestamp 1607319584
transform 1 0 3932 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_145
timestamp 1607319584
transform -1 0 3988 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_922
timestamp 1607319584
transform -1 0 4084 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_469
timestamp 1607319584
transform 1 0 4084 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_7_0
timestamp 1607319584
transform 1 0 4108 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_7_1
timestamp 1607319584
transform 1 0 4116 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_829
timestamp 1607319584
transform 1 0 4124 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_270
timestamp 1607319584
transform -1 0 4244 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_219
timestamp 1607319584
transform -1 0 4276 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_942
timestamp 1607319584
transform 1 0 4276 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_746
timestamp 1607319584
transform -1 0 4396 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_400
timestamp 1607319584
transform 1 0 4396 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_158
timestamp 1607319584
transform 1 0 4420 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_196
timestamp 1607319584
transform -1 0 4476 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_401
timestamp 1607319584
transform 1 0 4476 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_220
timestamp 1607319584
transform 1 0 4500 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_271
timestamp 1607319584
transform -1 0 4556 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_911
timestamp 1607319584
transform 1 0 4556 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_8_0
timestamp 1607319584
transform 1 0 4652 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_8_1
timestamp 1607319584
transform 1 0 4660 0 -1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_198
timestamp 1607319584
transform 1 0 4668 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_160
timestamp 1607319584
transform -1 0 4724 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_540
timestamp 1607319584
transform -1 0 4748 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_924
timestamp 1607319584
transform -1 0 4844 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_956
timestamp 1607319584
transform -1 0 4940 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_923
timestamp 1607319584
transform -1 0 5036 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_182
timestamp 1607319584
transform 1 0 5036 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_146
timestamp 1607319584
transform -1 0 5092 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_402
timestamp 1607319584
transform 1 0 5092 0 -1 505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_86
timestamp 1607319584
transform -1 0 5188 0 -1 505
box -2 -3 74 103
use FILL  FILL_5_1
timestamp 1607319584
transform -1 0 5196 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_676
timestamp 1607319584
transform 1 0 4 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_456
timestamp 1607319584
transform 1 0 100 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_455
timestamp 1607319584
transform -1 0 164 0 1 505
box -2 -3 34 103
use INVX1  INVX1_358
timestamp 1607319584
transform 1 0 164 0 1 505
box -2 -3 18 103
use INVX1  INVX1_231
timestamp 1607319584
transform 1 0 180 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_444
timestamp 1607319584
transform 1 0 196 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_443
timestamp 1607319584
transform -1 0 260 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_670
timestamp 1607319584
transform -1 0 356 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_345
timestamp 1607319584
transform 1 0 356 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_703
timestamp 1607319584
transform 1 0 452 0 1 505
box -2 -3 98 103
use FILL  FILL_5_0_0
timestamp 1607319584
transform 1 0 548 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1607319584
transform 1 0 556 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_425
timestamp 1607319584
transform 1 0 564 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_426
timestamp 1607319584
transform -1 0 628 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1698
timestamp 1607319584
transform -1 0 660 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_661
timestamp 1607319584
transform 1 0 660 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_501
timestamp 1607319584
transform -1 0 780 0 1 505
box -2 -3 26 103
use INVX1  INVX1_274
timestamp 1607319584
transform 1 0 780 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_1062
timestamp 1607319584
transform -1 0 828 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1674
timestamp 1607319584
transform -1 0 860 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1019
timestamp 1607319584
transform 1 0 860 0 1 505
box -2 -3 34 103
use INVX1  INVX1_424
timestamp 1607319584
transform 1 0 892 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_843
timestamp 1607319584
transform -1 0 940 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_266
timestamp 1607319584
transform 1 0 940 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_1211
timestamp 1607319584
transform -1 0 1020 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1126
timestamp 1607319584
transform -1 0 1052 0 1 505
box -2 -3 34 103
use FILL  FILL_5_1_0
timestamp 1607319584
transform 1 0 1052 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1607319584
transform 1 0 1060 0 1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_38
timestamp 1607319584
transform 1 0 1068 0 1 505
box -2 -3 50 103
use BUFX4  BUFX4_403
timestamp 1607319584
transform -1 0 1148 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_406
timestamp 1607319584
transform -1 0 1180 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_870
timestamp 1607319584
transform 1 0 1180 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_310
timestamp 1607319584
transform -1 0 1244 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_107
timestamp 1607319584
transform 1 0 1244 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_317
timestamp 1607319584
transform 1 0 1292 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_318
timestamp 1607319584
transform -1 0 1356 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_595
timestamp 1607319584
transform -1 0 1452 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_936
timestamp 1607319584
transform -1 0 1484 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_502
timestamp 1607319584
transform -1 0 1508 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_307
timestamp 1607319584
transform -1 0 1540 0 1 505
box -2 -3 34 103
use FILL  FILL_5_2_0
timestamp 1607319584
transform 1 0 1540 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1607319584
transform 1 0 1548 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_384
timestamp 1607319584
transform 1 0 1556 0 1 505
box -2 -3 98 103
use INVX1  INVX1_276
timestamp 1607319584
transform 1 0 1652 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_64
timestamp 1607319584
transform -1 0 1700 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_63
timestamp 1607319584
transform -1 0 1732 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_382
timestamp 1607319584
transform 1 0 1732 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_59
timestamp 1607319584
transform 1 0 1828 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_60
timestamp 1607319584
transform -1 0 1892 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_614
timestamp 1607319584
transform 1 0 1892 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_355
timestamp 1607319584
transform -1 0 2020 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_356
timestamp 1607319584
transform -1 0 2052 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_367
timestamp 1607319584
transform 1 0 2052 0 1 505
box -2 -3 34 103
use FILL  FILL_5_3_0
timestamp 1607319584
transform -1 0 2092 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1607319584
transform -1 0 2100 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_368
timestamp 1607319584
transform -1 0 2132 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_620
timestamp 1607319584
transform 1 0 2132 0 1 505
box -2 -3 98 103
use INVX1  INVX1_467
timestamp 1607319584
transform 1 0 2228 0 1 505
box -2 -3 18 103
use BUFX4  BUFX4_312
timestamp 1607319584
transform 1 0 2244 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1703
timestamp 1607319584
transform 1 0 2276 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1702
timestamp 1607319584
transform 1 0 2308 0 1 505
box -2 -3 34 103
use INVX1  INVX1_83
timestamp 1607319584
transform 1 0 2340 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_351
timestamp 1607319584
transform 1 0 2356 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_34
timestamp 1607319584
transform 1 0 2452 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_369
timestamp 1607319584
transform 1 0 2484 0 1 505
box -2 -3 98 103
use FILL  FILL_5_4_0
timestamp 1607319584
transform -1 0 2588 0 1 505
box -2 -3 10 103
use FILL  FILL_5_4_1
timestamp 1607319584
transform -1 0 2596 0 1 505
box -2 -3 10 103
use INVX1  INVX1_403
timestamp 1607319584
transform -1 0 2612 0 1 505
box -2 -3 18 103
use INVX1  INVX1_404
timestamp 1607319584
transform -1 0 2628 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_240
timestamp 1607319584
transform -1 0 2724 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_357
timestamp 1607319584
transform 1 0 2724 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_285
timestamp 1607319584
transform -1 0 2780 0 1 505
box -2 -3 34 103
use INVX1  INVX1_460
timestamp 1607319584
transform 1 0 2780 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_1248
timestamp 1607319584
transform 1 0 2796 0 1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_66
timestamp 1607319584
transform 1 0 2828 0 1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_355
timestamp 1607319584
transform 1 0 2900 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_283
timestamp 1607319584
transform -1 0 2956 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1120
timestamp 1607319584
transform 1 0 2956 0 1 505
box -2 -3 34 103
use INVX1  INVX1_74
timestamp 1607319584
transform 1 0 2988 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_236
timestamp 1607319584
transform -1 0 3100 0 1 505
box -2 -3 98 103
use FILL  FILL_5_5_0
timestamp 1607319584
transform 1 0 3100 0 1 505
box -2 -3 10 103
use FILL  FILL_5_5_1
timestamp 1607319584
transform 1 0 3108 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_353
timestamp 1607319584
transform 1 0 3116 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_281
timestamp 1607319584
transform -1 0 3172 0 1 505
box -2 -3 34 103
use INVX1  INVX1_15
timestamp 1607319584
transform 1 0 3172 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_1532
timestamp 1607319584
transform 1 0 3188 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_255
timestamp 1607319584
transform 1 0 3220 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1583
timestamp 1607319584
transform 1 0 3316 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1531
timestamp 1607319584
transform -1 0 3380 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1582
timestamp 1607319584
transform -1 0 3412 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1118
timestamp 1607319584
transform 1 0 3412 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1507
timestamp 1607319584
transform 1 0 3444 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_244
timestamp 1607319584
transform -1 0 3524 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_835
timestamp 1607319584
transform -1 0 3548 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_834
timestamp 1607319584
transform -1 0 3572 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_341
timestamp 1607319584
transform -1 0 3596 0 1 505
box -2 -3 26 103
use FILL  FILL_5_6_0
timestamp 1607319584
transform 1 0 3596 0 1 505
box -2 -3 10 103
use FILL  FILL_5_6_1
timestamp 1607319584
transform 1 0 3604 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_1117
timestamp 1607319584
transform 1 0 3612 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_211
timestamp 1607319584
transform 1 0 3644 0 1 505
box -2 -3 98 103
use INVX1  INVX1_393
timestamp 1607319584
transform -1 0 3756 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_1525
timestamp 1607319584
transform -1 0 3788 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1526
timestamp 1607319584
transform -1 0 3820 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1521
timestamp 1607319584
transform 1 0 3820 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_1522
timestamp 1607319584
transform 1 0 3852 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_177
timestamp 1607319584
transform -1 0 3908 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_209
timestamp 1607319584
transform -1 0 4004 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_1033
timestamp 1607319584
transform 1 0 4004 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_179
timestamp 1607319584
transform -1 0 4060 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_693
timestamp 1607319584
transform 1 0 4060 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_607
timestamp 1607319584
transform 1 0 4092 0 1 505
box -2 -3 26 103
use FILL  FILL_5_7_0
timestamp 1607319584
transform -1 0 4124 0 1 505
box -2 -3 10 103
use FILL  FILL_5_7_1
timestamp 1607319584
transform -1 0 4132 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_1161
timestamp 1607319584
transform -1 0 4164 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_694
timestamp 1607319584
transform -1 0 4196 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_533
timestamp 1607319584
transform -1 0 4220 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_140
timestamp 1607319584
transform 1 0 4220 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_112
timestamp 1607319584
transform -1 0 4276 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1607319584
transform -1 0 4372 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_174
timestamp 1607319584
transform 1 0 4372 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_969
timestamp 1607319584
transform -1 0 4428 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_175
timestamp 1607319584
transform 1 0 4428 0 1 505
box -2 -3 26 103
use INVX1  INVX1_5
timestamp 1607319584
transform -1 0 4468 0 1 505
box -2 -3 18 103
use BUFX4  BUFX4_65
timestamp 1607319584
transform -1 0 4500 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1607319584
transform 1 0 4500 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_704
timestamp 1607319584
transform 1 0 4596 0 1 505
box -2 -3 34 103
use FILL  FILL_5_8_0
timestamp 1607319584
transform 1 0 4628 0 1 505
box -2 -3 10 103
use FILL  FILL_5_8_1
timestamp 1607319584
transform 1 0 4636 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_703
timestamp 1607319584
transform 1 0 4644 0 1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_90
timestamp 1607319584
transform -1 0 4748 0 1 505
box -2 -3 74 103
use INVX1  INVX1_437
timestamp 1607319584
transform -1 0 4764 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_183
timestamp 1607319584
transform 1 0 4764 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_147
timestamp 1607319584
transform -1 0 4820 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_205
timestamp 1607319584
transform 1 0 4820 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_165
timestamp 1607319584
transform -1 0 4876 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_186
timestamp 1607319584
transform 1 0 4876 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_150
timestamp 1607319584
transform -1 0 4932 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_927
timestamp 1607319584
transform -1 0 5028 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_154
timestamp 1607319584
transform 1 0 5028 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_192
timestamp 1607319584
transform 1 0 5060 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_938
timestamp 1607319584
transform -1 0 5180 0 1 505
box -2 -3 98 103
use FILL  FILL_6_1
timestamp 1607319584
transform 1 0 5180 0 1 505
box -2 -3 10 103
use FILL  FILL_6_2
timestamp 1607319584
transform 1 0 5188 0 1 505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_96
timestamp 1607319584
transform -1 0 76 0 -1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_825
timestamp 1607319584
transform 1 0 76 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_108
timestamp 1607319584
transform 1 0 172 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1146
timestamp 1607319584
transform 1 0 204 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_591
timestamp 1607319584
transform -1 0 260 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1691
timestamp 1607319584
transform 1 0 260 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1690
timestamp 1607319584
transform 1 0 292 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_510
timestamp 1607319584
transform 1 0 324 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_509
timestamp 1607319584
transform -1 0 388 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_347
timestamp 1607319584
transform 1 0 388 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1694
timestamp 1607319584
transform 1 0 484 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1695
timestamp 1607319584
transform -1 0 548 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1607319584
transform -1 0 556 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1607319584
transform -1 0 564 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_363
timestamp 1607319584
transform -1 0 588 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_294
timestamp 1607319584
transform 1 0 588 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_337
timestamp 1607319584
transform 1 0 604 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1675
timestamp 1607319584
transform 1 0 700 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_348
timestamp 1607319584
transform 1 0 732 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1697
timestamp 1607319584
transform 1 0 828 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1696
timestamp 1607319584
transform -1 0 892 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_432
timestamp 1607319584
transform -1 0 916 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1212
timestamp 1607319584
transform 1 0 916 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_662
timestamp 1607319584
transform -1 0 972 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_385
timestamp 1607319584
transform -1 0 996 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_603
timestamp 1607319584
transform 1 0 996 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_1_0
timestamp 1607319584
transform -1 0 1100 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1607319584
transform -1 0 1108 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_333
timestamp 1607319584
transform -1 0 1140 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_380
timestamp 1607319584
transform -1 0 1164 0 -1 705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_79
timestamp 1607319584
transform 1 0 1164 0 -1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_596
timestamp 1607319584
transform 1 0 1236 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_320
timestamp 1607319584
transform 1 0 1332 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_319
timestamp 1607319584
transform -1 0 1396 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_708
timestamp 1607319584
transform -1 0 1420 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1063
timestamp 1607319584
transform 1 0 1420 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_618
timestamp 1607319584
transform 1 0 1452 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_2_0
timestamp 1607319584
transform 1 0 1548 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1607319584
transform 1 0 1556 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_364
timestamp 1607319584
transform 1 0 1564 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_363
timestamp 1607319584
transform 1 0 1596 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_503
timestamp 1607319584
transform 1 0 1628 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1064
timestamp 1607319584
transform -1 0 1684 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_448
timestamp 1607319584
transform 1 0 1684 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_347
timestamp 1607319584
transform 1 0 1708 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_348
timestamp 1607319584
transform -1 0 1772 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_610
timestamp 1607319584
transform -1 0 1868 0 -1 705
box -2 -3 98 103
use BUFX4  BUFX4_109
timestamp 1607319584
transform -1 0 1900 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_354
timestamp 1607319584
transform 1 0 1900 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_353
timestamp 1607319584
transform 1 0 1932 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_314
timestamp 1607319584
transform 1 0 1964 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_313
timestamp 1607319584
transform 1 0 1996 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_3_0
timestamp 1607319584
transform 1 0 2028 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1607319584
transform 1 0 2036 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_593
timestamp 1607319584
transform 1 0 2044 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1687
timestamp 1607319584
transform 1 0 2140 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_450
timestamp 1607319584
transform 1 0 2172 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_343
timestamp 1607319584
transform 1 0 2196 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1686
timestamp 1607319584
transform -1 0 2324 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_641
timestamp 1607319584
transform -1 0 2348 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_402
timestamp 1607319584
transform 1 0 2348 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_871
timestamp 1607319584
transform 1 0 2364 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_639
timestamp 1607319584
transform 1 0 2396 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_2
timestamp 1607319584
transform 1 0 2420 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1
timestamp 1607319584
transform 1 0 2452 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_353
timestamp 1607319584
transform 1 0 2484 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_4_0
timestamp 1607319584
transform -1 0 2588 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_4_1
timestamp 1607319584
transform -1 0 2596 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1191
timestamp 1607319584
transform -1 0 2628 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_33
timestamp 1607319584
transform -1 0 2660 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_50
timestamp 1607319584
transform 1 0 2660 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_377
timestamp 1607319584
transform 1 0 2692 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_49
timestamp 1607319584
transform -1 0 2820 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_404
timestamp 1607319584
transform 1 0 2820 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_405
timestamp 1607319584
transform 1 0 2852 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_562
timestamp 1607319584
transform -1 0 2908 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1119
timestamp 1607319584
transform -1 0 2940 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_245
timestamp 1607319584
transform 1 0 2940 0 -1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_287
timestamp 1607319584
transform -1 0 3012 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_991
timestamp 1607319584
transform 1 0 3012 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_424
timestamp 1607319584
transform -1 0 3068 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_90
timestamp 1607319584
transform -1 0 3100 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_5_0
timestamp 1607319584
transform 1 0 3100 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_5_1
timestamp 1607319584
transform 1 0 3108 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1562
timestamp 1607319584
transform 1 0 3116 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1563
timestamp 1607319584
transform -1 0 3180 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_245
timestamp 1607319584
transform 1 0 3180 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_494
timestamp 1607319584
transform -1 0 3300 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_241
timestamp 1607319584
transform 1 0 3300 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_632
timestamp 1607319584
transform -1 0 3420 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_9
timestamp 1607319584
transform 1 0 3420 0 -1 705
box -2 -3 18 103
use BUFX4  BUFX4_91
timestamp 1607319584
transform 1 0 3436 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1528
timestamp 1607319584
transform 1 0 3468 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1527
timestamp 1607319584
transform -1 0 3532 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_212
timestamp 1607319584
transform -1 0 3628 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_6_0
timestamp 1607319584
transform 1 0 3628 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_6_1
timestamp 1607319584
transform 1 0 3636 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_213
timestamp 1607319584
transform 1 0 3644 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1530
timestamp 1607319584
transform 1 0 3740 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1529
timestamp 1607319584
transform -1 0 3804 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_30
timestamp 1607319584
transform -1 0 3852 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_29
timestamp 1607319584
transform -1 0 3900 0 -1 705
box -2 -3 50 103
use NOR2X1  NOR2X1_346
timestamp 1607319584
transform 1 0 3900 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_275
timestamp 1607319584
transform -1 0 3956 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_221
timestamp 1607319584
transform 1 0 3956 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_608
timestamp 1607319584
transform 1 0 4052 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_7_0
timestamp 1607319584
transform -1 0 4084 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_7_1
timestamp 1607319584
transform -1 0 4092 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_906
timestamp 1607319584
transform -1 0 4188 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1092
timestamp 1607319584
transform -1 0 4220 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_115
timestamp 1607319584
transform 1 0 4220 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_304
timestamp 1607319584
transform -1 0 4268 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_821
timestamp 1607319584
transform -1 0 4364 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_539
timestamp 1607319584
transform 1 0 4364 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_133
timestamp 1607319584
transform 1 0 4388 0 -1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_970
timestamp 1607319584
transform 1 0 4436 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_182
timestamp 1607319584
transform -1 0 4484 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_953
timestamp 1607319584
transform -1 0 4580 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_162
timestamp 1607319584
transform -1 0 4612 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_747
timestamp 1607319584
transform 1 0 4612 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_8_0
timestamp 1607319584
transform 1 0 4636 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_8_1
timestamp 1607319584
transform 1 0 4644 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_676
timestamp 1607319584
transform 1 0 4652 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1225
timestamp 1607319584
transform -1 0 4708 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1099
timestamp 1607319584
transform -1 0 4740 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_168
timestamp 1607319584
transform -1 0 4772 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_959
timestamp 1607319584
transform 1 0 4772 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_333
timestamp 1607319584
transform 1 0 4868 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1607319584
transform -1 0 4988 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_221
timestamp 1607319584
transform 1 0 4988 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_272
timestamp 1607319584
transform -1 0 5044 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_717
timestamp 1607319584
transform 1 0 5044 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_311
timestamp 1607319584
transform -1 0 5092 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_933
timestamp 1607319584
transform -1 0 5188 0 -1 705
box -2 -3 98 103
use FILL  FILL_7_1
timestamp 1607319584
transform -1 0 5196 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_817
timestamp 1607319584
transform 1 0 4 0 1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_107
timestamp 1607319584
transform 1 0 100 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_134
timestamp 1607319584
transform -1 0 156 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_5
timestamp 1607319584
transform -1 0 204 0 1 705
box -2 -3 50 103
use NOR2X1  NOR2X1_136
timestamp 1607319584
transform 1 0 204 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_452
timestamp 1607319584
transform 1 0 228 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_342
timestamp 1607319584
transform 1 0 260 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_47
timestamp 1607319584
transform 1 0 292 0 1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_700
timestamp 1607319584
transform 1 0 364 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_504
timestamp 1607319584
transform 1 0 460 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_503
timestamp 1607319584
transform -1 0 524 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1607319584
transform 1 0 524 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1607319584
transform 1 0 532 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_511
timestamp 1607319584
transform 1 0 540 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_512
timestamp 1607319584
transform -1 0 604 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_704
timestamp 1607319584
transform 1 0 604 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_934
timestamp 1607319584
transform 1 0 700 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_220
timestamp 1607319584
transform -1 0 756 0 1 705
box -2 -3 26 103
use INVX1  INVX1_23
timestamp 1607319584
transform 1 0 756 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_202
timestamp 1607319584
transform 1 0 772 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_464
timestamp 1607319584
transform 1 0 820 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_680
timestamp 1607319584
transform 1 0 852 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_94
timestamp 1607319584
transform -1 0 972 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_998
timestamp 1607319584
transform -1 0 1004 0 1 705
box -2 -3 34 103
use INVX1  INVX1_167
timestamp 1607319584
transform 1 0 1004 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_97
timestamp 1607319584
transform -1 0 1044 0 1 705
box -2 -3 26 103
use FILL  FILL_7_1_0
timestamp 1607319584
transform 1 0 1044 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1607319584
transform 1 0 1052 0 1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_314
timestamp 1607319584
transform 1 0 1060 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_334
timestamp 1607319584
transform -1 0 1140 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_605
timestamp 1607319584
transform 1 0 1140 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_338
timestamp 1607319584
transform 1 0 1236 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_337
timestamp 1607319584
transform 1 0 1268 0 1 705
box -2 -3 34 103
use INVX1  INVX1_226
timestamp 1607319584
transform -1 0 1316 0 1 705
box -2 -3 18 103
use BUFX4  BUFX4_316
timestamp 1607319584
transform -1 0 1348 0 1 705
box -2 -3 34 103
use INVX2  INVX2_11
timestamp 1607319584
transform 1 0 1348 0 1 705
box -2 -3 18 103
use INVX1  INVX1_162
timestamp 1607319584
transform 1 0 1364 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_950
timestamp 1607319584
transform 1 0 1380 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1254
timestamp 1607319584
transform 1 0 1412 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_872
timestamp 1607319584
transform 1 0 1444 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_871
timestamp 1607319584
transform -1 0 1492 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_2
timestamp 1607319584
transform 1 0 1492 0 1 705
box -2 -3 26 103
use INVX1  INVX1_483
timestamp 1607319584
transform 1 0 1516 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_3
timestamp 1607319584
transform 1 0 1532 0 1 705
box -2 -3 26 103
use FILL  FILL_7_2_0
timestamp 1607319584
transform 1 0 1556 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1607319584
transform 1 0 1564 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_4
timestamp 1607319584
transform 1 0 1572 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_1
timestamp 1607319584
transform 1 0 1596 0 1 705
box -2 -3 26 103
use INVX2  INVX2_3
timestamp 1607319584
transform -1 0 1636 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_203
timestamp 1607319584
transform 1 0 1636 0 1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_204
timestamp 1607319584
transform 1 0 1684 0 1 705
box -2 -3 50 103
use BUFX4  BUFX4_382
timestamp 1607319584
transform -1 0 1764 0 1 705
box -2 -3 34 103
use INVX1  INVX1_99
timestamp 1607319584
transform 1 0 1764 0 1 705
box -2 -3 18 103
use INVX1  INVX1_339
timestamp 1607319584
transform -1 0 1796 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_312
timestamp 1607319584
transform -1 0 1820 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_632
timestamp 1607319584
transform -1 0 1916 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_613
timestamp 1607319584
transform 1 0 1916 0 1 705
box -2 -3 98 103
use BUFX4  BUFX4_102
timestamp 1607319584
transform -1 0 2044 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_387
timestamp 1607319584
transform -1 0 2076 0 1 705
box -2 -3 34 103
use FILL  FILL_7_3_0
timestamp 1607319584
transform 1 0 2076 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1607319584
transform 1 0 2084 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_330
timestamp 1607319584
transform 1 0 2092 0 1 705
box -2 -3 34 103
use INVX1  INVX1_50
timestamp 1607319584
transform 1 0 2124 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_601
timestamp 1607319584
transform 1 0 2140 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_329
timestamp 1607319584
transform -1 0 2268 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1015
timestamp 1607319584
transform -1 0 2300 0 1 705
box -2 -3 34 103
use INVX1  INVX1_227
timestamp 1607319584
transform -1 0 2316 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_345
timestamp 1607319584
transform 1 0 2316 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_346
timestamp 1607319584
transform -1 0 2380 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_378
timestamp 1607319584
transform 1 0 2380 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1190
timestamp 1607319584
transform 1 0 2404 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_59
timestamp 1607319584
transform -1 0 2484 0 1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_609
timestamp 1607319584
transform -1 0 2580 0 1 705
box -2 -3 98 103
use FILL  FILL_7_4_0
timestamp 1607319584
transform -1 0 2588 0 1 705
box -2 -3 10 103
use FILL  FILL_7_4_1
timestamp 1607319584
transform -1 0 2596 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_1192
timestamp 1607319584
transform -1 0 2628 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_63
timestamp 1607319584
transform -1 0 2652 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_49
timestamp 1607319584
transform -1 0 2684 0 1 705
box -2 -3 34 103
use INVX1  INVX1_22
timestamp 1607319584
transform 1 0 2684 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_585
timestamp 1607319584
transform 1 0 2700 0 1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_341
timestamp 1607319584
transform 1 0 2796 0 1 705
box -2 -3 50 103
use INVX1  INVX1_21
timestamp 1607319584
transform 1 0 2844 0 1 705
box -2 -3 18 103
use BUFX4  BUFX4_128
timestamp 1607319584
transform 1 0 2860 0 1 705
box -2 -3 34 103
use INVX1  INVX1_75
timestamp 1607319584
transform -1 0 2908 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_226
timestamp 1607319584
transform -1 0 3004 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_1540
timestamp 1607319584
transform 1 0 3004 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1539
timestamp 1607319584
transform -1 0 3068 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_149
timestamp 1607319584
transform -1 0 3116 0 1 705
box -2 -3 50 103
use FILL  FILL_7_5_0
timestamp 1607319584
transform -1 0 3124 0 1 705
box -2 -3 10 103
use FILL  FILL_7_5_1
timestamp 1607319584
transform -1 0 3132 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_837
timestamp 1607319584
transform -1 0 3156 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_836
timestamp 1607319584
transform -1 0 3180 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_839
timestamp 1607319584
transform -1 0 3204 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_459
timestamp 1607319584
transform 1 0 3204 0 1 705
box -2 -3 34 103
use INVX1  INVX1_268
timestamp 1607319584
transform 1 0 3236 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_1056
timestamp 1607319584
transform 1 0 3252 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1554
timestamp 1607319584
transform 1 0 3284 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1555
timestamp 1607319584
transform -1 0 3348 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_840
timestamp 1607319584
transform -1 0 3372 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1575
timestamp 1607319584
transform 1 0 3372 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1574
timestamp 1607319584
transform -1 0 3436 0 1 705
box -2 -3 34 103
use INVX1  INVX1_202
timestamp 1607319584
transform -1 0 3452 0 1 705
box -2 -3 18 103
use INVX1  INVX1_73
timestamp 1607319584
transform -1 0 3468 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_251
timestamp 1607319584
transform -1 0 3564 0 1 705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_76
timestamp 1607319584
transform 1 0 3564 0 1 705
box -2 -3 74 103
use FILL  FILL_7_6_0
timestamp 1607319584
transform -1 0 3644 0 1 705
box -2 -3 10 103
use FILL  FILL_7_6_1
timestamp 1607319584
transform -1 0 3652 0 1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_292
timestamp 1607319584
transform -1 0 3700 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_1181
timestamp 1607319584
transform -1 0 3732 0 1 705
box -2 -3 34 103
use INVX1  INVX1_138
timestamp 1607319584
transform 1 0 3732 0 1 705
box -2 -3 18 103
use INVX1  INVX1_266
timestamp 1607319584
transform 1 0 3748 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_21
timestamp 1607319584
transform 1 0 3764 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_492
timestamp 1607319584
transform -1 0 3836 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_331
timestamp 1607319584
transform 1 0 3836 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_905
timestamp 1607319584
transform -1 0 3892 0 1 705
box -2 -3 34 103
use INVX1  INVX1_117
timestamp 1607319584
transform -1 0 3908 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_201
timestamp 1607319584
transform -1 0 3932 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_190
timestamp 1607319584
transform -1 0 3956 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_64
timestamp 1607319584
transform 1 0 3956 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_199
timestamp 1607319584
transform -1 0 4012 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_181
timestamp 1607319584
transform 1 0 4012 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_713
timestamp 1607319584
transform -1 0 4092 0 1 705
box -2 -3 34 103
use FILL  FILL_7_7_0
timestamp 1607319584
transform 1 0 4092 0 1 705
box -2 -3 10 103
use FILL  FILL_7_7_1
timestamp 1607319584
transform 1 0 4100 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_920
timestamp 1607319584
transform 1 0 4108 0 1 705
box -2 -3 98 103
use INVX1  INVX1_502
timestamp 1607319584
transform 1 0 4204 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_618
timestamp 1607319584
transform 1 0 4220 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_145
timestamp 1607319584
transform -1 0 4276 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_480
timestamp 1607319584
transform -1 0 4300 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_1290
timestamp 1607319584
transform 1 0 4300 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_373
timestamp 1607319584
transform -1 0 4380 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_708
timestamp 1607319584
transform -1 0 4412 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_915
timestamp 1607319584
transform 1 0 4412 0 1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_19
timestamp 1607319584
transform 1 0 4508 0 1 705
box -2 -3 50 103
use NOR2X1  NOR2X1_202
timestamp 1607319584
transform 1 0 4556 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_188
timestamp 1607319584
transform -1 0 4604 0 1 705
box -2 -3 26 103
use INVX1  INVX1_503
timestamp 1607319584
transform -1 0 4620 0 1 705
box -2 -3 18 103
use FILL  FILL_7_8_0
timestamp 1607319584
transform -1 0 4628 0 1 705
box -2 -3 10 103
use FILL  FILL_7_8_1
timestamp 1607319584
transform -1 0 4636 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_936
timestamp 1607319584
transform -1 0 4732 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_208
timestamp 1607319584
transform -1 0 4756 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_200
timestamp 1607319584
transform -1 0 4780 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_161
timestamp 1607319584
transform -1 0 4812 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_945
timestamp 1607319584
transform -1 0 4908 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_266
timestamp 1607319584
transform 1 0 4908 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_215
timestamp 1607319584
transform -1 0 4964 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1607319584
transform 1 0 4964 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_186
timestamp 1607319584
transform -1 0 5084 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_931
timestamp 1607319584
transform 1 0 5084 0 1 705
box -2 -3 98 103
use INVX1  INVX1_183
timestamp 1607319584
transform -1 0 5196 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_660
timestamp 1607319584
transform 1 0 4 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_424
timestamp 1607319584
transform 1 0 100 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_423
timestamp 1607319584
transform -1 0 164 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_674
timestamp 1607319584
transform 1 0 164 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_451
timestamp 1607319584
transform -1 0 292 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_306
timestamp 1607319584
transform 1 0 292 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_384
timestamp 1607319584
transform -1 0 348 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_333
timestamp 1607319584
transform 1 0 348 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_692
timestamp 1607319584
transform 1 0 444 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_0_0
timestamp 1607319584
transform 1 0 540 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1607319584
transform 1 0 548 0 -1 905
box -2 -3 10 103
use INVX1  INVX1_273
timestamp 1607319584
transform 1 0 556 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1061
timestamp 1607319584
transform -1 0 604 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_489
timestamp 1607319584
transform 1 0 604 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_490
timestamp 1607319584
transform -1 0 668 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_693
timestamp 1607319584
transform 1 0 668 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_808
timestamp 1607319584
transform 1 0 764 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1607319584
transform -1 0 820 0 -1 905
box -2 -3 26 103
use INVX2  INVX2_4
timestamp 1607319584
transform -1 0 836 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_463
timestamp 1607319584
transform 1 0 836 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_93
timestamp 1607319584
transform 1 0 868 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_731
timestamp 1607319584
transform -1 0 916 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_95
timestamp 1607319584
transform -1 0 940 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_96
timestamp 1607319584
transform 1 0 940 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_455
timestamp 1607319584
transform -1 0 988 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_955
timestamp 1607319584
transform -1 0 1020 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_1_0
timestamp 1607319584
transform 1 0 1020 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1607319584
transform 1 0 1028 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_604
timestamp 1607319584
transform 1 0 1036 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_336
timestamp 1607319584
transform 1 0 1132 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_335
timestamp 1607319584
transform -1 0 1196 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_449
timestamp 1607319584
transform -1 0 1220 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1014
timestamp 1607319584
transform -1 0 1252 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_597
timestamp 1607319584
transform -1 0 1348 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_322
timestamp 1607319584
transform 1 0 1348 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_321
timestamp 1607319584
transform -1 0 1412 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_401
timestamp 1607319584
transform -1 0 1444 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_598
timestamp 1607319584
transform 1 0 1444 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_323
timestamp 1607319584
transform 1 0 1540 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_2_0
timestamp 1607319584
transform -1 0 1580 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1607319584
transform -1 0 1588 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_324
timestamp 1607319584
transform -1 0 1620 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_78
timestamp 1607319584
transform 1 0 1620 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_80
timestamp 1607319584
transform 1 0 1644 0 -1 905
box -2 -3 26 103
use BUFX4  BUFX4_381
timestamp 1607319584
transform -1 0 1700 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_392
timestamp 1607319584
transform 1 0 1700 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_391
timestamp 1607319584
transform -1 0 1764 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_887
timestamp 1607319584
transform 1 0 1764 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_571
timestamp 1607319584
transform 1 0 1796 0 -1 905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_60
timestamp 1607319584
transform 1 0 1820 0 -1 905
box -2 -3 74 103
use BUFX4  BUFX4_386
timestamp 1607319584
transform 1 0 1892 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_622
timestamp 1607319584
transform 1 0 1924 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_372
timestamp 1607319584
transform 1 0 2020 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_371
timestamp 1607319584
transform -1 0 2084 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_3_0
timestamp 1607319584
transform -1 0 2092 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1607319584
transform -1 0 2100 0 -1 905
box -2 -3 10 103
use INVX8  INVX8_15
timestamp 1607319584
transform -1 0 2140 0 -1 905
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_636
timestamp 1607319584
transform -1 0 2236 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_260
timestamp 1607319584
transform -1 0 2260 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_64
timestamp 1607319584
transform 1 0 2260 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_50
timestamp 1607319584
transform -1 0 2316 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_51
timestamp 1607319584
transform 1 0 2316 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_65
timestamp 1607319584
transform -1 0 2372 0 -1 905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_22
timestamp 1607319584
transform -1 0 2444 0 -1 905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_1021
timestamp 1607319584
transform 1 0 2444 0 -1 905
box -2 -3 98 103
use BUFX4  BUFX4_123
timestamp 1607319584
transform -1 0 2572 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_286
timestamp 1607319584
transform 1 0 2572 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_4_0
timestamp 1607319584
transform -1 0 2604 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_4_1
timestamp 1607319584
transform -1 0 2612 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_863
timestamp 1607319584
transform -1 0 2644 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_351
timestamp 1607319584
transform 1 0 2644 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_279
timestamp 1607319584
transform -1 0 2700 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_234
timestamp 1607319584
transform -1 0 2796 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_242
timestamp 1607319584
transform 1 0 2796 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1557
timestamp 1607319584
transform 1 0 2892 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1556
timestamp 1607319584
transform -1 0 2956 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_76
timestamp 1607319584
transform 1 0 2956 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_864
timestamp 1607319584
transform 1 0 2972 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_229
timestamp 1607319584
transform 1 0 3004 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_5_0
timestamp 1607319584
transform 1 0 3100 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_5_1
timestamp 1607319584
transform 1 0 3108 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_1546
timestamp 1607319584
transform 1 0 3116 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1545
timestamp 1607319584
transform -1 0 3180 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1542
timestamp 1607319584
transform 1 0 3180 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1541
timestamp 1607319584
transform -1 0 3244 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_267
timestamp 1607319584
transform 1 0 3244 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1055
timestamp 1607319584
transform 1 0 3260 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_197
timestamp 1607319584
transform 1 0 3292 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_356
timestamp 1607319584
transform 1 0 3340 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_928
timestamp 1607319584
transform -1 0 3396 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_140
timestamp 1607319584
transform -1 0 3412 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1559
timestamp 1607319584
transform 1 0 3412 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1558
timestamp 1607319584
transform -1 0 3476 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_350
timestamp 1607319584
transform -1 0 3500 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_243
timestamp 1607319584
transform -1 0 3596 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_6_0
timestamp 1607319584
transform 1 0 3596 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_6_1
timestamp 1607319584
transform 1 0 3604 0 -1 905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_5
timestamp 1607319584
transform 1 0 3612 0 -1 905
box -2 -3 74 103
use BUFX4  BUFX4_410
timestamp 1607319584
transform -1 0 3716 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_344
timestamp 1607319584
transform 1 0 3716 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_273
timestamp 1607319584
transform -1 0 3772 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1054
timestamp 1607319584
transform 1 0 3772 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_332
timestamp 1607319584
transform 1 0 3804 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1607319584
transform 1 0 3828 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_217
timestamp 1607319584
transform 1 0 3924 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_268
timestamp 1607319584
transform -1 0 3980 0 -1 905
box -2 -3 26 103
use BUFX4  BUFX4_131
timestamp 1607319584
transform 1 0 3980 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_470
timestamp 1607319584
transform -1 0 4036 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1034
timestamp 1607319584
transform -1 0 4068 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_246
timestamp 1607319584
transform -1 0 4084 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_709
timestamp 1607319584
transform 1 0 4084 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_7_0
timestamp 1607319584
transform -1 0 4124 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_7_1
timestamp 1607319584
transform -1 0 4132 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_916
timestamp 1607319584
transform -1 0 4228 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_687
timestamp 1607319584
transform 1 0 4228 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_472
timestamp 1607319584
transform 1 0 4252 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1042
timestamp 1607319584
transform -1 0 4308 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1607319584
transform -1 0 4404 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_222
timestamp 1607319584
transform 1 0 4404 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_273
timestamp 1607319584
transform -1 0 4460 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_609
timestamp 1607319584
transform 1 0 4460 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_20
timestamp 1607319584
transform 1 0 4484 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_549
timestamp 1607319584
transform 1 0 4532 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_18
timestamp 1607319584
transform 1 0 4556 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_1291
timestamp 1607319584
transform 1 0 4604 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_8_0
timestamp 1607319584
transform 1 0 4636 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_8_1
timestamp 1607319584
transform 1 0 4644 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_720
timestamp 1607319584
transform 1 0 4652 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_189
timestamp 1607319584
transform -1 0 4708 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_189
timestamp 1607319584
transform -1 0 4732 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_152
timestamp 1607319584
transform -1 0 4764 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_929
timestamp 1607319584
transform -1 0 4860 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_677
timestamp 1607319584
transform 1 0 4860 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_955
timestamp 1607319584
transform 1 0 4884 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1309
timestamp 1607319584
transform 1 0 4980 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_254
timestamp 1607319584
transform -1 0 5028 0 -1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1607319584
transform -1 0 5124 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_971
timestamp 1607319584
transform -1 0 5156 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_715
timestamp 1607319584
transform 1 0 5156 0 -1 905
box -2 -3 34 103
use FILL  FILL_9_1
timestamp 1607319584
transform -1 0 5196 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_664
timestamp 1607319584
transform 1 0 4 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_665
timestamp 1607319584
transform 1 0 100 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_434
timestamp 1607319584
transform 1 0 196 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_433
timestamp 1607319584
transform -1 0 260 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_663
timestamp 1607319584
transform -1 0 356 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_430
timestamp 1607319584
transform 1 0 356 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_429
timestamp 1607319584
transform -1 0 420 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_379
timestamp 1607319584
transform 1 0 420 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_488
timestamp 1607319584
transform 1 0 444 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_487
timestamp 1607319584
transform 1 0 476 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_500
timestamp 1607319584
transform -1 0 532 0 1 905
box -2 -3 26 103
use FILL  FILL_9_0_0
timestamp 1607319584
transform -1 0 540 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1607319584
transform -1 0 548 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_325
timestamp 1607319584
transform -1 0 644 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1670
timestamp 1607319584
transform -1 0 676 0 1 905
box -2 -3 34 103
use INVX1  INVX1_232
timestamp 1607319584
transform 1 0 676 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_339
timestamp 1607319584
transform -1 0 724 0 1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_6
timestamp 1607319584
transform 1 0 724 0 1 905
box -2 -3 74 103
use INVX1  INVX1_296
timestamp 1607319584
transform 1 0 796 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_479
timestamp 1607319584
transform 1 0 812 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_480
timestamp 1607319584
transform -1 0 876 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_688
timestamp 1607319584
transform 1 0 876 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1020
timestamp 1607319584
transform -1 0 1004 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1607319584
transform 1 0 1004 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1607319584
transform 1 0 1012 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_607
timestamp 1607319584
transform 1 0 1020 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_342
timestamp 1607319584
transform 1 0 1116 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_341
timestamp 1607319584
transform -1 0 1180 0 1 905
box -2 -3 34 103
use INVX8  INVX8_14
timestamp 1607319584
transform -1 0 1220 0 1 905
box -2 -3 42 103
use INVX1  INVX1_290
timestamp 1607319584
transform -1 0 1236 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_326
timestamp 1607319584
transform 1 0 1236 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_599
timestamp 1607319584
transform 1 0 1268 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_325
timestamp 1607319584
transform -1 0 1396 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_79
timestamp 1607319584
transform -1 0 1420 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_77
timestamp 1607319584
transform 1 0 1420 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_10
timestamp 1607319584
transform 1 0 1444 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_82
timestamp 1607319584
transform 1 0 1476 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_81
timestamp 1607319584
transform 1 0 1500 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_405
timestamp 1607319584
transform 1 0 1524 0 1 905
box -2 -3 34 103
use FILL  FILL_9_2_0
timestamp 1607319584
transform -1 0 1564 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1607319584
transform -1 0 1572 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_406
timestamp 1607319584
transform -1 0 1604 0 1 905
box -2 -3 34 103
use INVX1  INVX1_354
timestamp 1607319584
transform 1 0 1604 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_639
timestamp 1607319584
transform -1 0 1716 0 1 905
box -2 -3 98 103
use INVX1  INVX1_484
timestamp 1607319584
transform -1 0 1732 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_169
timestamp 1607319584
transform -1 0 1764 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1127
timestamp 1607319584
transform 1 0 1764 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_396
timestamp 1607319584
transform 1 0 1796 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_395
timestamp 1607319584
transform 1 0 1828 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_634
timestamp 1607319584
transform -1 0 1956 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_369
timestamp 1607319584
transform 1 0 1956 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_370
timestamp 1607319584
transform -1 0 2020 0 1 905
box -2 -3 34 103
use INVX1  INVX1_291
timestamp 1607319584
transform 1 0 2020 0 1 905
box -2 -3 18 103
use FILL  FILL_9_3_0
timestamp 1607319584
transform -1 0 2044 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1607319584
transform -1 0 2052 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_621
timestamp 1607319584
transform -1 0 2148 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_399
timestamp 1607319584
transform -1 0 2180 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_400
timestamp 1607319584
transform -1 0 2212 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_838
timestamp 1607319584
transform 1 0 2212 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_586
timestamp 1607319584
transform -1 0 2340 0 1 905
box -2 -3 98 103
use INVX1  INVX1_51
timestamp 1607319584
transform -1 0 2356 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_587
timestamp 1607319584
transform 1 0 2356 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_191
timestamp 1607319584
transform 1 0 2452 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_235
timestamp 1607319584
transform -1 0 2508 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_379
timestamp 1607319584
transform -1 0 2532 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_113
timestamp 1607319584
transform -1 0 2564 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_424
timestamp 1607319584
transform 1 0 2564 0 1 905
box -2 -3 34 103
use FILL  FILL_9_4_0
timestamp 1607319584
transform 1 0 2596 0 1 905
box -2 -3 10 103
use FILL  FILL_9_4_1
timestamp 1607319584
transform 1 0 2604 0 1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_299
timestamp 1607319584
transform 1 0 2612 0 1 905
box -2 -3 50 103
use BUFX4  BUFX4_17
timestamp 1607319584
transform 1 0 2660 0 1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_10
timestamp 1607319584
transform 1 0 2692 0 1 905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_237
timestamp 1607319584
transform 1 0 2764 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_282
timestamp 1607319584
transform 1 0 2860 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_354
timestamp 1607319584
transform 1 0 2892 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_342
timestamp 1607319584
transform -1 0 2964 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_53
timestamp 1607319584
transform 1 0 2964 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_493
timestamp 1607319584
transform -1 0 3036 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_227
timestamp 1607319584
transform 1 0 3036 0 1 905
box -2 -3 98 103
use FILL  FILL_9_5_0
timestamp 1607319584
transform -1 0 3140 0 1 905
box -2 -3 10 103
use FILL  FILL_9_5_1
timestamp 1607319584
transform -1 0 3148 0 1 905
box -2 -3 10 103
use INVX1  INVX1_139
timestamp 1607319584
transform -1 0 3164 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_247
timestamp 1607319584
transform 1 0 3164 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1567
timestamp 1607319584
transform 1 0 3260 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1566
timestamp 1607319584
transform -1 0 3324 0 1 905
box -2 -3 34 103
use INVX1  INVX1_396
timestamp 1607319584
transform 1 0 3324 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1184
timestamp 1607319584
transform 1 0 3340 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_293
timestamp 1607319584
transform -1 0 3420 0 1 905
box -2 -3 50 103
use BUFX4  BUFX4_92
timestamp 1607319584
transform 1 0 3420 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1513
timestamp 1607319584
transform 1 0 3452 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1514
timestamp 1607319584
transform -1 0 3516 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_205
timestamp 1607319584
transform 1 0 3516 0 1 905
box -2 -3 98 103
use FILL  FILL_9_6_0
timestamp 1607319584
transform 1 0 3612 0 1 905
box -2 -3 10 103
use FILL  FILL_9_6_1
timestamp 1607319584
transform 1 0 3620 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_219
timestamp 1607319584
transform 1 0 3628 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_906
timestamp 1607319584
transform 1 0 3724 0 1 905
box -2 -3 34 103
use INVX1  INVX1_118
timestamp 1607319584
transform -1 0 3772 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_707
timestamp 1607319584
transform 1 0 3772 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_247
timestamp 1607319584
transform 1 0 3804 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_914
timestamp 1607319584
transform -1 0 3924 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_182
timestamp 1607319584
transform 1 0 3924 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_402
timestamp 1607319584
transform -1 0 3980 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_850
timestamp 1607319584
transform -1 0 4012 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_273
timestamp 1607319584
transform -1 0 4036 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_267
timestamp 1607319584
transform 1 0 4036 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_216
timestamp 1607319584
transform -1 0 4092 0 1 905
box -2 -3 34 103
use FILL  FILL_9_7_0
timestamp 1607319584
transform -1 0 4100 0 1 905
box -2 -3 10 103
use FILL  FILL_9_7_1
timestamp 1607319584
transform -1 0 4108 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1607319584
transform -1 0 4204 0 1 905
box -2 -3 98 103
use INVX1  INVX1_62
timestamp 1607319584
transform -1 0 4220 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1607319584
transform -1 0 4316 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1306
timestamp 1607319584
transform 1 0 4316 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_767
timestamp 1607319584
transform -1 0 4372 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_177
timestamp 1607319584
transform 1 0 4372 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_1106
timestamp 1607319584
transform -1 0 4428 0 1 905
box -2 -3 34 103
use INVX1  INVX1_318
timestamp 1607319584
transform -1 0 4444 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_1310
timestamp 1607319584
transform 1 0 4444 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1607319584
transform -1 0 4572 0 1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_18
timestamp 1607319584
transform 1 0 4572 0 1 905
box -2 -3 74 103
use FILL  FILL_9_8_0
timestamp 1607319584
transform -1 0 4652 0 1 905
box -2 -3 10 103
use FILL  FILL_9_8_1
timestamp 1607319584
transform -1 0 4660 0 1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_86
timestamp 1607319584
transform -1 0 4708 0 1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_908
timestamp 1607319584
transform 1 0 4708 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_721
timestamp 1607319584
transform -1 0 4772 0 1 905
box -2 -3 34 103
use INVX1  INVX1_120
timestamp 1607319584
transform -1 0 4788 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_946
timestamp 1607319584
transform 1 0 4788 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_907
timestamp 1607319584
transform -1 0 4916 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_164
timestamp 1607319584
transform 1 0 4916 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_204
timestamp 1607319584
transform -1 0 4972 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_403
timestamp 1607319584
transform -1 0 4996 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_770
timestamp 1607319584
transform -1 0 5020 0 1 905
box -2 -3 26 103
use INVX1  INVX1_119
timestamp 1607319584
transform -1 0 5036 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_930
timestamp 1607319584
transform -1 0 5132 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_714
timestamp 1607319584
transform 1 0 5132 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_183
timestamp 1607319584
transform 1 0 5164 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1607319584
transform 1 0 5188 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_696
timestamp 1607319584
transform 1 0 4 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_432
timestamp 1607319584
transform -1 0 132 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_431
timestamp 1607319584
transform -1 0 164 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_488
timestamp 1607319584
transform 1 0 164 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_495
timestamp 1607319584
transform -1 0 212 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_496
timestamp 1607319584
transform -1 0 244 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_691
timestamp 1607319584
transform 1 0 244 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_486
timestamp 1607319584
transform 1 0 340 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_485
timestamp 1607319584
transform 1 0 372 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_440
timestamp 1607319584
transform 1 0 404 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_668
timestamp 1607319584
transform 1 0 436 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_0_0
timestamp 1607319584
transform -1 0 540 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1607319584
transform -1 0 548 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_439
timestamp 1607319584
transform -1 0 580 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_669
timestamp 1607319584
transform 1 0 580 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1020
timestamp 1607319584
transform 1 0 676 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_234
timestamp 1607319584
transform 1 0 772 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_190
timestamp 1607319584
transform -1 0 828 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1084
timestamp 1607319584
transform 1 0 828 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_168
timestamp 1607319584
transform 1 0 860 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_1276
timestamp 1607319584
transform 1 0 876 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_594
timestamp 1607319584
transform 1 0 908 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_453
timestamp 1607319584
transform -1 0 1028 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_730
timestamp 1607319584
transform -1 0 1052 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_1_0
timestamp 1607319584
transform 1 0 1052 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1607319584
transform 1 0 1060 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_316
timestamp 1607319584
transform 1 0 1068 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_315
timestamp 1607319584
transform -1 0 1132 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_327
timestamp 1607319584
transform 1 0 1132 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_328
timestamp 1607319584
transform -1 0 1196 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_600
timestamp 1607319584
transform 1 0 1196 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_518
timestamp 1607319584
transform -1 0 1316 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_329
timestamp 1607319584
transform 1 0 1316 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_302
timestamp 1607319584
transform -1 0 1444 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_658
timestamp 1607319584
transform 1 0 1444 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_623
timestamp 1607319584
transform -1 0 1564 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_2_0
timestamp 1607319584
transform -1 0 1572 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1607319584
transform -1 0 1580 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_373
timestamp 1607319584
transform -1 0 1612 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_374
timestamp 1607319584
transform -1 0 1644 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1142
timestamp 1607319584
transform 1 0 1644 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_587
timestamp 1607319584
transform 1 0 1676 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_606
timestamp 1607319584
transform -1 0 1796 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_339
timestamp 1607319584
transform -1 0 1828 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_340
timestamp 1607319584
transform -1 0 1860 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_313
timestamp 1607319584
transform -1 0 1884 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_572
timestamp 1607319584
transform -1 0 1908 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1128
timestamp 1607319584
transform 1 0 1908 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_251
timestamp 1607319584
transform -1 0 1988 0 -1 1105
box -2 -3 50 103
use BUFX4  BUFX4_172
timestamp 1607319584
transform -1 0 2020 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_375
timestamp 1607319584
transform 1 0 2020 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_519
timestamp 1607319584
transform -1 0 2076 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_3_0
timestamp 1607319584
transform -1 0 2084 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1607319584
transform -1 0 2092 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_376
timestamp 1607319584
transform -1 0 2124 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_624
timestamp 1607319584
transform 1 0 2124 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_709
timestamp 1607319584
transform -1 0 2244 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_383
timestamp 1607319584
transform 1 0 2244 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_384
timestamp 1607319584
transform -1 0 2308 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_628
timestamp 1607319584
transform 1 0 2308 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_382
timestamp 1607319584
transform 1 0 2404 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_381
timestamp 1607319584
transform 1 0 2436 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_164
timestamp 1607319584
transform 1 0 2468 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_952
timestamp 1607319584
transform 1 0 2484 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_119
timestamp 1607319584
transform -1 0 2564 0 -1 1105
box -2 -3 50 103
use FILL  FILL_10_4_0
timestamp 1607319584
transform -1 0 2572 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_4_1
timestamp 1607319584
transform -1 0 2580 0 -1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_120
timestamp 1607319584
transform -1 0 2628 0 -1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_118
timestamp 1607319584
transform -1 0 2676 0 -1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_949
timestamp 1607319584
transform -1 0 2708 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_218
timestamp 1607319584
transform -1 0 2732 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_579
timestamp 1607319584
transform -1 0 2828 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_187
timestamp 1607319584
transform 1 0 2828 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_231
timestamp 1607319584
transform -1 0 2884 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1017
timestamp 1607319584
transform -1 0 2980 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_197
timestamp 1607319584
transform -1 0 3012 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_254
timestamp 1607319584
transform -1 0 3044 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_171
timestamp 1607319584
transform -1 0 3076 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_227
timestamp 1607319584
transform 1 0 3076 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_5_0
timestamp 1607319584
transform -1 0 3116 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_5_1
timestamp 1607319584
transform -1 0 3124 0 -1 1105
box -2 -3 10 103
use BUFX4  BUFX4_213
timestamp 1607319584
transform -1 0 3156 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_274
timestamp 1607319584
transform 1 0 3156 0 -1 1105
box -2 -3 34 103
use INVX8  INVX8_3
timestamp 1607319584
transform 1 0 3188 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_862
timestamp 1607319584
transform 1 0 3228 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_285
timestamp 1607319584
transform 1 0 3260 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_218
timestamp 1607319584
transform -1 0 3380 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_343
timestamp 1607319584
transform 1 0 3380 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_272
timestamp 1607319584
transform -1 0 3436 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_861
timestamp 1607319584
transform 1 0 3436 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_284
timestamp 1607319584
transform -1 0 3492 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_207
timestamp 1607319584
transform 1 0 3492 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1518
timestamp 1607319584
transform 1 0 3588 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_6_0
timestamp 1607319584
transform 1 0 3620 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_6_1
timestamp 1607319584
transform 1 0 3628 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_1517
timestamp 1607319584
transform 1 0 3636 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_629
timestamp 1607319584
transform 1 0 3668 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_345
timestamp 1607319584
transform -1 0 3716 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_274
timestamp 1607319584
transform -1 0 3748 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_220
timestamp 1607319584
transform 1 0 3748 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_353
timestamp 1607319584
transform 1 0 3844 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_85
timestamp 1607319584
transform 1 0 3868 0 -1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_176
timestamp 1607319584
transform -1 0 3940 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_426
timestamp 1607319584
transform -1 0 3972 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_342
timestamp 1607319584
transform -1 0 3996 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_914
timestamp 1607319584
transform -1 0 4028 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1307
timestamp 1607319584
transform 1 0 4028 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_126
timestamp 1607319584
transform -1 0 4076 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_7_0
timestamp 1607319584
transform -1 0 4084 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_7_1
timestamp 1607319584
transform -1 0 4092 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1607319584
transform -1 0 4188 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1162
timestamp 1607319584
transform -1 0 4220 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1234
timestamp 1607319584
transform 1 0 4220 0 -1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_87
timestamp 1607319584
transform 1 0 4252 0 -1 1105
box -2 -3 74 103
use OAI21X1  OAI21X1_1312
timestamp 1607319584
transform 1 0 4324 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_446
timestamp 1607319584
transform -1 0 4372 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1607319584
transform -1 0 4468 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1607319584
transform -1 0 4564 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_610
timestamp 1607319584
transform 1 0 4564 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_167
timestamp 1607319584
transform 1 0 4588 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_207
timestamp 1607319584
transform 1 0 4620 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_8_0
timestamp 1607319584
transform -1 0 4652 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_8_1
timestamp 1607319584
transform -1 0 4660 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_958
timestamp 1607319584
transform -1 0 4756 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_16
timestamp 1607319584
transform 1 0 4756 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_334
timestamp 1607319584
transform 1 0 4788 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_134
timestamp 1607319584
transform 1 0 4812 0 -1 1105
box -2 -3 50 103
use NOR2X1  NOR2X1_203
timestamp 1607319584
transform 1 0 4860 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_954
timestamp 1607319584
transform -1 0 4980 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_972
timestamp 1607319584
transform -1 0 5012 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1607319584
transform -1 0 5108 0 -1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_14
timestamp 1607319584
transform -1 0 5180 0 -1 1105
box -2 -3 74 103
use FILL  FILL_11_1
timestamp 1607319584
transform -1 0 5188 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_2
timestamp 1607319584
transform -1 0 5196 0 -1 1105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_58
timestamp 1607319584
transform 1 0 4 0 1 1105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_690
timestamp 1607319584
transform 1 0 76 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_483
timestamp 1607319584
transform -1 0 204 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_484
timestamp 1607319584
transform -1 0 236 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_103
timestamp 1607319584
transform -1 0 252 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_337
timestamp 1607319584
transform -1 0 284 0 1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_70
timestamp 1607319584
transform 1 0 284 0 1 1105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_698
timestamp 1607319584
transform 1 0 356 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_486
timestamp 1607319584
transform 1 0 452 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_302
timestamp 1607319584
transform 1 0 468 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_230
timestamp 1607319584
transform 1 0 500 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_422
timestamp 1607319584
transform 1 0 516 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_0_0
timestamp 1607319584
transform 1 0 532 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1607319584
transform 1 0 540 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_442
timestamp 1607319584
transform 1 0 548 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_441
timestamp 1607319584
transform 1 0 580 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_867
timestamp 1607319584
transform 1 0 612 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_701
timestamp 1607319584
transform 1 0 636 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_506
timestamp 1607319584
transform 1 0 732 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_505
timestamp 1607319584
transform -1 0 796 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_524
timestamp 1607319584
transform -1 0 820 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_300
timestamp 1607319584
transform -1 0 852 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_218
timestamp 1607319584
transform -1 0 900 0 1 1105
box -2 -3 50 103
use BUFX4  BUFX4_83
timestamp 1607319584
transform -1 0 932 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_487
timestamp 1607319584
transform 1 0 932 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_170
timestamp 1607319584
transform 1 0 948 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_1018
timestamp 1607319584
transform 1 0 996 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1275
timestamp 1607319584
transform -1 0 1060 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_1_0
timestamp 1607319584
transform 1 0 1060 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1607319584
transform 1 0 1068 0 1 1105
box -2 -3 10 103
use BUFX4  BUFX4_85
timestamp 1607319584
transform 1 0 1076 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_98
timestamp 1607319584
transform 1 0 1108 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_421
timestamp 1607319584
transform -1 0 1156 0 1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_69
timestamp 1607319584
transform 1 0 1156 0 1 1105
box -2 -3 74 103
use OAI21X1  OAI21X1_1078
timestamp 1607319584
transform 1 0 1228 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_631
timestamp 1607319584
transform 1 0 1260 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_418
timestamp 1607319584
transform 1 0 1356 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_380
timestamp 1607319584
transform 1 0 1372 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_420
timestamp 1607319584
transform 1 0 1396 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_1208
timestamp 1607319584
transform 1 0 1412 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_389
timestamp 1607319584
transform -1 0 1476 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_390
timestamp 1607319584
transform -1 0 1508 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_377
timestamp 1607319584
transform 1 0 1508 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_378
timestamp 1607319584
transform -1 0 1572 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_2_0
timestamp 1607319584
transform -1 0 1580 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1607319584
transform -1 0 1588 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_625
timestamp 1607319584
transform -1 0 1684 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1271
timestamp 1607319584
transform 1 0 1684 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_726
timestamp 1607319584
transform 1 0 1716 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_71
timestamp 1607319584
transform -1 0 1788 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_888
timestamp 1607319584
transform -1 0 1820 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_100
timestamp 1607319584
transform -1 0 1836 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_380
timestamp 1607319584
transform 1 0 1836 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_379
timestamp 1607319584
transform -1 0 1900 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_414
timestamp 1607319584
transform -1 0 1932 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_626
timestamp 1607319584
transform -1 0 2028 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_380
timestamp 1607319584
transform -1 0 2060 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_3_0
timestamp 1607319584
transform 1 0 2060 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1607319584
transform 1 0 2068 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_362
timestamp 1607319584
transform 1 0 2076 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_361
timestamp 1607319584
transform 1 0 2108 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_617
timestamp 1607319584
transform -1 0 2236 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_228
timestamp 1607319584
transform -1 0 2252 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_415
timestamp 1607319584
transform 1 0 2252 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_627
timestamp 1607319584
transform -1 0 2380 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_398
timestamp 1607319584
transform 1 0 2380 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_397
timestamp 1607319584
transform 1 0 2412 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_382
timestamp 1607319584
transform 1 0 2444 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_635
timestamp 1607319584
transform -1 0 2564 0 1 1105
box -2 -3 98 103
use INVX8  INVX8_12
timestamp 1607319584
transform -1 0 2604 0 1 1105
box -2 -3 42 103
use FILL  FILL_11_4_0
timestamp 1607319584
transform -1 0 2612 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_4_1
timestamp 1607319584
transform -1 0 2620 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_307
timestamp 1607319584
transform -1 0 2652 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_26
timestamp 1607319584
transform -1 0 2700 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_807
timestamp 1607319584
transform 1 0 2700 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_161
timestamp 1607319584
transform -1 0 2748 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_229
timestamp 1607319584
transform 1 0 2748 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_186
timestamp 1607319584
transform -1 0 2804 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1009
timestamp 1607319584
transform -1 0 2900 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_258
timestamp 1607319584
transform -1 0 2932 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_280
timestamp 1607319584
transform 1 0 2932 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_352
timestamp 1607319584
transform -1 0 2988 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_235
timestamp 1607319584
transform 1 0 2988 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_355
timestamp 1607319584
transform -1 0 3108 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_5_0
timestamp 1607319584
transform -1 0 3116 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_5_1
timestamp 1607319584
transform -1 0 3124 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_927
timestamp 1607319584
transform -1 0 3156 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1607319584
transform -1 0 3172 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_54
timestamp 1607319584
transform -1 0 3220 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_52
timestamp 1607319584
transform -1 0 3268 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_246
timestamp 1607319584
transform -1 0 3316 0 1 1105
box -2 -3 50 103
use BUFX4  BUFX4_303
timestamp 1607319584
transform -1 0 3348 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_101
timestamp 1607319584
transform 1 0 3348 0 1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_204
timestamp 1607319584
transform -1 0 3492 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_1512
timestamp 1607319584
transform 1 0 3492 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_1511
timestamp 1607319584
transform -1 0 3556 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_257
timestamp 1607319584
transform 1 0 3556 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_208
timestamp 1607319584
transform -1 0 3612 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_6_0
timestamp 1607319584
transform 1 0 3612 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_6_1
timestamp 1607319584
transform 1 0 3620 0 1 1105
box -2 -3 10 103
use BUFX4  BUFX4_301
timestamp 1607319584
transform 1 0 3628 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_294
timestamp 1607319584
transform -1 0 3708 0 1 1105
box -2 -3 50 103
use INVX1  INVX1_265
timestamp 1607319584
transform 1 0 3708 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_354
timestamp 1607319584
transform -1 0 3748 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_926
timestamp 1607319584
transform 1 0 3748 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_87
timestamp 1607319584
transform -1 0 3828 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_100
timestamp 1607319584
transform -1 0 3876 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_925
timestamp 1607319584
transform -1 0 3908 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_186
timestamp 1607319584
transform -1 0 3940 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_457
timestamp 1607319584
transform -1 0 4036 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_768
timestamp 1607319584
transform 1 0 4036 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_279
timestamp 1607319584
transform 1 0 4060 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_178
timestamp 1607319584
transform -1 0 4132 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_7_0
timestamp 1607319584
transform 1 0 4132 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_7_1
timestamp 1607319584
transform 1 0 4140 0 1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_277
timestamp 1607319584
transform 1 0 4148 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_711
timestamp 1607319584
transform -1 0 4228 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_374
timestamp 1607319584
transform -1 0 4244 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_918
timestamp 1607319584
transform -1 0 4340 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_773
timestamp 1607319584
transform -1 0 4364 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_135
timestamp 1607319584
transform 1 0 4364 0 1 1105
box -2 -3 50 103
use AOI21X1  AOI21X1_212
timestamp 1607319584
transform 1 0 4412 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_261
timestamp 1607319584
transform -1 0 4468 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_771
timestamp 1607319584
transform -1 0 4492 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1163
timestamp 1607319584
transform -1 0 4524 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_278
timestamp 1607319584
transform 1 0 4524 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_1164
timestamp 1607319584
transform -1 0 4604 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_187
timestamp 1607319584
transform 1 0 4604 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_8_0
timestamp 1607319584
transform 1 0 4628 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_8_1
timestamp 1607319584
transform 1 0 4636 0 1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_325
timestamp 1607319584
transform 1 0 4644 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_718
timestamp 1607319584
transform -1 0 4724 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_375
timestamp 1607319584
transform -1 0 4740 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_934
timestamp 1607319584
transform -1 0 4836 0 1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_259
timestamp 1607319584
transform 1 0 4836 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_210
timestamp 1607319584
transform -1 0 4892 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_163
timestamp 1607319584
transform -1 0 4924 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_218
timestamp 1607319584
transform 1 0 4924 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_269
timestamp 1607319584
transform 1 0 4956 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_722
timestamp 1607319584
transform 1 0 4980 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_184
timestamp 1607319584
transform -1 0 5028 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_947
timestamp 1607319584
transform -1 0 5124 0 1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_23
timestamp 1607319584
transform 1 0 5124 0 1 1105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_657
timestamp 1607319584
transform 1 0 4 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_418
timestamp 1607319584
transform 1 0 100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_417
timestamp 1607319584
transform -1 0 164 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_316
timestamp 1607319584
transform -1 0 188 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_891
timestamp 1607319584
transform -1 0 220 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_264
timestamp 1607319584
transform 1 0 220 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_671
timestamp 1607319584
transform 1 0 244 0 -1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_219
timestamp 1607319584
transform -1 0 364 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_500
timestamp 1607319584
transform 1 0 364 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_499
timestamp 1607319584
transform 1 0 396 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_317
timestamp 1607319584
transform -1 0 452 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_660
timestamp 1607319584
transform -1 0 476 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1018
timestamp 1607319584
transform 1 0 476 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_0_0
timestamp 1607319584
transform 1 0 572 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1607319584
transform 1 0 580 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_1082
timestamp 1607319584
transform 1 0 588 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_522
timestamp 1607319584
transform -1 0 644 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_188
timestamp 1607319584
transform 1 0 644 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_232
timestamp 1607319584
transform 1 0 676 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_228
timestamp 1607319584
transform 1 0 700 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_818
timestamp 1607319584
transform -1 0 820 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_615
timestamp 1607319584
transform 1 0 820 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_900
timestamp 1607319584
transform 1 0 852 0 -1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_97
timestamp 1607319584
transform -1 0 956 0 -1 1305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_615
timestamp 1607319584
transform 1 0 956 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_1_0
timestamp 1607319584
transform -1 0 1060 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1607319584
transform -1 0 1068 0 -1 1305
box -2 -3 10 103
use BUFX4  BUFX4_308
timestamp 1607319584
transform -1 0 1100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_357
timestamp 1607319584
transform 1 0 1100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_358
timestamp 1607319584
transform -1 0 1164 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_419
timestamp 1607319584
transform 1 0 1164 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_656
timestamp 1607319584
transform -1 0 1204 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1671
timestamp 1607319584
transform 1 0 1204 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_326
timestamp 1607319584
transform 1 0 1236 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_337
timestamp 1607319584
transform -1 0 1348 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_1207
timestamp 1607319584
transform 1 0 1348 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_657
timestamp 1607319584
transform 1 0 1380 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_311
timestamp 1607319584
transform 1 0 1404 0 -1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_221
timestamp 1607319584
transform -1 0 1476 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1006
timestamp 1607319584
transform -1 0 1572 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_2_0
timestamp 1607319584
transform 1 0 1572 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1607319584
transform 1 0 1580 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_225
timestamp 1607319584
transform 1 0 1588 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_183
timestamp 1607319584
transform -1 0 1644 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1272
timestamp 1607319584
transform -1 0 1676 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_56
timestamp 1607319584
transform 1 0 1676 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_70
timestamp 1607319584
transform 1 0 1708 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_592
timestamp 1607319584
transform -1 0 1828 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_629
timestamp 1607319584
transform 1 0 1828 0 -1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_55
timestamp 1607319584
transform 1 0 1924 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_69
timestamp 1607319584
transform 1 0 1956 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_588
timestamp 1607319584
transform 1 0 1980 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_710
timestamp 1607319584
transform -1 0 2028 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1256
timestamp 1607319584
transform -1 0 2060 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_3_0
timestamp 1607319584
transform 1 0 2060 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1607319584
transform 1 0 2068 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_1079
timestamp 1607319584
transform 1 0 2076 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_383
timestamp 1607319584
transform 1 0 2108 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_451
timestamp 1607319584
transform -1 0 2164 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_261
timestamp 1607319584
transform -1 0 2188 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_310
timestamp 1607319584
transform 1 0 2188 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1255
timestamp 1607319584
transform -1 0 2244 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_404
timestamp 1607319584
transform 1 0 2244 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_403
timestamp 1607319584
transform -1 0 2308 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_638
timestamp 1607319584
transform -1 0 2404 0 -1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_61
timestamp 1607319584
transform -1 0 2428 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_298
timestamp 1607319584
transform -1 0 2476 0 -1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_589
timestamp 1607319584
transform -1 0 2572 0 -1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_220
timestamp 1607319584
transform -1 0 2596 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_4_0
timestamp 1607319584
transform -1 0 2604 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_4_1
timestamp 1607319584
transform -1 0 2612 0 -1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_178
timestamp 1607319584
transform -1 0 2644 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_300
timestamp 1607319584
transform 1 0 2644 0 -1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_1001
timestamp 1607319584
transform -1 0 2788 0 -1 1305
box -2 -3 98 103
use BUFX4  BUFX4_219
timestamp 1607319584
transform 1 0 2788 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_219
timestamp 1607319584
transform 1 0 2820 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_260
timestamp 1607319584
transform 1 0 2844 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_225
timestamp 1607319584
transform 1 0 2876 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_255
timestamp 1607319584
transform 1 0 2908 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_838
timestamp 1607319584
transform 1 0 2940 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1553
timestamp 1607319584
transform -1 0 2996 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_233
timestamp 1607319584
transform 1 0 2996 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_5_0
timestamp 1607319584
transform 1 0 3092 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_5_1
timestamp 1607319584
transform 1 0 3100 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_14
timestamp 1607319584
transform 1 0 3108 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_800
timestamp 1607319584
transform 1 0 3124 0 -1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_3
timestamp 1607319584
transform -1 0 3196 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_246
timestamp 1607319584
transform -1 0 3220 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_211
timestamp 1607319584
transform -1 0 3244 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_810
timestamp 1607319584
transform -1 0 3268 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_265
timestamp 1607319584
transform 1 0 3268 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_195
timestamp 1607319584
transform 1 0 3292 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_209
timestamp 1607319584
transform 1 0 3324 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_258
timestamp 1607319584
transform -1 0 3380 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_375
timestamp 1607319584
transform 1 0 3380 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_990
timestamp 1607319584
transform -1 0 3444 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_423
timestamp 1607319584
transform 1 0 3444 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_272
timestamp 1607319584
transform 1 0 3468 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1607319584
transform -1 0 3588 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_849
timestamp 1607319584
transform -1 0 3620 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_6_0
timestamp 1607319584
transform 1 0 3620 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_6_1
timestamp 1607319584
transform 1 0 3628 0 -1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_43
timestamp 1607319584
transform 1 0 3636 0 -1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_491
timestamp 1607319584
transform -1 0 3708 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1053
timestamp 1607319584
transform -1 0 3740 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_196
timestamp 1607319584
transform 1 0 3740 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_801
timestamp 1607319584
transform -1 0 3820 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_248
timestamp 1607319584
transform -1 0 3844 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_102
timestamp 1607319584
transform 1 0 3844 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_185
timestamp 1607319584
transform 1 0 3892 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_146
timestamp 1607319584
transform -1 0 3956 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_147
timestamp 1607319584
transform 1 0 3956 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_461
timestamp 1607319584
transform -1 0 4084 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_1036
timestamp 1607319584
transform 1 0 4084 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_7_0
timestamp 1607319584
transform 1 0 4116 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_7_1
timestamp 1607319584
transform 1 0 4124 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_180
timestamp 1607319584
transform 1 0 4132 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1607319584
transform -1 0 4252 0 -1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_229
timestamp 1607319584
transform 1 0 4252 0 -1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_209
timestamp 1607319584
transform 1 0 4300 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_169
timestamp 1607319584
transform -1 0 4356 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1098
timestamp 1607319584
transform -1 0 4388 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_310
timestamp 1607319584
transform 1 0 4388 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_710
timestamp 1607319584
transform 1 0 4404 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_179
timestamp 1607319584
transform 1 0 4436 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_548
timestamp 1607319584
transform 1 0 4460 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_940
timestamp 1607319584
transform -1 0 4580 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_181
timestamp 1607319584
transform 1 0 4580 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_712
timestamp 1607319584
transform -1 0 4636 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_8_0
timestamp 1607319584
transform 1 0 4636 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_8_1
timestamp 1607319584
transform 1 0 4644 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_438
timestamp 1607319584
transform 1 0 4652 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_1226
timestamp 1607319584
transform 1 0 4668 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_410
timestamp 1607319584
transform 1 0 4700 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_679
timestamp 1607319584
transform 1 0 4724 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_411
timestamp 1607319584
transform 1 0 4748 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_233
timestamp 1607319584
transform 1 0 4772 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1607319584
transform -1 0 4892 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1607319584
transform -1 0 4988 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_191
timestamp 1607319584
transform 1 0 4988 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1170
timestamp 1607319584
transform -1 0 5044 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1311
timestamp 1607319584
transform -1 0 5076 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_382
timestamp 1607319584
transform -1 0 5092 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1607319584
transform 1 0 5092 0 -1 1305
box -2 -3 98 103
use FILL  FILL_13_1
timestamp 1607319584
transform -1 0 5196 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_672
timestamp 1607319584
transform 1 0 4 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_448
timestamp 1607319584
transform -1 0 132 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_447
timestamp 1607319584
transform -1 0 164 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_54
timestamp 1607319584
transform 1 0 164 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_666
timestamp 1607319584
transform 1 0 180 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_436
timestamp 1607319584
transform 1 0 276 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_435
timestamp 1607319584
transform -1 0 340 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_446
timestamp 1607319584
transform 1 0 340 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_445
timestamp 1607319584
transform -1 0 404 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_438
timestamp 1607319584
transform 1 0 404 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_667
timestamp 1607319584
transform 1 0 436 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_0_0
timestamp 1607319584
transform -1 0 540 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1607319584
transform -1 0 548 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_1210
timestamp 1607319584
transform -1 0 580 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_997
timestamp 1607319584
transform -1 0 612 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_209
timestamp 1607319584
transform -1 0 628 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_324
timestamp 1607319584
transform -1 0 724 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_1669
timestamp 1607319584
transform 1 0 724 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_866
timestamp 1607319584
transform -1 0 780 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_112
timestamp 1607319584
transform 1 0 780 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_501
timestamp 1607319584
transform 1 0 796 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_142
timestamp 1607319584
transform 1 0 828 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_729
timestamp 1607319584
transform -1 0 876 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_124
timestamp 1607319584
transform -1 0 908 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1274
timestamp 1607319584
transform -1 0 940 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_154
timestamp 1607319584
transform 1 0 940 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_362
timestamp 1607319584
transform -1 0 1036 0 1 1305
box -2 -3 50 103
use FILL  FILL_13_1_0
timestamp 1607319584
transform 1 0 1036 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1607319584
transform 1 0 1044 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_777
timestamp 1607319584
transform 1 0 1052 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_776
timestamp 1607319584
transform 1 0 1084 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_993
timestamp 1607319584
transform 1 0 1116 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_868
timestamp 1607319584
transform 1 0 1212 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_15
timestamp 1607319584
transform 1 0 1236 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1125
timestamp 1607319584
transform -1 0 1300 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_250
timestamp 1607319584
transform -1 0 1348 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_1206
timestamp 1607319584
transform -1 0 1380 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_377
timestamp 1607319584
transform -1 0 1412 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_408
timestamp 1607319584
transform 1 0 1412 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_640
timestamp 1607319584
transform 1 0 1444 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_727
timestamp 1607319584
transform -1 0 1564 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_2_0
timestamp 1607319584
transform 1 0 1564 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1607319584
transform 1 0 1572 0 1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_252
timestamp 1607319584
transform 1 0 1580 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_388
timestamp 1607319584
transform 1 0 1628 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_359
timestamp 1607319584
transform -1 0 1708 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_387
timestamp 1607319584
transform -1 0 1740 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1607319584
transform 1 0 1740 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_384
timestamp 1607319584
transform 1 0 1764 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_386
timestamp 1607319584
transform 1 0 1796 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_385
timestamp 1607319584
transform 1 0 1828 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_591
timestamp 1607319584
transform 1 0 1860 0 1 1305
box -2 -3 98 103
use INVX1  INVX1_355
timestamp 1607319584
transform -1 0 1972 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_167
timestamp 1607319584
transform -1 0 2020 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_347
timestamp 1607319584
transform -1 0 2068 0 1 1305
box -2 -3 50 103
use FILL  FILL_13_3_0
timestamp 1607319584
transform -1 0 2076 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1607319584
transform -1 0 2084 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_1016
timestamp 1607319584
transform -1 0 2116 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_327
timestamp 1607319584
transform 1 0 2116 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_1672
timestamp 1607319584
transform -1 0 2244 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_401
timestamp 1607319584
transform 1 0 2244 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_1189
timestamp 1607319584
transform 1 0 2260 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_1666
timestamp 1607319584
transform -1 0 2324 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_809
timestamp 1607319584
transform -1 0 2356 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1607319584
transform -1 0 2372 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_321
timestamp 1607319584
transform -1 0 2468 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_517
timestamp 1607319584
transform -1 0 2492 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_67
timestamp 1607319584
transform 1 0 2492 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_53
timestamp 1607319584
transform -1 0 2548 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_25
timestamp 1607319584
transform 1 0 2548 0 1 1305
box -2 -3 50 103
use FILL  FILL_13_4_0
timestamp 1607319584
transform -1 0 2604 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_4_1
timestamp 1607319584
transform -1 0 2612 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_71
timestamp 1607319584
transform -1 0 2636 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_27
timestamp 1607319584
transform 1 0 2636 0 1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_233
timestamp 1607319584
transform 1 0 2684 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_189
timestamp 1607319584
transform -1 0 2740 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1019
timestamp 1607319584
transform -1 0 2836 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_806
timestamp 1607319584
transform 1 0 2836 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_197
timestamp 1607319584
transform 1 0 2868 0 1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1607319584
transform 1 0 2900 0 1 1305
box -2 -3 42 103
use NAND3X1  NAND3X1_2
timestamp 1607319584
transform 1 0 2940 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1607319584
transform 1 0 2972 0 1 1305
box -2 -3 98 103
use INVX1  INVX1_319
timestamp 1607319584
transform -1 0 3084 0 1 1305
box -2 -3 18 103
use FILL  FILL_13_5_0
timestamp 1607319584
transform -1 0 3092 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_5_1
timestamp 1607319584
transform -1 0 3100 0 1 1305
box -2 -3 10 103
use BUFX4  BUFX4_190
timestamp 1607319584
transform -1 0 3132 0 1 1305
box -2 -3 34 103
use OR2X2  OR2X2_1
timestamp 1607319584
transform 1 0 3132 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_320
timestamp 1607319584
transform -1 0 3188 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_212
timestamp 1607319584
transform -1 0 3212 0 1 1305
box -2 -3 26 103
use INVX4  INVX4_2
timestamp 1607319584
transform 1 0 3212 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_298
timestamp 1607319584
transform 1 0 3236 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_774
timestamp 1607319584
transform 1 0 3260 0 1 1305
box -2 -3 26 103
use INVX8  INVX8_4
timestamp 1607319584
transform -1 0 3324 0 1 1305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1607319584
transform 1 0 3324 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_341
timestamp 1607319584
transform 1 0 3420 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_459
timestamp 1607319584
transform 1 0 3444 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_452
timestamp 1607319584
transform -1 0 3636 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_6_0
timestamp 1607319584
transform -1 0 3644 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_6_1
timestamp 1607319584
transform -1 0 3652 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_1298
timestamp 1607319584
transform -1 0 3684 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_61
timestamp 1607319584
transform -1 0 3700 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1607319584
transform -1 0 3796 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_200
timestamp 1607319584
transform -1 0 3828 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_198
timestamp 1607319584
transform 1 0 3828 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_196
timestamp 1607319584
transform -1 0 3908 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_462
timestamp 1607319584
transform -1 0 4004 0 1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_91
timestamp 1607319584
transform -1 0 4052 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_913
timestamp 1607319584
transform -1 0 4084 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_182
timestamp 1607319584
transform -1 0 4132 0 1 1305
box -2 -3 50 103
use FILL  FILL_13_7_0
timestamp 1607319584
transform 1 0 4132 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_7_1
timestamp 1607319584
transform 1 0 4140 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_471
timestamp 1607319584
transform 1 0 4148 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_1035
timestamp 1607319584
transform -1 0 4204 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_125
timestamp 1607319584
transform 1 0 4204 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_1299
timestamp 1607319584
transform 1 0 4220 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_758
timestamp 1607319584
transform -1 0 4276 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_960
timestamp 1607319584
transform -1 0 4372 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_917
timestamp 1607319584
transform -1 0 4468 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_194
timestamp 1607319584
transform 1 0 4468 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_156
timestamp 1607319584
transform -1 0 4524 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_190
timestamp 1607319584
transform 1 0 4524 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_919
timestamp 1607319584
transform 1 0 4548 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_8_0
timestamp 1607319584
transform 1 0 4644 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_8_1
timestamp 1607319584
transform 1 0 4652 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_716
timestamp 1607319584
transform 1 0 4660 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_247
timestamp 1607319584
transform -1 0 4708 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_932
timestamp 1607319584
transform 1 0 4708 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_725
timestamp 1607319584
transform 1 0 4804 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_376
timestamp 1607319584
transform -1 0 4852 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_950
timestamp 1607319584
transform -1 0 4948 0 1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_213
timestamp 1607319584
transform 1 0 4948 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_262
timestamp 1607319584
transform 1 0 4980 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_159
timestamp 1607319584
transform 1 0 5004 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_772
timestamp 1607319584
transform 1 0 5036 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_197
timestamp 1607319584
transform -1 0 5084 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_943
timestamp 1607319584
transform -1 0 5180 0 1 1305
box -2 -3 98 103
use FILL  FILL_14_1
timestamp 1607319584
transform 1 0 5180 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1607319584
transform 1 0 5188 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_658
timestamp 1607319584
transform 1 0 4 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_420
timestamp 1607319584
transform 1 0 100 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_419
timestamp 1607319584
transform -1 0 164 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_184
timestamp 1607319584
transform 1 0 164 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_386
timestamp 1607319584
transform -1 0 220 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_308
timestamp 1607319584
transform -1 0 252 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_842
timestamp 1607319584
transform -1 0 284 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_335
timestamp 1607319584
transform 1 0 284 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_315
timestamp 1607319584
transform -1 0 404 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_104
timestamp 1607319584
transform 1 0 404 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_892
timestamp 1607319584
transform 1 0 420 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_437
timestamp 1607319584
transform 1 0 452 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_659
timestamp 1607319584
transform 1 0 484 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_0_0
timestamp 1607319584
transform 1 0 580 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1607319584
transform 1 0 588 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_422
timestamp 1607319584
transform 1 0 596 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_421
timestamp 1607319584
transform -1 0 660 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_338
timestamp 1607319584
transform -1 0 684 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_110
timestamp 1607319584
transform 1 0 684 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_138
timestamp 1607319584
transform -1 0 740 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_384
timestamp 1607319584
transform -1 0 764 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_476
timestamp 1607319584
transform 1 0 764 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_502
timestamp 1607319584
transform 1 0 788 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_699
timestamp 1607319584
transform 1 0 820 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_386
timestamp 1607319584
transform -1 0 940 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_956
timestamp 1607319584
transform 1 0 940 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_602
timestamp 1607319584
transform 1 0 972 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_1_0
timestamp 1607319584
transform 1 0 1068 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1607319584
transform 1 0 1076 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_331
timestamp 1607319584
transform 1 0 1084 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_332
timestamp 1607319584
transform -1 0 1148 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_311
timestamp 1607319584
transform -1 0 1172 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_886
timestamp 1607319584
transform -1 0 1204 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_419
timestamp 1607319584
transform 1 0 1204 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_638
timestamp 1607319584
transform -1 0 1260 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_284
timestamp 1607319584
transform -1 0 1292 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_608
timestamp 1607319584
transform 1 0 1292 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_344
timestamp 1607319584
transform 1 0 1388 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_725
timestamp 1607319584
transform 1 0 1420 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_343
timestamp 1607319584
transform -1 0 1476 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_613
timestamp 1607319584
transform 1 0 1476 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_407
timestamp 1607319584
transform 1 0 1500 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_283
timestamp 1607319584
transform 1 0 1532 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_2_0
timestamp 1607319584
transform 1 0 1564 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1607319584
transform 1 0 1572 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_630
timestamp 1607319584
transform 1 0 1580 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_724
timestamp 1607319584
transform 1 0 1676 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_70
timestamp 1607319584
transform -1 0 1748 0 -1 1505
box -2 -3 50 103
use BUFX4  BUFX4_87
timestamp 1607319584
transform 1 0 1748 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_885
timestamp 1607319584
transform 1 0 1780 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_583
timestamp 1607319584
transform -1 0 1908 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_292
timestamp 1607319584
transform 1 0 1908 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_655
timestamp 1607319584
transform 1 0 1924 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_1143
timestamp 1607319584
transform 1 0 1948 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_637
timestamp 1607319584
transform -1 0 2076 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_3_0
timestamp 1607319584
transform 1 0 2076 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1607319584
transform 1 0 2084 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_402
timestamp 1607319584
transform 1 0 2092 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_401
timestamp 1607319584
transform -1 0 2156 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_839
timestamp 1607319584
transform -1 0 2188 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_869
timestamp 1607319584
transform 1 0 2188 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_1077
timestamp 1607319584
transform -1 0 2244 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_309
timestamp 1607319584
transform 1 0 2244 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_289
timestamp 1607319584
transform -1 0 2292 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_581
timestamp 1607319584
transform -1 0 2388 0 -1 1505
box -2 -3 98 103
use BUFX4  BUFX4_235
timestamp 1607319584
transform -1 0 2420 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_193
timestamp 1607319584
transform -1 0 2452 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1023
timestamp 1607319584
transform -1 0 2548 0 -1 1505
box -2 -3 98 103
use BUFX4  BUFX4_204
timestamp 1607319584
transform 1 0 2548 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_4_0
timestamp 1607319584
transform -1 0 2588 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_4_1
timestamp 1607319584
transform -1 0 2596 0 -1 1505
box -2 -3 10 103
use BUFX4  BUFX4_268
timestamp 1607319584
transform -1 0 2628 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_259
timestamp 1607319584
transform 1 0 2628 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_246
timestamp 1607319584
transform 1 0 2652 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_261
timestamp 1607319584
transform 1 0 2684 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1607319584
transform 1 0 2716 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_291
timestamp 1607319584
transform 1 0 2812 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1607319584
transform 1 0 2836 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_292
timestamp 1607319584
transform 1 0 2932 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_237
timestamp 1607319584
transform -1 0 2988 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_398
timestamp 1607319584
transform -1 0 3020 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_620
timestamp 1607319584
transform -1 0 3044 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_296
timestamp 1607319584
transform 1 0 3044 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_765
timestamp 1607319584
transform 1 0 3068 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_5_0
timestamp 1607319584
transform 1 0 3092 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_5_1
timestamp 1607319584
transform 1 0 3100 0 -1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_294
timestamp 1607319584
transform 1 0 3108 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_755
timestamp 1607319584
transform 1 0 3132 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_285
timestamp 1607319584
transform 1 0 3156 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_254
timestamp 1607319584
transform 1 0 3180 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_264
timestamp 1607319584
transform -1 0 3228 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_439
timestamp 1607319584
transform 1 0 3228 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_460
timestamp 1607319584
transform -1 0 3348 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_422
timestamp 1607319584
transform 1 0 3348 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_191
timestamp 1607319584
transform -1 0 3404 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_192
timestamp 1607319584
transform -1 0 3436 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_370
timestamp 1607319584
transform 1 0 3436 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_190
timestamp 1607319584
transform 1 0 3460 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_189
timestamp 1607319584
transform -1 0 3524 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_12
timestamp 1607319584
transform -1 0 3548 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_175
timestamp 1607319584
transform -1 0 3580 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_176
timestamp 1607319584
transform -1 0 3612 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_6_0
timestamp 1607319584
transform 1 0 3612 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_6_1
timestamp 1607319584
transform 1 0 3620 0 -1 1505
box -2 -3 10 103
use BUFX4  BUFX4_282
timestamp 1607319584
transform 1 0 3628 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_715
timestamp 1607319584
transform 1 0 3660 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_229
timestamp 1607319584
transform 1 0 3684 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_199
timestamp 1607319584
transform 1 0 3708 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_464
timestamp 1607319584
transform -1 0 3836 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_577
timestamp 1607319584
transform 1 0 3836 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_195
timestamp 1607319584
transform 1 0 3860 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_193
timestamp 1607319584
transform 1 0 3892 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_194
timestamp 1607319584
transform -1 0 3956 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_508
timestamp 1607319584
transform 1 0 3956 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_248
timestamp 1607319584
transform -1 0 3996 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_948
timestamp 1607319584
transform -1 0 4092 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_479
timestamp 1607319584
transform 1 0 4092 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_7_0
timestamp 1607319584
transform 1 0 4116 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_7_1
timestamp 1607319584
transform 1 0 4124 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1607319584
transform 1 0 4132 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_317
timestamp 1607319584
transform 1 0 4228 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_748
timestamp 1607319584
transform 1 0 4244 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_235
timestamp 1607319584
transform -1 0 4316 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_1105
timestamp 1607319584
transform 1 0 4316 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_260
timestamp 1607319584
transform -1 0 4372 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_211
timestamp 1607319584
transform -1 0 4404 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1607319584
transform -1 0 4500 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1301
timestamp 1607319584
transform 1 0 4500 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_760
timestamp 1607319584
transform -1 0 4556 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_957
timestamp 1607319584
transform -1 0 4652 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_8_0
timestamp 1607319584
transform 1 0 4652 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_8_1
timestamp 1607319584
transform 1 0 4660 0 -1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_185
timestamp 1607319584
transform 1 0 4668 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_206
timestamp 1607319584
transform 1 0 4692 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_166
timestamp 1607319584
transform -1 0 4748 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_283
timestamp 1607319584
transform 1 0 4748 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_1169
timestamp 1607319584
transform 1 0 4796 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_194
timestamp 1607319584
transform -1 0 4852 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_617
timestamp 1607319584
transform 1 0 4852 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_15
timestamp 1607319584
transform -1 0 4908 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1227
timestamp 1607319584
transform -1 0 4940 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_678
timestamp 1607319584
transform 1 0 4940 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_477
timestamp 1607319584
transform 1 0 4964 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_719
timestamp 1607319584
transform 1 0 5060 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_935
timestamp 1607319584
transform -1 0 5188 0 -1 1505
box -2 -3 98 103
use FILL  FILL_15_1
timestamp 1607319584
transform -1 0 5196 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1002
timestamp 1607319584
transform 1 0 4 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_179
timestamp 1607319584
transform 1 0 100 0 1 1505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_85
timestamp 1607319584
transform 1 0 4 0 -1 1705
box -2 -3 74 103
use AOI21X1  AOI21X1_181
timestamp 1607319584
transform 1 0 76 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_221
timestamp 1607319584
transform -1 0 156 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1007
timestamp 1607319584
transform 1 0 156 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_223
timestamp 1607319584
transform -1 0 132 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_331
timestamp 1607319584
transform 1 0 132 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_226
timestamp 1607319584
transform 1 0 252 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_779
timestamp 1607319584
transform 1 0 276 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_994
timestamp 1607319584
transform 1 0 228 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_778
timestamp 1607319584
transform -1 0 340 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_102
timestamp 1607319584
transform 1 0 340 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_890
timestamp 1607319584
transform 1 0 356 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_338
timestamp 1607319584
transform -1 0 420 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_123
timestamp 1607319584
transform 1 0 324 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_997
timestamp 1607319584
transform 1 0 340 0 -1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_185
timestamp 1607319584
transform 1 0 420 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_227
timestamp 1607319584
transform -1 0 476 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1008
timestamp 1607319584
transform 1 0 476 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_785
timestamp 1607319584
transform 1 0 436 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_784
timestamp 1607319584
transform -1 0 500 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_315
timestamp 1607319584
transform 1 0 500 0 -1 1705
box -2 -3 18 103
use FILL  FILL_15_0_0
timestamp 1607319584
transform -1 0 580 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1607319584
transform -1 0 588 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_751
timestamp 1607319584
transform -1 0 612 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_507
timestamp 1607319584
transform 1 0 516 0 -1 1705
box -2 -3 18 103
use FILL  FILL_16_0_0
timestamp 1607319584
transform 1 0 532 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1607319584
transform 1 0 540 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_1295
timestamp 1607319584
transform 1 0 548 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_911
timestamp 1607319584
transform 1 0 580 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_337
timestamp 1607319584
transform -1 0 636 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_166
timestamp 1607319584
transform 1 0 636 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_865
timestamp 1607319584
transform -1 0 676 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_827
timestamp 1607319584
transform 1 0 676 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1668
timestamp 1607319584
transform -1 0 644 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_912
timestamp 1607319584
transform 1 0 644 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_89
timestamp 1607319584
transform 1 0 676 0 -1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_1005
timestamp 1607319584
transform -1 0 868 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_954
timestamp 1607319584
transform 1 0 724 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_682
timestamp 1607319584
transform -1 0 780 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_194
timestamp 1607319584
transform 1 0 780 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_182
timestamp 1607319584
transform 1 0 868 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_224
timestamp 1607319584
transform -1 0 924 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_238
timestamp 1607319584
transform -1 0 836 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1024
timestamp 1607319584
transform 1 0 836 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_544
timestamp 1607319584
transform -1 0 948 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_361
timestamp 1607319584
transform -1 0 996 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_864
timestamp 1607319584
transform -1 0 1020 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_1103
timestamp 1607319584
transform 1 0 932 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_752
timestamp 1607319584
transform -1 0 988 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1667
timestamp 1607319584
transform -1 0 1020 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_363
timestamp 1607319584
transform 1 0 1020 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_1_0
timestamp 1607319584
transform 1 0 1068 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1607319584
transform 1 0 1076 0 1 1505
box -2 -3 10 103
use BUFX4  BUFX4_149
timestamp 1607319584
transform 1 0 1084 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_395
timestamp 1607319584
transform -1 0 1044 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_1_0
timestamp 1607319584
transform 1 0 1044 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1607319584
transform 1 0 1052 0 -1 1705
box -2 -3 10 103
use INVX1  INVX1_81
timestamp 1607319584
transform 1 0 1060 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_334
timestamp 1607319584
transform 1 0 1076 0 -1 1705
box -2 -3 98 103
use BUFX4  BUFX4_117
timestamp 1607319584
transform -1 0 1148 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_122
timestamp 1607319584
transform -1 0 1196 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_569
timestamp 1607319584
transform 1 0 1196 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_230
timestamp 1607319584
transform 1 0 1172 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_869
timestamp 1607319584
transform 1 0 1196 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_633
timestamp 1607319584
transform 1 0 1220 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_262
timestamp 1607319584
transform 1 0 1316 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_293
timestamp 1607319584
transform 1 0 1228 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_303
timestamp 1607319584
transform 1 0 1252 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_381
timestamp 1607319584
transform -1 0 1308 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_378
timestamp 1607319584
transform -1 0 1340 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_393
timestamp 1607319584
transform -1 0 1372 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_394
timestamp 1607319584
transform -1 0 1404 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_482
timestamp 1607319584
transform 1 0 1404 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_328
timestamp 1607319584
transform 1 0 1340 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1270
timestamp 1607319584
transform 1 0 1420 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_870
timestamp 1607319584
transform -1 0 1476 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_840
timestamp 1607319584
transform -1 0 1508 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_52
timestamp 1607319584
transform -1 0 1524 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_1673
timestamp 1607319584
transform -1 0 1468 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1253
timestamp 1607319584
transform 1 0 1468 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_346
timestamp 1607319584
transform -1 0 1548 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_358
timestamp 1607319584
transform -1 0 1572 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_2_0
timestamp 1607319584
transform 1 0 1572 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1607319584
transform 1 0 1580 0 1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_360
timestamp 1607319584
transform 1 0 1588 0 1 1505
box -2 -3 50 103
use FILL  FILL_16_2_0
timestamp 1607319584
transform 1 0 1548 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1607319584
transform 1 0 1556 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_580
timestamp 1607319584
transform 1 0 1564 0 -1 1705
box -2 -3 98 103
use BUFX4  BUFX4_385
timestamp 1607319584
transform -1 0 1668 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1269
timestamp 1607319584
transform -1 0 1700 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_72
timestamp 1607319584
transform 1 0 1700 0 1 1505
box -2 -3 50 103
use INVX1  INVX1_225
timestamp 1607319584
transform 1 0 1660 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_72
timestamp 1607319584
transform 1 0 1676 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_308
timestamp 1607319584
transform -1 0 1732 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_312
timestamp 1607319584
transform -1 0 1796 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_310
timestamp 1607319584
transform -1 0 1844 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_1013
timestamp 1607319584
transform 1 0 1732 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_166
timestamp 1607319584
transform 1 0 1764 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_348
timestamp 1607319584
transform 1 0 1812 0 -1 1705
box -2 -3 50 103
use INVX1  INVX1_356
timestamp 1607319584
transform 1 0 1844 0 1 1505
box -2 -3 18 103
use INVX1  INVX1_417
timestamp 1607319584
transform 1 0 1860 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_311
timestamp 1607319584
transform -1 0 1908 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1205
timestamp 1607319584
transform 1 0 1908 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1607319584
transform 1 0 1860 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_236
timestamp 1607319584
transform -1 0 1908 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_192
timestamp 1607319584
transform -1 0 1940 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1080
timestamp 1607319584
transform 1 0 1940 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_520
timestamp 1607319584
transform 1 0 1972 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_214
timestamp 1607319584
transform -1 0 2044 0 1 1505
box -2 -3 50 103
use BUFX4  BUFX4_188
timestamp 1607319584
transform -1 0 1972 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_184
timestamp 1607319584
transform 1 0 1972 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_205
timestamp 1607319584
transform -1 0 2036 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_215
timestamp 1607319584
transform -1 0 2092 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_3_0
timestamp 1607319584
transform -1 0 2100 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1607319584
transform -1 0 2108 0 1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_35
timestamp 1607319584
transform -1 0 2156 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_216
timestamp 1607319584
transform 1 0 2036 0 -1 1705
box -2 -3 50 103
use FILL  FILL_16_3_0
timestamp 1607319584
transform 1 0 2084 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1607319584
transform 1 0 2092 0 -1 1705
box -2 -3 10 103
use BUFX4  BUFX4_306
timestamp 1607319584
transform 1 0 2100 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_36
timestamp 1607319584
transform -1 0 2204 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_34
timestamp 1607319584
transform -1 0 2252 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_863
timestamp 1607319584
transform 1 0 2132 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_589
timestamp 1607319584
transform -1 0 2180 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_222
timestamp 1607319584
transform -1 0 2204 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_180
timestamp 1607319584
transform -1 0 2236 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_73
timestamp 1607319584
transform 1 0 2252 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_837
timestamp 1607319584
transform 1 0 2276 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_272
timestamp 1607319584
transform -1 0 2340 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_49
timestamp 1607319584
transform -1 0 2252 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_577
timestamp 1607319584
transform -1 0 2348 0 -1 1705
box -2 -3 98 103
use BUFX4  BUFX4_29
timestamp 1607319584
transform 1 0 2340 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_218
timestamp 1607319584
transform -1 0 2404 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_237
timestamp 1607319584
transform -1 0 2428 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_305
timestamp 1607319584
transform 1 0 2348 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_683
timestamp 1607319584
transform 1 0 2380 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_407
timestamp 1607319584
transform 1 0 2404 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_271
timestamp 1607319584
transform -1 0 2460 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_182
timestamp 1607319584
transform -1 0 2492 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_468
timestamp 1607319584
transform 1 0 2492 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_444
timestamp 1607319584
transform -1 0 2444 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_545
timestamp 1607319584
transform 1 0 2444 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1015
timestamp 1607319584
transform -1 0 2564 0 -1 1705
box -2 -3 98 103
use FILL  FILL_15_4_0
timestamp 1607319584
transform 1 0 2588 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_4_1
timestamp 1607319584
transform 1 0 2596 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_218
timestamp 1607319584
transform 1 0 2604 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_204
timestamp 1607319584
transform -1 0 2652 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_413
timestamp 1607319584
transform 1 0 2564 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_4_0
timestamp 1607319584
transform 1 0 2596 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_4_1
timestamp 1607319584
transform 1 0 2604 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_26
timestamp 1607319584
transform 1 0 2612 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_234
timestamp 1607319584
transform 1 0 2652 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_212
timestamp 1607319584
transform 1 0 2684 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_24
timestamp 1607319584
transform 1 0 2716 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_470
timestamp 1607319584
transform 1 0 2636 0 -1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_236
timestamp 1607319584
transform 1 0 2748 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1006
timestamp 1607319584
transform 1 0 2780 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_160
timestamp 1607319584
transform -1 0 2860 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_206
timestamp 1607319584
transform -1 0 2764 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_346
timestamp 1607319584
transform 1 0 2764 0 -1 1705
box -2 -3 18 103
use CLKBUF1  CLKBUF1_3
timestamp 1607319584
transform 1 0 2780 0 -1 1705
box -2 -3 74 103
use NAND2X1  NAND2X1_209
timestamp 1607319584
transform -1 0 2884 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_310
timestamp 1607319584
transform -1 0 2908 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_210
timestamp 1607319584
transform -1 0 2932 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_275
timestamp 1607319584
transform -1 0 2956 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_551
timestamp 1607319584
transform -1 0 2876 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1607319584
transform -1 0 2972 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_308
timestamp 1607319584
transform 1 0 2956 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_274
timestamp 1607319584
transform -1 0 3004 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_295
timestamp 1607319584
transform 1 0 3004 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_764
timestamp 1607319584
transform -1 0 3052 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_780
timestamp 1607319584
transform 1 0 2972 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1318
timestamp 1607319584
transform -1 0 3028 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_550
timestamp 1607319584
transform -1 0 3052 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_255
timestamp 1607319584
transform 1 0 3052 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_5_0
timestamp 1607319584
transform -1 0 3084 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_5_1
timestamp 1607319584
transform -1 0 3092 0 1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_150
timestamp 1607319584
transform -1 0 3140 0 1 1505
box -2 -3 50 103
use CLKBUF1  CLKBUF1_56
timestamp 1607319584
transform -1 0 3124 0 -1 1705
box -2 -3 74 103
use FILL  FILL_16_5_0
timestamp 1607319584
transform -1 0 3132 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_5_1
timestamp 1607319584
transform -1 0 3140 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_148
timestamp 1607319584
transform -1 0 3188 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_1005
timestamp 1607319584
transform -1 0 3220 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_463
timestamp 1607319584
transform 1 0 3220 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_245
timestamp 1607319584
transform -1 0 3164 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_440
timestamp 1607319584
transform 1 0 3164 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_476
timestamp 1607319584
transform -1 0 3284 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_989
timestamp 1607319584
transform -1 0 3348 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_1172
timestamp 1607319584
transform -1 0 3316 0 -1 1705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_50
timestamp 1607319584
transform 1 0 3316 0 -1 1705
box -2 -3 74 103
use OAI21X1  OAI21X1_198
timestamp 1607319584
transform 1 0 3348 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_197
timestamp 1607319584
transform -1 0 3412 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_217
timestamp 1607319584
transform -1 0 3428 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_455
timestamp 1607319584
transform -1 0 3524 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_646
timestamp 1607319584
transform -1 0 3412 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_153
timestamp 1607319584
transform 1 0 3412 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_941
timestamp 1607319584
transform 1 0 3428 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_181
timestamp 1607319584
transform -1 0 3556 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_409
timestamp 1607319584
transform -1 0 3476 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_451
timestamp 1607319584
transform -1 0 3572 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_182
timestamp 1607319584
transform -1 0 3588 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_133
timestamp 1607319584
transform -1 0 3620 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_6_0
timestamp 1607319584
transform 1 0 3620 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_6_1
timestamp 1607319584
transform 1 0 3628 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_454
timestamp 1607319584
transform 1 0 3636 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_174
timestamp 1607319584
transform 1 0 3572 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_6_0
timestamp 1607319584
transform -1 0 3612 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_6_1
timestamp 1607319584
transform -1 0 3620 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_173
timestamp 1607319584
transform -1 0 3652 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_180
timestamp 1607319584
transform -1 0 3764 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_132
timestamp 1607319584
transform 1 0 3652 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_817
timestamp 1607319584
transform -1 0 3716 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_32
timestamp 1607319584
transform -1 0 3732 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_179
timestamp 1607319584
transform -1 0 3764 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_345
timestamp 1607319584
transform 1 0 3764 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_1133
timestamp 1607319584
transform 1 0 3780 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_285
timestamp 1607319584
transform -1 0 3860 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_284
timestamp 1607319584
transform -1 0 3812 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_187
timestamp 1607319584
transform 1 0 3812 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_21
timestamp 1607319584
transform 1 0 3860 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_1
timestamp 1607319584
transform 1 0 3884 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_22
timestamp 1607319584
transform -1 0 3924 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_183
timestamp 1607319584
transform -1 0 3972 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_188
timestamp 1607319584
transform -1 0 3876 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_458
timestamp 1607319584
transform 1 0 3876 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_723
timestamp 1607319584
transform -1 0 4004 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_375
timestamp 1607319584
transform -1 0 4052 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_301
timestamp 1607319584
transform -1 0 3996 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_203
timestamp 1607319584
transform 1 0 3996 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1171
timestamp 1607319584
transform -1 0 4060 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1302
timestamp 1607319584
transform -1 0 4084 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_187
timestamp 1607319584
transform -1 0 4132 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_7_0
timestamp 1607319584
transform -1 0 4140 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_7_1
timestamp 1607319584
transform -1 0 4148 0 1 1505
box -2 -3 10 103
use BUFX4  BUFX4_269
timestamp 1607319584
transform -1 0 4092 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_273
timestamp 1607319584
transform -1 0 4124 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_7_0
timestamp 1607319584
transform 1 0 4124 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_7_1
timestamp 1607319584
transform 1 0 4132 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_374
timestamp 1607319584
transform 1 0 4140 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_1041
timestamp 1607319584
transform -1 0 4180 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_450
timestamp 1607319584
transform -1 0 4276 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_1292
timestamp 1607319584
transform -1 0 4220 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_171
timestamp 1607319584
transform 1 0 4220 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_178
timestamp 1607319584
transform 1 0 4276 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_281
timestamp 1607319584
transform 1 0 4308 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_1069
timestamp 1607319584
transform 1 0 4324 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_172
timestamp 1607319584
transform -1 0 4284 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_177
timestamp 1607319584
transform 1 0 4284 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1607319584
transform 1 0 4316 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_208
timestamp 1607319584
transform 1 0 4356 0 1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_453
timestamp 1607319584
transform -1 0 4500 0 1 1505
box -2 -3 98 103
use BUFX4  BUFX4_233
timestamp 1607319584
transform 1 0 4348 0 -1 1705
box -2 -3 34 103
use INVX4  INVX4_1
timestamp 1607319584
transform -1 0 4404 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_327
timestamp 1607319584
transform -1 0 4452 0 -1 1705
box -2 -3 50 103
use INVX1  INVX1_253
timestamp 1607319584
transform -1 0 4516 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1607319584
transform -1 0 4612 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_326
timestamp 1607319584
transform 1 0 4452 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_139
timestamp 1607319584
transform 1 0 4500 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_541
timestamp 1607319584
transform 1 0 4548 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_27
timestamp 1607319584
transform 1 0 4612 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_8_0
timestamp 1607319584
transform -1 0 4644 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_8_1
timestamp 1607319584
transform -1 0 4652 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_1228
timestamp 1607319584
transform -1 0 4604 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_978
timestamp 1607319584
transform -1 0 4636 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_8_0
timestamp 1607319584
transform -1 0 4644 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_8_1
timestamp 1607319584
transform -1 0 4652 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_205
timestamp 1607319584
transform -1 0 4684 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_469
timestamp 1607319584
transform 1 0 4684 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_977
timestamp 1607319584
transform -1 0 4684 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_819
timestamp 1607319584
transform -1 0 4716 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_759
timestamp 1607319584
transform 1 0 4716 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1300
timestamp 1607319584
transform -1 0 4772 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_282
timestamp 1607319584
transform 1 0 4780 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_1070
timestamp 1607319584
transform 1 0 4796 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_769
timestamp 1607319584
transform 1 0 4828 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_189
timestamp 1607319584
transform -1 0 4788 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1607319584
transform -1 0 4884 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_19
timestamp 1607319584
transform -1 0 4876 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_479
timestamp 1607319584
transform -1 0 4972 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_647
timestamp 1607319584
transform 1 0 4884 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_381
timestamp 1607319584
transform -1 0 4924 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_1308
timestamp 1607319584
transform -1 0 4956 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_13
timestamp 1607319584
transform 1 0 4972 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_17
timestamp 1607319584
transform -1 0 5028 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_509
timestamp 1607319584
transform -1 0 5052 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_1319
timestamp 1607319584
transform 1 0 5052 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1607319584
transform -1 0 5052 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_781
timestamp 1607319584
transform 1 0 5052 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_383
timestamp 1607319584
transform -1 0 5100 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1607319584
transform -1 0 5196 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_190
timestamp 1607319584
transform -1 0 5092 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1607319584
transform -1 0 5188 0 -1 1705
box -2 -3 98 103
use FILL  FILL_17_1
timestamp 1607319584
transform -1 0 5196 0 -1 1705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_73
timestamp 1607319584
transform 1 0 4 0 1 1705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_1004
timestamp 1607319584
transform 1 0 76 0 1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_304
timestamp 1607319584
transform -1 0 204 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_382
timestamp 1607319584
transform -1 0 228 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1000
timestamp 1607319584
transform 1 0 228 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_791
timestamp 1607319584
transform 1 0 324 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_790
timestamp 1607319584
transform -1 0 388 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_332
timestamp 1607319584
transform 1 0 388 0 1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_305
timestamp 1607319584
transform 1 0 484 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_383
timestamp 1607319584
transform -1 0 540 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_0_0
timestamp 1607319584
transform -1 0 548 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1607319584
transform -1 0 556 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_431
timestamp 1607319584
transform -1 0 580 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_323
timestamp 1607319584
transform 1 0 580 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_145
timestamp 1607319584
transform -1 0 692 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_362
timestamp 1607319584
transform -1 0 716 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_933
timestamp 1607319584
transform 1 0 716 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_999
timestamp 1607319584
transform 1 0 748 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_443
timestamp 1607319584
transform 1 0 844 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_1231
timestamp 1607319584
transform 1 0 860 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_106
timestamp 1607319584
transform 1 0 892 0 1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_1296
timestamp 1607319584
transform 1 0 940 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_322
timestamp 1607319584
transform 1 0 972 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_1_0
timestamp 1607319584
transform -1 0 1076 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1607319584
transform -1 0 1084 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_964
timestamp 1607319584
transform -1 0 1116 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_438
timestamp 1607319584
transform 1 0 1116 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_377
timestamp 1607319584
transform -1 0 1196 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_58
timestamp 1607319584
transform -1 0 1244 0 1 1705
box -2 -3 50 103
use AOI21X1  AOI21X1_307
timestamp 1607319584
transform 1 0 1244 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_385
timestamp 1607319584
transform 1 0 1276 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_330
timestamp 1607319584
transform -1 0 1396 0 1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_309
timestamp 1607319584
transform 1 0 1396 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_387
timestamp 1607319584
transform -1 0 1452 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_465
timestamp 1607319584
transform 1 0 1452 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_707
timestamp 1607319584
transform 1 0 1468 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_336
timestamp 1607319584
transform -1 0 1588 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_2_0
timestamp 1607319584
transform -1 0 1596 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1607319584
transform -1 0 1604 0 1 1705
box -2 -3 10 103
use INVX1  INVX1_176
timestamp 1607319584
transform -1 0 1620 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_819
timestamp 1607319584
transform -1 0 1716 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_616
timestamp 1607319584
transform 1 0 1716 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1607319584
transform 1 0 1748 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_306
timestamp 1607319584
transform -1 0 1804 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_97
timestamp 1607319584
transform -1 0 1820 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_578
timestamp 1607319584
transform -1 0 1916 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_168
timestamp 1607319584
transform 1 0 1916 0 1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_1022
timestamp 1607319584
transform -1 0 2060 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_3_0
timestamp 1607319584
transform -1 0 2068 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1607319584
transform -1 0 2076 0 1 1705
box -2 -3 10 103
use BUFX4  BUFX4_189
timestamp 1607319584
transform -1 0 2108 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_256
timestamp 1607319584
transform -1 0 2140 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_26
timestamp 1607319584
transform 1 0 2140 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_208
timestamp 1607319584
transform 1 0 2172 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_143
timestamp 1607319584
transform -1 0 2228 0 1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_329
timestamp 1607319584
transform 1 0 2228 0 1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_1003
timestamp 1607319584
transform -1 0 2372 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_69
timestamp 1607319584
transform -1 0 2396 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1232
timestamp 1607319584
transform -1 0 2428 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_233
timestamp 1607319584
transform 1 0 2428 0 1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_1104
timestamp 1607319584
transform -1 0 2508 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_797
timestamp 1607319584
transform 1 0 2508 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_795
timestamp 1607319584
transform 1 0 2540 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_316
timestamp 1607319584
transform -1 0 2588 0 1 1705
box -2 -3 18 103
use FILL  FILL_17_4_0
timestamp 1607319584
transform -1 0 2596 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_4_1
timestamp 1607319584
transform -1 0 2604 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1013
timestamp 1607319584
transform -1 0 2700 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_28
timestamp 1607319584
transform 1 0 2700 0 1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_256
timestamp 1607319584
transform 1 0 2724 0 1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_1134
timestamp 1607319584
transform 1 0 2772 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1607319584
transform 1 0 2804 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_320
timestamp 1607319584
transform 1 0 2900 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_1108
timestamp 1607319584
transform -1 0 2948 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1326
timestamp 1607319584
transform 1 0 2948 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_228
timestamp 1607319584
transform 1 0 2980 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_281
timestamp 1607319584
transform -1 0 3036 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1107
timestamp 1607319584
transform -1 0 3068 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_236
timestamp 1607319584
transform 1 0 3068 0 1 1705
box -2 -3 50 103
use FILL  FILL_17_5_0
timestamp 1607319584
transform 1 0 3116 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_5_1
timestamp 1607319584
transform 1 0 3124 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_284
timestamp 1607319584
transform 1 0 3132 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_509
timestamp 1607319584
transform -1 0 3172 0 1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_237
timestamp 1607319584
transform -1 0 3220 0 1 1705
box -2 -3 50 103
use NOR2X1  NOR2X1_16
timestamp 1607319584
transform 1 0 3220 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1607319584
transform -1 0 3276 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1607319584
transform -1 0 3372 0 1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_214
timestamp 1607319584
transform -1 0 3404 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_263
timestamp 1607319584
transform 1 0 3404 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1197
timestamp 1607319584
transform -1 0 3460 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_304
timestamp 1607319584
transform 1 0 3460 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_761
timestamp 1607319584
transform 1 0 3508 0 1 1705
box -2 -3 26 103
use BUFX4  BUFX4_122
timestamp 1607319584
transform 1 0 3532 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1261
timestamp 1607319584
transform -1 0 3596 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_473
timestamp 1607319584
transform -1 0 3612 0 1 1705
box -2 -3 18 103
use FILL  FILL_17_6_0
timestamp 1607319584
transform 1 0 3612 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_6_1
timestamp 1607319584
transform 1 0 3620 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_757
timestamp 1607319584
transform 1 0 3628 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_456
timestamp 1607319584
transform -1 0 3748 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_184
timestamp 1607319584
transform 1 0 3748 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_183
timestamp 1607319584
transform -1 0 3812 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_134
timestamp 1607319584
transform 1 0 3812 0 1 1705
box -2 -3 34 103
use INVX8  INVX8_8
timestamp 1607319584
transform 1 0 3844 0 1 1705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1607319584
transform 1 0 3884 0 1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_229
timestamp 1607319584
transform 1 0 3980 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_282
timestamp 1607319584
transform 1 0 4012 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_619
timestamp 1607319584
transform -1 0 4060 0 1 1705
box -2 -3 26 103
use BUFX4  BUFX4_275
timestamp 1607319584
transform 1 0 4060 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_7_0
timestamp 1607319584
transform 1 0 4092 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_7_1
timestamp 1607319584
transform 1 0 4100 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_952
timestamp 1607319584
transform 1 0 4108 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_504
timestamp 1607319584
transform 1 0 4204 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_727
timestamp 1607319584
transform -1 0 4252 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_89
timestamp 1607319584
transform 1 0 4252 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_877
timestamp 1607319584
transform 1 0 4268 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_231
timestamp 1607319584
transform 1 0 4300 0 1 1705
box -2 -3 50 103
use BUFX4  BUFX4_251
timestamp 1607319584
transform 1 0 4348 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_395
timestamp 1607319584
transform 1 0 4380 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_169
timestamp 1607319584
transform 1 0 4412 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_170
timestamp 1607319584
transform -1 0 4476 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_449
timestamp 1607319584
transform -1 0 4572 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_777
timestamp 1607319584
transform 1 0 4572 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1315
timestamp 1607319584
transform -1 0 4628 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_8_0
timestamp 1607319584
transform -1 0 4636 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_8_1
timestamp 1607319584
transform -1 0 4644 0 1 1705
box -2 -3 10 103
use INVX1  INVX1_127
timestamp 1607319584
transform -1 0 4660 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1607319584
transform -1 0 4756 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1305
timestamp 1607319584
transform -1 0 4788 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_1303
timestamp 1607319584
transform -1 0 4820 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_34
timestamp 1607319584
transform -1 0 4836 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1607319584
transform 1 0 4836 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_1198
timestamp 1607319584
transform -1 0 4964 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1607319584
transform -1 0 5060 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_29
timestamp 1607319584
transform 1 0 5060 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_207
timestamp 1607319584
transform -1 0 5116 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_256
timestamp 1607319584
transform 1 0 5116 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_207
timestamp 1607319584
transform -1 0 5172 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_34
timestamp 1607319584
transform 1 0 5172 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_984
timestamp 1607319584
transform -1 0 100 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_775
timestamp 1607319584
transform -1 0 132 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_774
timestamp 1607319584
transform -1 0 164 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_506
timestamp 1607319584
transform 1 0 164 0 -1 1905
box -2 -3 18 103
use BUFX4  BUFX4_443
timestamp 1607319584
transform -1 0 212 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_782
timestamp 1607319584
transform 1 0 212 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_783
timestamp 1607319584
transform -1 0 276 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_992
timestamp 1607319584
transform 1 0 276 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_251
timestamp 1607319584
transform 1 0 372 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_1294
timestamp 1607319584
transform 1 0 388 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_750
timestamp 1607319584
transform -1 0 444 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_475
timestamp 1607319584
transform -1 0 468 0 -1 1905
box -2 -3 26 103
use BUFX4  BUFX4_442
timestamp 1607319584
transform 1 0 468 0 -1 1905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_59
timestamp 1607319584
transform 1 0 500 0 -1 1905
box -2 -3 74 103
use FILL  FILL_18_0_0
timestamp 1607319584
transform -1 0 580 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1607319584
transform -1 0 588 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_124
timestamp 1607319584
transform -1 0 604 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_1010
timestamp 1607319584
transform -1 0 700 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_792
timestamp 1607319584
transform 1 0 700 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_252
timestamp 1607319584
transform 1 0 732 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_789
timestamp 1607319584
transform 1 0 748 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1040
timestamp 1607319584
transform -1 0 812 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_788
timestamp 1607319584
transform -1 0 844 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1016
timestamp 1607319584
transform 1 0 844 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_508
timestamp 1607319584
transform 1 0 940 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_798
timestamp 1607319584
transform 1 0 956 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1273
timestamp 1607319584
transform -1 0 1020 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_780
timestamp 1607319584
transform 1 0 1020 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_1_0
timestamp 1607319584
transform -1 0 1060 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1607319584
transform -1 0 1068 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_781
timestamp 1607319584
transform -1 0 1100 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_995
timestamp 1607319584
transform 1 0 1100 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_787
timestamp 1607319584
transform 1 0 1196 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_786
timestamp 1607319584
transform 1 0 1228 0 -1 1905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_83
timestamp 1607319584
transform 1 0 1260 0 -1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_998
timestamp 1607319584
transform 1 0 1332 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_187
timestamp 1607319584
transform 1 0 1428 0 -1 1905
box -2 -3 18 103
use INVX1  INVX1_379
timestamp 1607319584
transform 1 0 1444 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_1167
timestamp 1607319584
transform 1 0 1460 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1141
timestamp 1607319584
transform 1 0 1492 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_262
timestamp 1607319584
transform 1 0 1524 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_2_0
timestamp 1607319584
transform -1 0 1580 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1607319584
transform -1 0 1588 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_353
timestamp 1607319584
transform -1 0 1604 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_584
timestamp 1607319584
transform 1 0 1604 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_481
timestamp 1607319584
transform 1 0 1700 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_312
timestamp 1607319584
transform 1 0 1716 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_76
timestamp 1607319584
transform -1 0 1772 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_156
timestamp 1607319584
transform 1 0 1772 0 -1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_614
timestamp 1607319584
transform 1 0 1820 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_1144
timestamp 1607319584
transform 1 0 1844 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_263
timestamp 1607319584
transform -1 0 1924 0 -1 1905
box -2 -3 50 103
use BUFX4  BUFX4_198
timestamp 1607319584
transform -1 0 1956 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_366
timestamp 1607319584
transform 1 0 1956 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_183
timestamp 1607319584
transform -1 0 2020 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_211
timestamp 1607319584
transform -1 0 2052 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_210
timestamp 1607319584
transform -1 0 2084 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_3_0
timestamp 1607319584
transform 1 0 2084 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1607319584
transform 1 0 2092 0 -1 1905
box -2 -3 10 103
use BUFX4  BUFX4_247
timestamp 1607319584
transform 1 0 2100 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_60
timestamp 1607319584
transform 1 0 2132 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_975
timestamp 1607319584
transform 1 0 2180 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_406
timestamp 1607319584
transform -1 0 2236 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1011
timestamp 1607319584
transform 1 0 2236 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_188
timestamp 1607319584
transform 1 0 2332 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_793
timestamp 1607319584
transform 1 0 2348 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_203
timestamp 1607319584
transform -1 0 2404 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_976
timestamp 1607319584
transform 1 0 2404 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1607319584
transform 1 0 2436 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_208
timestamp 1607319584
transform -1 0 2492 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_474
timestamp 1607319584
transform -1 0 2508 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_472
timestamp 1607319584
transform -1 0 2604 0 -1 1905
box -2 -3 98 103
use FILL  FILL_18_4_0
timestamp 1607319584
transform 1 0 2604 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_4_1
timestamp 1607319584
transform 1 0 2612 0 -1 1905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_40
timestamp 1607319584
transform 1 0 2620 0 -1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_478
timestamp 1607319584
transform 1 0 2692 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_578
timestamp 1607319584
transform -1 0 2812 0 -1 1905
box -2 -3 26 103
use INVX8  INVX8_11
timestamp 1607319584
transform 1 0 2812 0 -1 1905
box -2 -3 42 103
use AOI21X1  AOI21X1_230
timestamp 1607319584
transform 1 0 2852 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_283
timestamp 1607319584
transform -1 0 2908 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1607319584
transform -1 0 3004 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_445
timestamp 1607319584
transform 1 0 3004 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_688
timestamp 1607319584
transform 1 0 3020 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_7
timestamp 1607319584
transform -1 0 3076 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_763
timestamp 1607319584
transform 1 0 3076 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_5_0
timestamp 1607319584
transform -1 0 3108 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_5_1
timestamp 1607319584
transform -1 0 3116 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_1304
timestamp 1607319584
transform -1 0 3148 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1233
timestamp 1607319584
transform 1 0 3148 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_686
timestamp 1607319584
transform 1 0 3180 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1607319584
transform 1 0 3204 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_384
timestamp 1607319584
transform 1 0 3300 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_1327
timestamp 1607319584
transform 1 0 3316 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_475
timestamp 1607319584
transform 1 0 3348 0 -1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1607319584
transform 1 0 3444 0 -1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_287
timestamp 1607319584
transform 1 0 3540 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_232
timestamp 1607319584
transform -1 0 3596 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_275
timestamp 1607319584
transform -1 0 3620 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_6_0
timestamp 1607319584
transform 1 0 3620 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_6_1
timestamp 1607319584
transform 1 0 3628 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_1314
timestamp 1607319584
transform 1 0 3636 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_63
timestamp 1607319584
transform -1 0 3684 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1607319584
transform -1 0 3780 0 -1 1905
box -2 -3 98 103
use BUFX4  BUFX4_194
timestamp 1607319584
transform -1 0 3812 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_285
timestamp 1607319584
transform 1 0 3812 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_785
timestamp 1607319584
transform 1 0 3844 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_489
timestamp 1607319584
transform -1 0 3964 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_192
timestamp 1607319584
transform -1 0 3988 0 -1 1905
box -2 -3 26 103
use BUFX4  BUFX4_201
timestamp 1607319584
transform -1 0 4020 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_241
timestamp 1607319584
transform 1 0 4020 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_239
timestamp 1607319584
transform -1 0 4084 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_196
timestamp 1607319584
transform 1 0 4084 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_343
timestamp 1607319584
transform 1 0 4108 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_7_0
timestamp 1607319584
transform -1 0 4140 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_7_1
timestamp 1607319584
transform -1 0 4148 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_915
timestamp 1607319584
transform -1 0 4180 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_199
timestamp 1607319584
transform -1 0 4212 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1607319584
transform -1 0 4308 0 -1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_278
timestamp 1607319584
transform 1 0 4308 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1607319584
transform 1 0 4332 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_1297
timestamp 1607319584
transform 1 0 4428 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_756
timestamp 1607319584
transform -1 0 4484 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_230
timestamp 1607319584
transform 1 0 4484 0 -1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_234
timestamp 1607319584
transform 1 0 4532 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_1100
timestamp 1607319584
transform -1 0 4588 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_766
timestamp 1607319584
transform 1 0 4588 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_440
timestamp 1607319584
transform -1 0 4628 0 -1 1905
box -2 -3 18 103
use FILL  FILL_18_8_0
timestamp 1607319584
transform -1 0 4636 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_8_1
timestamp 1607319584
transform -1 0 4644 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_951
timestamp 1607319584
transform -1 0 4740 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_726
timestamp 1607319584
transform 1 0 4740 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_762
timestamp 1607319584
transform 1 0 4772 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_13
timestamp 1607319584
transform 1 0 4796 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_9
timestamp 1607319584
transform -1 0 4852 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_473
timestamp 1607319584
transform -1 0 4948 0 -1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_10
timestamp 1607319584
transform 1 0 4948 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1607319584
transform 1 0 4980 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_35
timestamp 1607319584
transform 1 0 5076 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1607319584
transform 1 0 5092 0 -1 1905
box -2 -3 98 103
use FILL  FILL_19_1
timestamp 1607319584
transform -1 0 5196 0 -1 1905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_65
timestamp 1607319584
transform 1 0 4 0 1 1905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_67
timestamp 1607319584
transform 1 0 76 0 1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_979
timestamp 1607319584
transform 1 0 148 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_765
timestamp 1607319584
transform 1 0 244 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_764
timestamp 1607319584
transform -1 0 308 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_996
timestamp 1607319584
transform 1 0 308 0 1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_218
timestamp 1607319584
transform 1 0 404 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_177
timestamp 1607319584
transform -1 0 460 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1039
timestamp 1607319584
transform 1 0 460 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_0_0
timestamp 1607319584
transform 1 0 492 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1607319584
transform 1 0 500 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_971
timestamp 1607319584
transform 1 0 508 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_749
timestamp 1607319584
transform 1 0 604 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_748
timestamp 1607319584
transform -1 0 668 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1012
timestamp 1607319584
transform 1 0 668 0 1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_202
timestamp 1607319584
transform -1 0 788 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_794
timestamp 1607319584
transform 1 0 788 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_204
timestamp 1607319584
transform -1 0 844 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_185
timestamp 1607319584
transform -1 0 892 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_376
timestamp 1607319584
transform 1 0 892 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_201
timestamp 1607319584
transform 1 0 940 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_208
timestamp 1607319584
transform -1 0 988 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_313
timestamp 1607319584
transform 1 0 988 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_728
timestamp 1607319584
transform -1 0 1060 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_1_0
timestamp 1607319584
transform -1 0 1068 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1607319584
transform -1 0 1076 0 1 1905
box -2 -3 10 103
use BUFX4  BUFX4_400
timestamp 1607319584
transform -1 0 1108 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_315
timestamp 1607319584
transform 1 0 1108 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_378
timestamp 1607319584
transform 1 0 1156 0 1 1905
box -2 -3 50 103
use INVX1  INVX1_186
timestamp 1607319584
transform 1 0 1204 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_974
timestamp 1607319584
transform 1 0 1220 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_136
timestamp 1607319584
transform -1 0 1300 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_973
timestamp 1607319584
transform 1 0 1300 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_404
timestamp 1607319584
transform -1 0 1356 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_108
timestamp 1607319584
transform 1 0 1356 0 1 1905
box -2 -3 50 103
use INVX1  INVX1_485
timestamp 1607319584
transform -1 0 1420 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_416
timestamp 1607319584
transform 1 0 1420 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_91
timestamp 1607319584
transform -1 0 1476 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_281
timestamp 1607319584
transform -1 0 1508 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_648
timestamp 1607319584
transform -1 0 1604 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_2_0
timestamp 1607319584
transform -1 0 1612 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1607319584
transform -1 0 1620 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_582
timestamp 1607319584
transform -1 0 1716 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_310
timestamp 1607319584
transform 1 0 1716 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_74
timestamp 1607319584
transform -1 0 1772 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_281
timestamp 1607319584
transform 1 0 1772 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_1168
timestamp 1607319584
transform -1 0 1852 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_206
timestamp 1607319584
transform 1 0 1852 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_796
timestamp 1607319584
transform -1 0 1908 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_380
timestamp 1607319584
transform -1 0 1924 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_1014
timestamp 1607319584
transform 1 0 1924 0 1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_264
timestamp 1607319584
transform 1 0 2020 0 1 1905
box -2 -3 50 103
use FILL  FILL_19_3_0
timestamp 1607319584
transform 1 0 2068 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1607319584
transform 1 0 2076 0 1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_330
timestamp 1607319584
transform 1 0 2084 0 1 1905
box -2 -3 50 103
use BUFX4  BUFX4_264
timestamp 1607319584
transform -1 0 2164 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_35
timestamp 1607319584
transform -1 0 2196 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_33
timestamp 1607319584
transform 1 0 2196 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_265
timestamp 1607319584
transform 1 0 2228 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_217
timestamp 1607319584
transform -1 0 2292 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_830
timestamp 1607319584
transform -1 0 2388 0 1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_141
timestamp 1607319584
transform 1 0 2388 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_113
timestamp 1607319584
transform -1 0 2444 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_137
timestamp 1607319584
transform -1 0 2492 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_138
timestamp 1607319584
transform 1 0 2492 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_207
timestamp 1607319584
transform -1 0 2564 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_205
timestamp 1607319584
transform -1 0 2588 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_4_0
timestamp 1607319584
transform -1 0 2596 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_4_1
timestamp 1607319584
transform -1 0 2604 0 1 1905
box -2 -3 10 103
use BUFX4  BUFX4_34
timestamp 1607319584
transform -1 0 2636 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1262
timestamp 1607319584
transform 1 0 2636 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_352
timestamp 1607319584
transform -1 0 2716 0 1 1905
box -2 -3 50 103
use BUFX4  BUFX4_32
timestamp 1607319584
transform 1 0 2716 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_716
timestamp 1607319584
transform 1 0 2748 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_480
timestamp 1607319584
transform -1 0 2868 0 1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_20
timestamp 1607319584
transform 1 0 2868 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1607319584
transform -1 0 2924 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1607319584
transform 1 0 2924 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_14
timestamp 1607319584
transform -1 0 2980 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_788
timestamp 1607319584
transform -1 0 3004 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1607319584
transform 1 0 3004 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_5_0
timestamp 1607319584
transform -1 0 3108 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_5_1
timestamp 1607319584
transform -1 0 3116 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_1235
timestamp 1607319584
transform -1 0 3148 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1607319584
transform -1 0 3180 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_43
timestamp 1607319584
transform 1 0 3180 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_213
timestamp 1607319584
transform 1 0 3212 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_447
timestamp 1607319584
transform -1 0 3252 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1607319584
transform -1 0 3348 0 1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_789
timestamp 1607319584
transform -1 0 3372 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_1320
timestamp 1607319584
transform 1 0 3372 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_782
timestamp 1607319584
transform -1 0 3428 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_333
timestamp 1607319584
transform -1 0 3476 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_331
timestamp 1607319584
transform 1 0 3476 0 1 1905
box -2 -3 50 103
use AOI21X1  AOI21X1_11
timestamp 1607319584
transform 1 0 3524 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_15
timestamp 1607319584
transform 1 0 3556 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_852
timestamp 1607319584
transform 1 0 3580 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_6_0
timestamp 1607319584
transform 1 0 3612 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_6_1
timestamp 1607319584
transform 1 0 3620 0 1 1905
box -2 -3 10 103
use BUFX4  BUFX4_376
timestamp 1607319584
transform 1 0 3628 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_45
timestamp 1607319584
transform 1 0 3660 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_44
timestamp 1607319584
transform -1 0 3756 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_851
timestamp 1607319584
transform 1 0 3756 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_244
timestamp 1607319584
transform 1 0 3788 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_274
timestamp 1607319584
transform -1 0 3836 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_776
timestamp 1607319584
transform -1 0 3860 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_423
timestamp 1607319584
transform 1 0 3860 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_1323
timestamp 1607319584
transform -1 0 3924 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1607319584
transform 1 0 3924 0 1 1905
box -2 -3 98 103
use INVX1  INVX1_128
timestamp 1607319584
transform 1 0 4020 0 1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_17
timestamp 1607319584
transform 1 0 4036 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_23
timestamp 1607319584
transform 1 0 4068 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_93
timestamp 1607319584
transform 1 0 4092 0 1 1905
box -2 -3 50 103
use FILL  FILL_19_7_0
timestamp 1607319584
transform 1 0 4140 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_7_1
timestamp 1607319584
transform 1 0 4148 0 1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_92
timestamp 1607319584
transform 1 0 4156 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_916
timestamp 1607319584
transform 1 0 4204 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_344
timestamp 1607319584
transform -1 0 4260 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1607319584
transform 1 0 4260 0 1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_225
timestamp 1607319584
transform -1 0 4388 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_201
timestamp 1607319584
transform -1 0 4420 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_33
timestamp 1607319584
transform 1 0 4420 0 1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_232
timestamp 1607319584
transform 1 0 4436 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_818
timestamp 1607319584
transform 1 0 4460 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_231
timestamp 1607319584
transform -1 0 4516 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_255
timestamp 1607319584
transform -1 0 4532 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1607319584
transform -1 0 4628 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_8_0
timestamp 1607319584
transform 1 0 4628 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_8_1
timestamp 1607319584
transform 1 0 4636 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_1317
timestamp 1607319584
transform 1 0 4644 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_779
timestamp 1607319584
transform -1 0 4700 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_64
timestamp 1607319584
transform 1 0 4700 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_195
timestamp 1607319584
transform 1 0 4748 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_878
timestamp 1607319584
transform 1 0 4772 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_302
timestamp 1607319584
transform 1 0 4804 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_193
timestamp 1607319584
transform 1 0 4828 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_724
timestamp 1607319584
transform -1 0 4884 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_312
timestamp 1607319584
transform -1 0 4900 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_949
timestamp 1607319584
transform -1 0 4996 0 1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_14
timestamp 1607319584
transform -1 0 5020 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_474
timestamp 1607319584
transform -1 0 5116 0 1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_223
timestamp 1607319584
transform 1 0 5116 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_276
timestamp 1607319584
transform -1 0 5172 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_235
timestamp 1607319584
transform 1 0 5172 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_965
timestamp 1607319584
transform -1 0 100 0 -1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_174
timestamp 1607319584
transform 1 0 100 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_215
timestamp 1607319584
transform -1 0 156 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_737
timestamp 1607319584
transform -1 0 188 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_736
timestamp 1607319584
transform -1 0 220 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_313
timestamp 1607319584
transform 1 0 220 0 -1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_981
timestamp 1607319584
transform 1 0 236 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_976
timestamp 1607319584
transform 1 0 332 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_769
timestamp 1607319584
transform 1 0 428 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_768
timestamp 1607319584
transform 1 0 460 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_759
timestamp 1607319584
transform 1 0 492 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_314
timestamp 1607319584
transform 1 0 524 0 -1 2105
box -2 -3 18 103
use FILL  FILL_20_0_0
timestamp 1607319584
transform 1 0 540 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1607319584
transform 1 0 548 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_1102
timestamp 1607319584
transform 1 0 556 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_973
timestamp 1607319584
transform 1 0 588 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_753
timestamp 1607319584
transform 1 0 684 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_752
timestamp 1607319584
transform -1 0 748 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_542
timestamp 1607319584
transform -1 0 772 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_1101
timestamp 1607319584
transform 1 0 772 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_200
timestamp 1607319584
transform -1 0 828 0 -1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_186
timestamp 1607319584
transform 1 0 828 0 -1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_970
timestamp 1607319584
transform 1 0 876 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_747
timestamp 1607319584
transform 1 0 972 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_746
timestamp 1607319584
transform -1 0 1036 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_335
timestamp 1607319584
transform -1 0 1060 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_1_0
timestamp 1607319584
transform -1 0 1068 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1607319584
transform -1 0 1076 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_909
timestamp 1607319584
transform -1 0 1108 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_88
timestamp 1607319584
transform 1 0 1108 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_90
timestamp 1607319584
transform 1 0 1156 0 -1 2105
box -2 -3 50 103
use BUFX4  BUFX4_441
timestamp 1607319584
transform 1 0 1204 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_754
timestamp 1607319584
transform 1 0 1236 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_185
timestamp 1607319584
transform 1 0 1268 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_755
timestamp 1607319584
transform -1 0 1316 0 -1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_76
timestamp 1607319584
transform 1 0 1316 0 -1 2105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_974
timestamp 1607319584
transform 1 0 1356 0 -1 2105
box -2 -3 98 103
use INVX8  INVX8_6
timestamp 1607319584
transform -1 0 1492 0 -1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_18
timestamp 1607319584
transform -1 0 1532 0 -1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_611
timestamp 1607319584
transform -1 0 1556 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_2_0
timestamp 1607319584
transform -1 0 1564 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1607319584
transform -1 0 1572 0 -1 2105
box -2 -3 10 103
use AOI22X1  AOI22X1_58
timestamp 1607319584
transform -1 0 1612 0 -1 2105
box -2 -3 42 103
use MUX2X1  MUX2X1_282
timestamp 1607319584
transform 1 0 1612 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_753
timestamp 1607319584
transform 1 0 1660 0 -1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_79
timestamp 1607319584
transform -1 0 1724 0 -1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_736
timestamp 1607319584
transform -1 0 1748 0 -1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_78
timestamp 1607319584
transform -1 0 1788 0 -1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_38
timestamp 1607319584
transform -1 0 1828 0 -1 2105
box -2 -3 42 103
use MUX2X1  MUX2X1_232
timestamp 1607319584
transform -1 0 1876 0 -1 2105
box -2 -3 50 103
use BUFX4  BUFX4_266
timestamp 1607319584
transform -1 0 1908 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_220
timestamp 1607319584
transform 1 0 1908 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_195
timestamp 1607319584
transform -1 0 1972 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_257
timestamp 1607319584
transform 1 0 1972 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_237
timestamp 1607319584
transform -1 0 2036 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_229
timestamp 1607319584
transform 1 0 2036 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_3_0
timestamp 1607319584
transform -1 0 2076 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1607319584
transform -1 0 2084 0 -1 2105
box -2 -3 10 103
use AOI22X1  AOI22X1_68
timestamp 1607319584
transform -1 0 2124 0 -1 2105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_814
timestamp 1607319584
transform 1 0 2124 0 -1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_104
timestamp 1607319584
transform -1 0 2252 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_38
timestamp 1607319584
transform -1 0 2284 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_39
timestamp 1607319584
transform -1 0 2316 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_602
timestamp 1607319584
transform 1 0 2316 0 -1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_28
timestamp 1607319584
transform 1 0 2340 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_234
timestamp 1607319584
transform 1 0 2388 0 -1 2105
box -2 -3 50 103
use INVX1  INVX1_11
timestamp 1607319584
transform 1 0 2436 0 -1 2105
box -2 -3 18 103
use OAI22X1  OAI22X1_2
timestamp 1607319584
transform -1 0 2492 0 -1 2105
box -2 -3 42 103
use INVX1  INVX1_10
timestamp 1607319584
transform -1 0 2508 0 -1 2105
box -2 -3 18 103
use AOI22X1  AOI22X1_28
timestamp 1607319584
transform -1 0 2548 0 -1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_48
timestamp 1607319584
transform -1 0 2588 0 -1 2105
box -2 -3 42 103
use FILL  FILL_20_4_0
timestamp 1607319584
transform 1 0 2588 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_4_1
timestamp 1607319584
transform 1 0 2596 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1607319584
transform 1 0 2604 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_448
timestamp 1607319584
transform 1 0 2700 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_790
timestamp 1607319584
transform 1 0 2716 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_1328
timestamp 1607319584
transform -1 0 2772 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_173
timestamp 1607319584
transform -1 0 2796 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_786
timestamp 1607319584
transform 1 0 2796 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_1236
timestamp 1607319584
transform 1 0 2820 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_1324
timestamp 1607319584
transform -1 0 2884 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1607319584
transform 1 0 2884 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_192
timestamp 1607319584
transform 1 0 2980 0 -1 2105
box -2 -3 18 103
use BUFX4  BUFX4_13
timestamp 1607319584
transform 1 0 2996 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_332
timestamp 1607319584
transform -1 0 3076 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_784
timestamp 1607319584
transform 1 0 3076 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_5_0
timestamp 1607319584
transform -1 0 3108 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_5_1
timestamp 1607319584
transform -1 0 3116 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_1322
timestamp 1607319584
transform -1 0 3148 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1607319584
transform 1 0 3148 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_64
timestamp 1607319584
transform 1 0 3244 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_251
timestamp 1607319584
transform 1 0 3260 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_505
timestamp 1607319584
transform -1 0 3380 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_33
timestamp 1607319584
transform 1 0 3380 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1607319584
transform -1 0 3436 0 -1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_5
timestamp 1607319584
transform -1 0 3476 0 -1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_371
timestamp 1607319584
transform 1 0 3476 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_467
timestamp 1607319584
transform -1 0 3596 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_6_0
timestamp 1607319584
transform 1 0 3596 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_6_1
timestamp 1607319584
transform 1 0 3604 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_487
timestamp 1607319584
transform 1 0 3612 0 -1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_648
timestamp 1607319584
transform 1 0 3708 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1607319584
transform 1 0 3732 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_277
timestamp 1607319584
transform 1 0 3828 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_224
timestamp 1607319584
transform -1 0 3884 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_226
timestamp 1607319584
transform -1 0 3908 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_29
timestamp 1607319584
transform 1 0 3908 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1607319584
transform -1 0 3964 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_495
timestamp 1607319584
transform -1 0 4060 0 -1 2105
box -2 -3 98 103
use INVX2  INVX2_6
timestamp 1607319584
transform 1 0 4060 0 -1 2105
box -2 -3 18 103
use AOI21X1  AOI21X1_233
timestamp 1607319584
transform 1 0 4076 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_288
timestamp 1607319584
transform -1 0 4132 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_7_0
timestamp 1607319584
transform 1 0 4132 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_7_1
timestamp 1607319584
transform 1 0 4140 0 -1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_787
timestamp 1607319584
transform 1 0 4148 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1607319584
transform -1 0 4268 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_465
timestamp 1607319584
transform 1 0 4268 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_31
timestamp 1607319584
transform 1 0 4364 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_201
timestamp 1607319584
transform 1 0 4380 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1607319584
transform -1 0 4436 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_816
timestamp 1607319584
transform 1 0 4436 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_228
timestamp 1607319584
transform 1 0 4468 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_1043
timestamp 1607319584
transform 1 0 4492 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_481
timestamp 1607319584
transform 1 0 4524 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_280
timestamp 1607319584
transform 1 0 4548 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_227
timestamp 1607319584
transform -1 0 4604 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_236
timestamp 1607319584
transform 1 0 4604 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_8_0
timestamp 1607319584
transform -1 0 4636 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_8_1
timestamp 1607319584
transform -1 0 4644 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_202
timestamp 1607319584
transform -1 0 4676 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_466
timestamp 1607319584
transform 1 0 4676 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_90
timestamp 1607319584
transform 1 0 4772 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_620
timestamp 1607319584
transform -1 0 4820 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_432
timestamp 1607319584
transform -1 0 4836 0 -1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_823
timestamp 1607319584
transform -1 0 4932 0 -1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_778
timestamp 1607319584
transform 1 0 4932 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_24
timestamp 1607319584
transform 1 0 4956 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_18
timestamp 1607319584
transform -1 0 5012 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_618
timestamp 1607319584
transform 1 0 5012 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_226
timestamp 1607319584
transform 1 0 5036 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_279
timestamp 1607319584
transform -1 0 5092 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_412
timestamp 1607319584
transform 1 0 5092 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_979
timestamp 1607319584
transform -1 0 5148 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_1316
timestamp 1607319584
transform -1 0 5180 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_191
timestamp 1607319584
transform -1 0 5196 0 -1 2105
box -2 -3 18 103
use BUFX2  BUFX2_8
timestamp 1607319584
transform -1 0 28 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1032
timestamp 1607319584
transform -1 0 124 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_978
timestamp 1607319584
transform 1 0 124 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_763
timestamp 1607319584
transform 1 0 220 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_762
timestamp 1607319584
transform -1 0 284 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_989
timestamp 1607319584
transform 1 0 284 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_972
timestamp 1607319584
transform 1 0 380 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_751
timestamp 1607319584
transform 1 0 476 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_750
timestamp 1607319584
transform -1 0 540 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_0_0
timestamp 1607319584
transform 1 0 540 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1607319584
transform 1 0 548 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_758
timestamp 1607319584
transform 1 0 556 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_543
timestamp 1607319584
transform -1 0 612 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_473
timestamp 1607319584
transform -1 0 636 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_71
timestamp 1607319584
transform -1 0 660 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_74
timestamp 1607319584
transform -1 0 708 0 1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_967
timestamp 1607319584
transform 1 0 708 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_741
timestamp 1607319584
transform 1 0 804 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_740
timestamp 1607319584
transform -1 0 868 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_199
timestamp 1607319584
transform 1 0 868 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_122
timestamp 1607319584
transform 1 0 892 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_198
timestamp 1607319584
transform 1 0 908 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_730
timestamp 1607319584
transform 1 0 932 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_731
timestamp 1607319584
transform -1 0 996 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_962
timestamp 1607319584
transform 1 0 996 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_1_0
timestamp 1607319584
transform -1 0 1100 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1607319584
transform -1 0 1108 0 1 2105
box -2 -3 10 103
use INVX1  INVX1_121
timestamp 1607319584
transform -1 0 1124 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_910
timestamp 1607319584
transform 1 0 1124 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_963
timestamp 1607319584
transform 1 0 1156 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_405
timestamp 1607319584
transform -1 0 1276 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_267
timestamp 1607319584
transform 1 0 1276 0 1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_171
timestamp 1607319584
transform -1 0 1372 0 1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_169
timestamp 1607319584
transform -1 0 1420 0 1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_452
timestamp 1607319584
transform -1 0 1444 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_1017
timestamp 1607319584
transform -1 0 1476 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_229
timestamp 1607319584
transform -1 0 1492 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_412
timestamp 1607319584
transform 1 0 1492 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_87
timestamp 1607319584
transform -1 0 1548 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_2_0
timestamp 1607319584
transform -1 0 1556 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1607319584
transform -1 0 1564 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_644
timestamp 1607319584
transform -1 0 1660 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_83
timestamp 1607319584
transform -1 0 1684 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_754
timestamp 1607319584
transform -1 0 1708 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_324
timestamp 1607319584
transform -1 0 1740 0 1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_75
timestamp 1607319584
transform -1 0 1780 0 1 2105
box -2 -3 42 103
use INVX1  INVX1_496
timestamp 1607319584
transform -1 0 1796 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_824
timestamp 1607319584
transform -1 0 1892 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_621
timestamp 1607319584
transform 1 0 1892 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_322
timestamp 1607319584
transform -1 0 1948 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_15
timestamp 1607319584
transform 1 0 1948 0 1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_148
timestamp 1607319584
transform -1 0 2012 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_214
timestamp 1607319584
transform -1 0 2044 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_68
timestamp 1607319584
transform -1 0 2068 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_3_0
timestamp 1607319584
transform -1 0 2076 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1607319584
transform -1 0 2084 0 1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_862
timestamp 1607319584
transform -1 0 2108 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_72
timestamp 1607319584
transform -1 0 2148 0 1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_719
timestamp 1607319584
transform 1 0 2148 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_74
timestamp 1607319584
transform -1 0 2212 0 1 2105
box -2 -3 42 103
use NOR2X1  NOR2X1_130
timestamp 1607319584
transform 1 0 2212 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_37
timestamp 1607319584
transform -1 0 2268 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_31
timestamp 1607319584
transform -1 0 2300 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_231
timestamp 1607319584
transform 1 0 2300 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_1156
timestamp 1607319584
transform -1 0 2364 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_368
timestamp 1607319584
transform -1 0 2380 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_822
timestamp 1607319584
transform -1 0 2476 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_619
timestamp 1607319584
transform 1 0 2476 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_146
timestamp 1607319584
transform -1 0 2532 0 1 2105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_30
timestamp 1607319584
transform 1 0 2532 0 1 2105
box -2 -3 74 103
use FILL  FILL_21_4_0
timestamp 1607319584
transform 1 0 2604 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_4_1
timestamp 1607319584
transform 1 0 2612 0 1 2105
box -2 -3 10 103
use BUFX4  BUFX4_75
timestamp 1607319584
transform 1 0 2620 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_78
timestamp 1607319584
transform 1 0 2652 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_36
timestamp 1607319584
transform 1 0 2684 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_325
timestamp 1607319584
transform 1 0 2716 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1607319584
transform 1 0 2748 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_689
timestamp 1607319584
transform -1 0 2868 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_293
timestamp 1607319584
transform 1 0 2868 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_238
timestamp 1607319584
transform -1 0 2924 0 1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_6
timestamp 1607319584
transform 1 0 2924 0 1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_71
timestamp 1607319584
transform -1 0 3004 0 1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_702
timestamp 1607319584
transform -1 0 3028 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_200
timestamp 1607319584
transform 1 0 3028 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_230
timestamp 1607319584
transform -1 0 3084 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_5_0
timestamp 1607319584
transform -1 0 3092 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_5_1
timestamp 1607319584
transform -1 0 3100 0 1 2105
box -2 -3 10 103
use AOI22X1  AOI22X1_3
timestamp 1607319584
transform -1 0 3140 0 1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_441
timestamp 1607319584
transform 1 0 3140 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_492
timestamp 1607319584
transform -1 0 3260 0 1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_20
timestamp 1607319584
transform 1 0 3260 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_26
timestamp 1607319584
transform 1 0 3292 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_70
timestamp 1607319584
transform -1 0 3356 0 1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_814
timestamp 1607319584
transform 1 0 3356 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_4
timestamp 1607319584
transform 1 0 3388 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_227
timestamp 1607319584
transform 1 0 3420 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_112
timestamp 1607319584
transform 1 0 3444 0 1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_942
timestamp 1607319584
transform -1 0 3524 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_154
timestamp 1607319584
transform 1 0 3524 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_203
timestamp 1607319584
transform 1 0 3540 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_25
timestamp 1607319584
transform -1 0 3596 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_6_0
timestamp 1607319584
transform 1 0 3596 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_6_1
timestamp 1607319584
transform 1 0 3604 0 1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_306
timestamp 1607319584
transform 1 0 3612 0 1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_305
timestamp 1607319584
transform 1 0 3660 0 1 2105
box -2 -3 50 103
use INVX1  INVX1_411
timestamp 1607319584
transform 1 0 3708 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_1199
timestamp 1607319584
transform -1 0 3756 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_215
timestamp 1607319584
transform 1 0 3756 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_37
timestamp 1607319584
transform -1 0 3812 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_815
timestamp 1607319584
transform -1 0 3844 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_31
timestamp 1607319584
transform 1 0 3844 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_209
timestamp 1607319584
transform -1 0 3900 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_30
timestamp 1607319584
transform -1 0 3916 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_481
timestamp 1607319584
transform -1 0 4012 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_980
timestamp 1607319584
transform 1 0 4012 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_413
timestamp 1607319584
transform 1 0 4044 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_189
timestamp 1607319584
transform -1 0 4116 0 1 2105
box -2 -3 50 103
use FILL  FILL_21_7_0
timestamp 1607319584
transform -1 0 4124 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_7_1
timestamp 1607319584
transform -1 0 4132 0 1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_140
timestamp 1607319584
transform -1 0 4180 0 1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_141
timestamp 1607319584
transform -1 0 4228 0 1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_1325
timestamp 1607319584
transform -1 0 4260 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_256
timestamp 1607319584
transform 1 0 4260 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_1044
timestamp 1607319584
transform 1 0 4276 0 1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_188
timestamp 1607319584
transform -1 0 4356 0 1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_482
timestamp 1607319584
transform 1 0 4356 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1607319584
transform -1 0 4476 0 1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_235
timestamp 1607319584
transform 1 0 4476 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_290
timestamp 1607319584
transform 1 0 4508 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1607319584
transform -1 0 4628 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_8_0
timestamp 1607319584
transform -1 0 4636 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_8_1
timestamp 1607319584
transform -1 0 4644 0 1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_24
timestamp 1607319584
transform -1 0 4668 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_66
timestamp 1607319584
transform -1 0 4716 0 1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_32
timestamp 1607319584
transform 1 0 4716 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_210
timestamp 1607319584
transform -1 0 4772 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_147
timestamp 1607319584
transform 1 0 4772 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_879
timestamp 1607319584
transform 1 0 4796 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_303
timestamp 1607319584
transform 1 0 4828 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_91
timestamp 1607319584
transform -1 0 4868 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_482
timestamp 1607319584
transform -1 0 4964 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_490
timestamp 1607319584
transform -1 0 5060 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_140
timestamp 1607319584
transform -1 0 5092 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1607319584
transform -1 0 5188 0 1 2105
box -2 -3 98 103
use FILL  FILL_22_1
timestamp 1607319584
transform 1 0 5188 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_980
timestamp 1607319584
transform -1 0 100 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_767
timestamp 1607319584
transform 1 0 100 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_766
timestamp 1607319584
transform -1 0 164 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_440
timestamp 1607319584
transform -1 0 196 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_964
timestamp 1607319584
transform 1 0 196 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_735
timestamp 1607319584
transform 1 0 292 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_734
timestamp 1607319584
transform -1 0 356 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_968
timestamp 1607319584
transform 1 0 356 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_249
timestamp 1607319584
transform 1 0 452 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_505
timestamp 1607319584
transform 1 0 468 0 -1 2305
box -2 -3 18 103
use BUFX4  BUFX4_439
timestamp 1607319584
transform 1 0 484 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1037
timestamp 1607319584
transform 1 0 516 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_0_0
timestamp 1607319584
transform 1 0 548 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1607319584
transform 1 0 556 0 -1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_749
timestamp 1607319584
transform 1 0 564 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1293
timestamp 1607319584
transform 1 0 588 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_24
timestamp 1607319584
transform 1 0 620 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_773
timestamp 1607319584
transform 1 0 668 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_772
timestamp 1607319584
transform 1 0 700 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_975
timestamp 1607319584
transform 1 0 732 0 -1 2305
box -2 -3 98 103
use INVX2  INVX2_5
timestamp 1607319584
transform 1 0 828 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_770
timestamp 1607319584
transform 1 0 844 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_771
timestamp 1607319584
transform -1 0 908 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_265
timestamp 1607319584
transform 1 0 908 0 -1 2305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_982
timestamp 1607319584
transform 1 0 956 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_1_0
timestamp 1607319584
transform -1 0 1060 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1607319584
transform -1 0 1068 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_409
timestamp 1607319584
transform -1 0 1100 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_378
timestamp 1607319584
transform 1 0 1100 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_733
timestamp 1607319584
transform 1 0 1116 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_732
timestamp 1607319584
transform 1 0 1148 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1166
timestamp 1607319584
transform 1 0 1180 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_197
timestamp 1607319584
transform -1 0 1236 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_738
timestamp 1607319584
transform 1 0 1236 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_739
timestamp 1607319584
transform -1 0 1300 0 -1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_56
timestamp 1607319584
transform -1 0 1340 0 -1 2305
box -2 -3 42 103
use AOI22X1  AOI22X1_36
timestamp 1607319584
transform 1 0 1340 0 -1 2305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_966
timestamp 1607319584
transform 1 0 1380 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_377
timestamp 1607319584
transform 1 0 1476 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_339
timestamp 1607319584
transform 1 0 1492 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1165
timestamp 1607319584
transform 1 0 1516 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_615
timestamp 1607319584
transform 1 0 1548 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_2_0
timestamp 1607319584
transform 1 0 1572 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1607319584
transform 1 0 1580 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_280
timestamp 1607319584
transform 1 0 1588 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_598
timestamp 1607319584
transform -1 0 1660 0 -1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_66
timestamp 1607319584
transform 1 0 1660 0 -1 2305
box -2 -3 42 103
use OAI21X1  OAI21X1_1284
timestamp 1607319584
transform -1 0 1732 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_740
timestamp 1607319584
transform -1 0 1756 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_290
timestamp 1607319584
transform -1 0 1788 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_143
timestamp 1607319584
transform -1 0 1812 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_460
timestamp 1607319584
transform -1 0 1836 0 -1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_35
timestamp 1607319584
transform 1 0 1836 0 -1 2305
box -2 -3 42 103
use AOI22X1  AOI22X1_19
timestamp 1607319584
transform -1 0 1916 0 -1 2305
box -2 -3 42 103
use BUFX4  BUFX4_322
timestamp 1607319584
transform -1 0 1948 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_124
timestamp 1607319584
transform 1 0 1948 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_667
timestamp 1607319584
transform -1 0 1996 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_135
timestamp 1607319584
transform 1 0 1996 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_6
timestamp 1607319584
transform -1 0 2052 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_133
timestamp 1607319584
transform 1 0 2052 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_3_0
timestamp 1607319584
transform -1 0 2084 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1607319584
transform -1 0 2092 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_292
timestamp 1607319584
transform -1 0 2124 0 -1 2305
box -2 -3 34 103
use INVX8  INVX8_9
timestamp 1607319584
transform -1 0 2164 0 -1 2305
box -2 -3 42 103
use MUX2X1  MUX2X1_272
timestamp 1607319584
transform -1 0 2212 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_601
timestamp 1607319584
transform -1 0 2236 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1155
timestamp 1607319584
transform -1 0 2268 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_289
timestamp 1607319584
transform 1 0 2268 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_7
timestamp 1607319584
transform 1 0 2300 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_367
timestamp 1607319584
transform -1 0 2348 0 -1 2305
box -2 -3 18 103
use BUFX4  BUFX4_77
timestamp 1607319584
transform 1 0 2348 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_5
timestamp 1607319584
transform -1 0 2412 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1607319584
transform 1 0 2412 0 -1 2305
box -2 -3 34 103
use INVX8  INVX8_16
timestamp 1607319584
transform 1 0 2444 0 -1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_408
timestamp 1607319584
transform 1 0 2484 0 -1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_49
timestamp 1607319584
transform 1 0 2508 0 -1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_546
timestamp 1607319584
transform -1 0 2572 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_4_0
timestamp 1607319584
transform -1 0 2580 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_4_1
timestamp 1607319584
transform -1 0 2588 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_63
timestamp 1607319584
transform -1 0 2620 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_72
timestamp 1607319584
transform -1 0 2652 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_62
timestamp 1607319584
transform -1 0 2684 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_49
timestamp 1607319584
transform -1 0 2716 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_51
timestamp 1607319584
transform 1 0 2716 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_73
timestamp 1607319584
transform 1 0 2748 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_48
timestamp 1607319584
transform -1 0 2812 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_162
timestamp 1607319584
transform -1 0 2860 0 -1 2305
box -2 -3 50 103
use INVX8  INVX8_1
timestamp 1607319584
transform -1 0 2900 0 -1 2305
box -2 -3 42 103
use NOR2X1  NOR2X1_32
timestamp 1607319584
transform -1 0 2924 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_29
timestamp 1607319584
transform 1 0 2924 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_199
timestamp 1607319584
transform 1 0 2940 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_31
timestamp 1607319584
transform -1 0 2996 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_291
timestamp 1607319584
transform 1 0 2996 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_11
timestamp 1607319584
transform -1 0 3052 0 -1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_161
timestamp 1607319584
transform -1 0 3100 0 -1 2305
box -2 -3 50 103
use FILL  FILL_22_5_0
timestamp 1607319584
transform 1 0 3100 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_5_1
timestamp 1607319584
transform 1 0 3108 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_68
timestamp 1607319584
transform 1 0 3116 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1007
timestamp 1607319584
transform -1 0 3180 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_219
timestamp 1607319584
transform -1 0 3196 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_484
timestamp 1607319584
transform -1 0 3292 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_212
timestamp 1607319584
transform 1 0 3292 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_34
timestamp 1607319584
transform -1 0 3348 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1008
timestamp 1607319584
transform -1 0 3380 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_220
timestamp 1607319584
transform 1 0 3380 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_500
timestamp 1607319584
transform -1 0 3492 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_220
timestamp 1607319584
transform 1 0 3492 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1607319584
transform -1 0 3548 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_21
timestamp 1607319584
transform 1 0 3548 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_22
timestamp 1607319584
transform -1 0 3596 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_6_0
timestamp 1607319584
transform -1 0 3604 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_6_1
timestamp 1607319584
transform -1 0 3612 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_135
timestamp 1607319584
transform -1 0 3644 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_50
timestamp 1607319584
transform 1 0 3644 0 -1 2305
box -2 -3 34 103
use INVX8  INVX8_7
timestamp 1607319584
transform 1 0 3676 0 -1 2305
box -2 -3 42 103
use MUX2X1  MUX2X1_224
timestamp 1607319584
transform -1 0 3764 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_547
timestamp 1607319584
transform -1 0 3788 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1091
timestamp 1607319584
transform -1 0 3820 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_532
timestamp 1607319584
transform -1 0 3844 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_129
timestamp 1607319584
transform 1 0 3844 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_103
timestamp 1607319584
transform -1 0 3900 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_303
timestamp 1607319584
transform -1 0 3916 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_813
timestamp 1607319584
transform -1 0 4012 0 -1 2305
box -2 -3 98 103
use BUFX4  BUFX4_136
timestamp 1607319584
transform -1 0 4044 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_138
timestamp 1607319584
transform -1 0 4076 0 -1 2305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_2
timestamp 1607319584
transform -1 0 4148 0 -1 2305
box -2 -3 74 103
use FILL  FILL_22_7_0
timestamp 1607319584
transform -1 0 4156 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_7_1
timestamp 1607319584
transform -1 0 4164 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_444
timestamp 1607319584
transform -1 0 4196 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_448
timestamp 1607319584
transform 1 0 4196 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_446
timestamp 1607319584
transform -1 0 4260 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_1200
timestamp 1607319584
transform -1 0 4292 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_649
timestamp 1607319584
transform 1 0 4292 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_412
timestamp 1607319584
transform 1 0 4316 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_223
timestamp 1607319584
transform 1 0 4332 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_45
timestamp 1607319584
transform -1 0 4388 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_445
timestamp 1607319584
transform -1 0 4420 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_783
timestamp 1607319584
transform 1 0 4420 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_1321
timestamp 1607319584
transform -1 0 4476 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_202
timestamp 1607319584
transform -1 0 4508 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_36
timestamp 1607319584
transform -1 0 4524 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1607319584
transform -1 0 4620 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_8_0
timestamp 1607319584
transform 1 0 4620 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_8_1
timestamp 1607319584
transform 1 0 4628 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_65
timestamp 1607319584
transform 1 0 4636 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_144
timestamp 1607319584
transform 1 0 4684 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_617
timestamp 1607319584
transform -1 0 4740 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_820
timestamp 1607319584
transform 1 0 4740 0 -1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_153
timestamp 1607319584
transform -1 0 4868 0 -1 2305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_71
timestamp 1607319584
transform -1 0 4940 0 -1 2305
box -2 -3 74 103
use BUFX4  BUFX4_139
timestamp 1607319584
transform -1 0 4972 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_501
timestamp 1607319584
transform 1 0 4972 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_221
timestamp 1607319584
transform 1 0 5068 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_188
timestamp 1607319584
transform -1 0 5124 0 -1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_44
timestamp 1607319584
transform -1 0 5196 0 -1 2305
box -2 -3 74 103
use BUFX2  BUFX2_6
timestamp 1607319584
transform -1 0 28 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1030
timestamp 1607319584
transform -1 0 124 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_761
timestamp 1607319584
transform 1 0 124 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_760
timestamp 1607319584
transform 1 0 156 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_977
timestamp 1607319584
transform 1 0 188 0 1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_23
timestamp 1607319584
transform -1 0 332 0 1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_743
timestamp 1607319584
transform 1 0 332 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_742
timestamp 1607319584
transform 1 0 364 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_969
timestamp 1607319584
transform 1 0 396 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_745
timestamp 1607319584
transform 1 0 492 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_0_0
timestamp 1607319584
transform -1 0 532 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1607319584
transform -1 0 540 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_744
timestamp 1607319584
transform -1 0 572 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_22
timestamp 1607319584
transform -1 0 620 0 1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_728
timestamp 1607319584
transform 1 0 620 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_983
timestamp 1607319584
transform 1 0 652 0 1 2305
box -2 -3 98 103
use INVX1  INVX1_442
timestamp 1607319584
transform 1 0 748 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_72
timestamp 1607319584
transform -1 0 788 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_757
timestamp 1607319584
transform 1 0 788 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_756
timestamp 1607319584
transform -1 0 852 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_680
timestamp 1607319584
transform -1 0 876 0 1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_217
timestamp 1607319584
transform 1 0 876 0 1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_219
timestamp 1607319584
transform 1 0 924 0 1 2305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_656
timestamp 1607319584
transform 1 0 972 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_1_0
timestamp 1607319584
transform 1 0 1068 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1607319584
transform 1 0 1076 0 1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_80
timestamp 1607319584
transform 1 0 1084 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_64
timestamp 1607319584
transform -1 0 1140 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_336
timestamp 1607319584
transform -1 0 1164 0 1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_121
timestamp 1607319584
transform -1 0 1212 0 1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_612
timestamp 1607319584
transform -1 0 1236 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_455
timestamp 1607319584
transform -1 0 1268 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_37
timestamp 1607319584
transform -1 0 1316 0 1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_841
timestamp 1607319584
transform -1 0 1348 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_123
timestamp 1607319584
transform 1 0 1348 0 1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_39
timestamp 1607319584
transform 1 0 1396 0 1 2305
box -2 -3 50 103
use INVX1  INVX1_53
timestamp 1607319584
transform -1 0 1460 0 1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_641
timestamp 1607319584
transform -1 0 1556 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_2_0
timestamp 1607319584
transform 1 0 1556 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1607319584
transform 1 0 1564 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_409
timestamp 1607319584
transform 1 0 1572 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1607319584
transform -1 0 1628 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_59
timestamp 1607319584
transform -1 0 1668 0 1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_616
timestamp 1607319584
transform -1 0 1692 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_239
timestamp 1607319584
transform 1 0 1692 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_16
timestamp 1607319584
transform 1 0 1716 0 1 2305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_832
timestamp 1607319584
transform -1 0 1852 0 1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_115
timestamp 1607319584
transform -1 0 1884 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_241
timestamp 1607319584
transform 1 0 1884 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_9
timestamp 1607319584
transform -1 0 1924 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_7
timestamp 1607319584
transform 1 0 1924 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_242
timestamp 1607319584
transform 1 0 1940 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_240
timestamp 1607319584
transform -1 0 1988 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_65
timestamp 1607319584
transform 1 0 1988 0 1 2305
box -2 -3 42 103
use AOI22X1  AOI22X1_55
timestamp 1607319584
transform 1 0 2028 0 1 2305
box -2 -3 42 103
use FILL  FILL_23_3_0
timestamp 1607319584
transform -1 0 2076 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1607319584
transform -1 0 2084 0 1 2305
box -2 -3 10 103
use BUFX4  BUFX4_157
timestamp 1607319584
transform -1 0 2116 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_352
timestamp 1607319584
transform -1 0 2148 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_46
timestamp 1607319584
transform 1 0 2148 0 1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_529
timestamp 1607319584
transform -1 0 2212 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_45
timestamp 1607319584
transform -1 0 2252 0 1 2305
box -2 -3 42 103
use BUFX4  BUFX4_351
timestamp 1607319584
transform -1 0 2284 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_54
timestamp 1607319584
transform -1 0 2324 0 1 2305
box -2 -3 42 103
use OAI21X1  OAI21X1_612
timestamp 1607319584
transform 1 0 2324 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_139
timestamp 1607319584
transform -1 0 2380 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_806
timestamp 1607319584
transform -1 0 2476 0 1 2305
box -2 -3 98 103
use BUFX4  BUFX4_4
timestamp 1607319584
transform -1 0 2508 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_29
timestamp 1607319584
transform 1 0 2508 0 1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_409
timestamp 1607319584
transform -1 0 2572 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_4_0
timestamp 1607319584
transform 1 0 2572 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_4_1
timestamp 1607319584
transform 1 0 2580 0 1 2305
box -2 -3 10 103
use BUFX4  BUFX4_1
timestamp 1607319584
transform 1 0 2588 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1607319584
transform 1 0 2620 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_354
timestamp 1607319584
transform -1 0 2700 0 1 2305
box -2 -3 50 103
use BUFX4  BUFX4_61
timestamp 1607319584
transform -1 0 2732 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_60
timestamp 1607319584
transform 1 0 2732 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_258
timestamp 1607319584
transform 1 0 2764 0 1 2305
box -2 -3 50 103
use BUFX4  BUFX4_74
timestamp 1607319584
transform -1 0 2844 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_497
timestamp 1607319584
transform 1 0 2844 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_217
timestamp 1607319584
transform 1 0 2940 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1607319584
transform -1 0 2996 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_288
timestamp 1607319584
transform 1 0 2996 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1607319584
transform 1 0 3028 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_349
timestamp 1607319584
transform -1 0 3092 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_5_0
timestamp 1607319584
transform -1 0 3100 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_5_1
timestamp 1607319584
transform -1 0 3108 0 1 2305
box -2 -3 10 103
use BUFX4  BUFX4_156
timestamp 1607319584
transform -1 0 3140 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_323
timestamp 1607319584
transform -1 0 3172 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_42
timestamp 1607319584
transform 1 0 3172 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_564
timestamp 1607319584
transform -1 0 3228 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_50
timestamp 1607319584
transform 1 0 3228 0 1 2305
box -2 -3 42 103
use AOI22X1  AOI22X1_51
timestamp 1607319584
transform -1 0 3308 0 1 2305
box -2 -3 42 103
use AOI22X1  AOI22X1_42
timestamp 1607319584
transform -1 0 3348 0 1 2305
box -2 -3 42 103
use AOI21X1  AOI21X1_28
timestamp 1607319584
transform 1 0 3348 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1607319584
transform -1 0 3404 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_442
timestamp 1607319584
transform -1 0 3428 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_508
timestamp 1607319584
transform -1 0 3524 0 1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_114
timestamp 1607319584
transform 1 0 3524 0 1 2305
box -2 -3 50 103
use NOR2X1  NOR2X1_30
timestamp 1607319584
transform -1 0 3596 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_6_0
timestamp 1607319584
transform -1 0 3604 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_6_1
timestamp 1607319584
transform -1 0 3612 0 1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_24
timestamp 1607319584
transform -1 0 3644 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_496
timestamp 1607319584
transform -1 0 3740 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_20
timestamp 1607319584
transform -1 0 3764 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_512
timestamp 1607319584
transform 1 0 3764 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_44
timestamp 1607319584
transform -1 0 3828 0 1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_138
timestamp 1607319584
transform 1 0 3828 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_611
timestamp 1607319584
transform -1 0 3884 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_805
timestamp 1607319584
transform 1 0 3884 0 1 2305
box -2 -3 98 103
use AOI22X1  AOI22X1_41
timestamp 1607319584
transform -1 0 4020 0 1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_495
timestamp 1607319584
transform -1 0 4044 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_40
timestamp 1607319584
transform -1 0 4084 0 1 2305
box -2 -3 42 103
use BUFX4  BUFX4_263
timestamp 1607319584
transform -1 0 4116 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_7_0
timestamp 1607319584
transform 1 0 4116 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_7_1
timestamp 1607319584
transform 1 0 4124 0 1 2305
box -2 -3 10 103
use BUFX4  BUFX4_276
timestamp 1607319584
transform 1 0 4132 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_822
timestamp 1607319584
transform -1 0 4196 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_289
timestamp 1607319584
transform -1 0 4220 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_234
timestamp 1607319584
transform -1 0 4252 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1607319584
transform 1 0 4252 0 1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_210
timestamp 1607319584
transform 1 0 4348 0 1 2305
box -2 -3 50 103
use BUFX4  BUFX4_277
timestamp 1607319584
transform 1 0 4396 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_39
timestamp 1607319584
transform 1 0 4428 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_31
timestamp 1607319584
transform -1 0 4484 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_238
timestamp 1607319584
transform 1 0 4484 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_821
timestamp 1607319584
transform 1 0 4508 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_511
timestamp 1607319584
transform -1 0 4636 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_8_0
timestamp 1607319584
transform -1 0 4644 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_8_1
timestamp 1607319584
transform -1 0 4652 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_503
timestamp 1607319584
transform -1 0 4748 0 1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_209
timestamp 1607319584
transform 1 0 4748 0 1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_1072
timestamp 1607319584
transform 1 0 4796 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_240
timestamp 1607319584
transform -1 0 4844 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_1220
timestamp 1607319584
transform 1 0 4844 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_511
timestamp 1607319584
transform -1 0 4900 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_671
timestamp 1607319584
transform 1 0 4900 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_831
timestamp 1607319584
transform -1 0 5020 0 1 2305
box -2 -3 98 103
use INVX1  INVX1_284
timestamp 1607319584
transform 1 0 5020 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_142
timestamp 1607319584
transform 1 0 5036 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_439
timestamp 1607319584
transform -1 0 5076 0 1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_114
timestamp 1607319584
transform -1 0 5108 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1607319584
transform -1 0 5132 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_237
timestamp 1607319584
transform 1 0 5132 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_231
timestamp 1607319584
transform 1 0 5156 0 1 2305
box -2 -3 34 103
use FILL  FILL_24_1
timestamp 1607319584
transform 1 0 5188 0 1 2305
box -2 -3 10 103
use BUFX2  BUFX2_2
timestamp 1607319584
transform -1 0 28 0 -1 2505
box -2 -3 26 103
use BUFX2  BUFX2_4
timestamp 1607319584
transform -1 0 52 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1028
timestamp 1607319584
transform -1 0 148 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1026
timestamp 1607319584
transform -1 0 244 0 -1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_211
timestamp 1607319584
transform -1 0 268 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_985
timestamp 1607319584
transform -1 0 364 0 -1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_210
timestamp 1607319584
transform 1 0 364 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_987
timestamp 1607319584
transform 1 0 388 0 -1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_213
timestamp 1607319584
transform 1 0 484 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_250
timestamp 1607319584
transform 1 0 508 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_0_0
timestamp 1607319584
transform 1 0 524 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_0_1
timestamp 1607319584
transform 1 0 532 0 -1 2505
box -2 -3 10 103
use MUX2X1  MUX2X1_184
timestamp 1607319584
transform 1 0 540 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_1038
timestamp 1607319584
transform 1 0 588 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_474
timestamp 1607319584
transform -1 0 644 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_729
timestamp 1607319584
transform 1 0 644 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_961
timestamp 1607319584
transform 1 0 676 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_1230
timestamp 1607319584
transform 1 0 772 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_75
timestamp 1607319584
transform 1 0 804 0 -1 2505
box -2 -3 50 103
use INVX1  INVX1_441
timestamp 1607319584
transform 1 0 852 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_1229
timestamp 1607319584
transform 1 0 868 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_62
timestamp 1607319584
transform 1 0 900 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_78
timestamp 1607319584
transform 1 0 932 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_649
timestamp 1607319584
transform 1 0 956 0 -1 2505
box -2 -3 98 103
use FILL  FILL_24_1_0
timestamp 1607319584
transform 1 0 1052 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_1_1
timestamp 1607319584
transform 1 0 1060 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_986
timestamp 1607319584
transform 1 0 1068 0 -1 2505
box -2 -3 98 103
use BUFX4  BUFX4_141
timestamp 1607319584
transform 1 0 1164 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_328
timestamp 1607319584
transform -1 0 1244 0 -1 2505
box -2 -3 50 103
use BUFX4  BUFX4_103
timestamp 1607319584
transform -1 0 1276 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_263
timestamp 1607319584
transform -1 0 1300 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_143
timestamp 1607319584
transform 1 0 1300 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_145
timestamp 1607319584
transform -1 0 1364 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_144
timestamp 1607319584
transform 1 0 1364 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_816
timestamp 1607319584
transform 1 0 1396 0 -1 2505
box -2 -3 98 103
use AOI21X1  AOI21X1_106
timestamp 1607319584
transform 1 0 1492 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_132
timestamp 1607319584
transform 1 0 1524 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_2_0
timestamp 1607319584
transform -1 0 1556 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_2_1
timestamp 1607319584
transform -1 0 1564 0 -1 2505
box -2 -3 10 103
use BUFX4  BUFX4_353
timestamp 1607319584
transform -1 0 1596 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1607319584
transform 1 0 1596 0 -1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_243
timestamp 1607319584
transform -1 0 1636 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_12
timestamp 1607319584
transform -1 0 1652 0 -1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_253
timestamp 1607319584
transform -1 0 1676 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_469
timestamp 1607319584
transform 1 0 1676 0 -1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_249
timestamp 1607319584
transform -1 0 1716 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_252
timestamp 1607319584
transform -1 0 1740 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_98
timestamp 1607319584
transform -1 0 1764 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_160
timestamp 1607319584
transform -1 0 1796 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_477
timestamp 1607319584
transform 1 0 1796 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_39
timestamp 1607319584
transform 1 0 1820 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_478
timestamp 1607319584
transform -1 0 1884 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1257
timestamp 1607319584
transform -1 0 1916 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_340
timestamp 1607319584
transform -1 0 1940 0 -1 2505
box -2 -3 26 103
use INVX8  INVX8_13
timestamp 1607319584
transform 1 0 1940 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_69
timestamp 1607319584
transform 1 0 1980 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_685
timestamp 1607319584
transform -1 0 2044 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_684
timestamp 1607319584
transform 1 0 2044 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_3_0
timestamp 1607319584
transform -1 0 2076 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_3_1
timestamp 1607319584
transform -1 0 2084 0 -1 2505
box -2 -3 10 103
use BUFX4  BUFX4_159
timestamp 1607319584
transform -1 0 2116 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_8
timestamp 1607319584
transform 1 0 2116 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_73
timestamp 1607319584
transform 1 0 2156 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_5
timestamp 1607319584
transform 1 0 2196 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_32
timestamp 1607319584
transform -1 0 2260 0 -1 2505
box -2 -3 42 103
use AOI21X1  AOI21X1_32
timestamp 1607319584
transform 1 0 2260 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_53
timestamp 1607319584
transform 1 0 2292 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_26
timestamp 1607319584
transform 1 0 2332 0 -1 2505
box -2 -3 42 103
use BUFX4  BUFX4_320
timestamp 1607319584
transform 1 0 2372 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_33
timestamp 1607319584
transform 1 0 2404 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_443
timestamp 1607319584
transform 1 0 2444 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_34
timestamp 1607319584
transform -1 0 2508 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_391
timestamp 1607319584
transform -1 0 2532 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_350
timestamp 1607319584
transform 1 0 2532 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_25
timestamp 1607319584
transform -1 0 2604 0 -1 2505
box -2 -3 42 103
use FILL  FILL_24_4_0
timestamp 1607319584
transform -1 0 2612 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_4_1
timestamp 1607319584
transform -1 0 2620 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_1264
timestamp 1607319584
transform -1 0 2652 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_353
timestamp 1607319584
transform -1 0 2700 0 -1 2505
box -2 -3 50 103
use AOI22X1  AOI22X1_47
timestamp 1607319584
transform -1 0 2740 0 -1 2505
box -2 -3 42 103
use BUFX4  BUFX4_158
timestamp 1607319584
transform -1 0 2772 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_225
timestamp 1607319584
transform 1 0 2772 0 -1 2505
box -2 -3 50 103
use MUX2X1  MUX2X1_257
timestamp 1607319584
transform 1 0 2820 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_1136
timestamp 1607319584
transform -1 0 2900 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_305
timestamp 1607319584
transform 1 0 2900 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_14
timestamp 1607319584
transform -1 0 2964 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_374
timestamp 1607319584
transform 1 0 2964 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_24
timestamp 1607319584
transform -1 0 3028 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_23
timestamp 1607319584
transform 1 0 3028 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_13
timestamp 1607319584
transform 1 0 3068 0 -1 2505
box -2 -3 42 103
use FILL  FILL_24_5_0
timestamp 1607319584
transform -1 0 3116 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_5_1
timestamp 1607319584
transform -1 0 3124 0 -1 2505
box -2 -3 10 103
use AOI22X1  AOI22X1_62
timestamp 1607319584
transform -1 0 3164 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_650
timestamp 1607319584
transform 1 0 3164 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_63
timestamp 1607319584
transform 1 0 3188 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_11
timestamp 1607319584
transform -1 0 3268 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_288
timestamp 1607319584
transform -1 0 3292 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1263
timestamp 1607319584
transform 1 0 3292 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_10
timestamp 1607319584
transform -1 0 3364 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_64
timestamp 1607319584
transform -1 0 3404 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_31
timestamp 1607319584
transform -1 0 3444 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_426
timestamp 1607319584
transform -1 0 3468 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1135
timestamp 1607319584
transform -1 0 3500 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_347
timestamp 1607319584
transform -1 0 3516 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_214
timestamp 1607319584
transform 1 0 3516 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_36
timestamp 1607319584
transform -1 0 3572 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_717
timestamp 1607319584
transform -1 0 3596 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_6_0
timestamp 1607319584
transform 1 0 3596 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_6_1
timestamp 1607319584
transform 1 0 3604 0 -1 2505
box -2 -3 10 103
use NAND3X1  NAND3X1_1
timestamp 1607319584
transform 1 0 3612 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_486
timestamp 1607319584
transform 1 0 3644 0 -1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_841
timestamp 1607319584
transform -1 0 3764 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_354
timestamp 1607319584
transform 1 0 3764 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_250
timestamp 1607319584
transform 1 0 3796 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_321
timestamp 1607319584
transform 1 0 3820 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_43
timestamp 1607319584
transform 1 0 3852 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_61
timestamp 1607319584
transform -1 0 3932 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_633
timestamp 1607319584
transform -1 0 3956 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_60
timestamp 1607319584
transform 1 0 3956 0 -1 2505
box -2 -3 42 103
use BUFX4  BUFX4_155
timestamp 1607319584
transform 1 0 3996 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_21
timestamp 1607319584
transform -1 0 4068 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_357
timestamp 1607319584
transform -1 0 4092 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_20
timestamp 1607319584
transform -1 0 4132 0 -1 2505
box -2 -3 42 103
use FILL  FILL_24_7_0
timestamp 1607319584
transform -1 0 4140 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_7_1
timestamp 1607319584
transform -1 0 4148 0 -1 2505
box -2 -3 10 103
use AOI22X1  AOI22X1_30
timestamp 1607319584
transform -1 0 4188 0 -1 2505
box -2 -3 42 103
use BUFX4  BUFX4_270
timestamp 1607319584
transform -1 0 4220 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_807
timestamp 1607319584
transform 1 0 4220 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_1219
timestamp 1607319584
transform -1 0 4348 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_431
timestamp 1607319584
transform -1 0 4364 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_613
timestamp 1607319584
transform 1 0 4364 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_140
timestamp 1607319584
transform -1 0 4420 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_202
timestamp 1607319584
transform 1 0 4420 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_943
timestamp 1607319584
transform -1 0 4484 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_113
timestamp 1607319584
transform 1 0 4484 0 -1 2505
box -2 -3 50 103
use NAND2X1  NAND2X1_33
timestamp 1607319584
transform 1 0 4532 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_944
timestamp 1607319584
transform -1 0 4588 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_211
timestamp 1607319584
transform -1 0 4620 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_155
timestamp 1607319584
transform -1 0 4636 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_8_0
timestamp 1607319584
transform 1 0 4636 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_8_1
timestamp 1607319584
transform 1 0 4644 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_483
timestamp 1607319584
transform 1 0 4652 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_1071
timestamp 1607319584
transform 1 0 4748 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_35
timestamp 1607319584
transform 1 0 4780 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_27
timestamp 1607319584
transform -1 0 4836 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_510
timestamp 1607319584
transform -1 0 4860 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_41
timestamp 1607319584
transform 1 0 4860 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_37
timestamp 1607319584
transform 1 0 4884 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_509
timestamp 1607319584
transform -1 0 5004 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_493
timestamp 1607319584
transform -1 0 5100 0 -1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_139
timestamp 1607319584
transform 1 0 5100 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_111
timestamp 1607319584
transform -1 0 5156 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_26
timestamp 1607319584
transform 1 0 5156 0 -1 2505
box -2 -3 34 103
use FILL  FILL_25_1
timestamp 1607319584
transform -1 0 5196 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_988
timestamp 1607319584
transform 1 0 4 0 1 2505
box -2 -3 98 103
use AOI21X1  AOI21X1_173
timestamp 1607319584
transform -1 0 132 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_214
timestamp 1607319584
transform -1 0 156 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_991
timestamp 1607319584
transform 1 0 156 0 1 2505
box -2 -3 98 103
use AOI21X1  AOI21X1_170
timestamp 1607319584
transform -1 0 284 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_652
timestamp 1607319584
transform 1 0 284 0 1 2505
box -2 -3 98 103
use AOI21X1  AOI21X1_60
timestamp 1607319584
transform 1 0 380 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_76
timestamp 1607319584
transform 1 0 412 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_172
timestamp 1607319584
transform 1 0 436 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_889
timestamp 1607319584
transform -1 0 500 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_383
timestamp 1607319584
transform -1 0 524 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_0_0
timestamp 1607319584
transform -1 0 532 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_0_1
timestamp 1607319584
transform -1 0 540 0 1 2505
box -2 -3 10 103
use MUX2X1  MUX2X1_73
timestamp 1607319584
transform -1 0 588 0 1 2505
box -2 -3 50 103
use BUFX4  BUFX4_142
timestamp 1607319584
transform 1 0 588 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_681
timestamp 1607319584
transform -1 0 644 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_654
timestamp 1607319584
transform -1 0 740 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_590
timestamp 1607319584
transform 1 0 740 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1209
timestamp 1607319584
transform 1 0 764 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_953
timestamp 1607319584
transform -1 0 828 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_1145
timestamp 1607319584
transform -1 0 860 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_73
timestamp 1607319584
transform -1 0 884 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_57
timestamp 1607319584
transform -1 0 916 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_357
timestamp 1607319584
transform -1 0 932 0 1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_646
timestamp 1607319584
transform -1 0 1028 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_414
timestamp 1607319584
transform 1 0 1028 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_1_0
timestamp 1607319584
transform 1 0 1060 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_1_1
timestamp 1607319584
transform 1 0 1068 0 1 2505
box -2 -3 10 103
use AOI21X1  AOI21X1_171
timestamp 1607319584
transform 1 0 1076 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_212
timestamp 1607319584
transform -1 0 1132 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_89
timestamp 1607319584
transform -1 0 1156 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_57
timestamp 1607319584
transform -1 0 1196 0 1 2505
box -2 -3 42 103
use MUX2X1  MUX2X1_273
timestamp 1607319584
transform 1 0 1196 0 1 2505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_808
timestamp 1607319584
transform 1 0 1244 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_495
timestamp 1607319584
transform 1 0 1340 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_614
timestamp 1607319584
transform 1 0 1356 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_141
timestamp 1607319584
transform -1 0 1412 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_311
timestamp 1607319584
transform 1 0 1412 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_739
timestamp 1607319584
transform 1 0 1444 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1283
timestamp 1607319584
transform -1 0 1500 0 1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_368
timestamp 1607319584
transform 1 0 1500 0 1 2505
box -2 -3 50 103
use FILL  FILL_25_2_0
timestamp 1607319584
transform 1 0 1548 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_2_1
timestamp 1607319584
transform 1 0 1556 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_392
timestamp 1607319584
transform 1 0 1564 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_13
timestamp 1607319584
transform 1 0 1660 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_72
timestamp 1607319584
transform -1 0 1716 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_53
timestamp 1607319584
transform -1 0 1748 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_55
timestamp 1607319584
transform -1 0 1780 0 1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_349
timestamp 1607319584
transform -1 0 1828 0 1 2505
box -2 -3 50 103
use MUX2X1  MUX2X1_351
timestamp 1607319584
transform 1 0 1828 0 1 2505
box -2 -3 50 103
use NAND2X1  NAND2X1_711
timestamp 1607319584
transform 1 0 1876 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_27
timestamp 1607319584
transform 1 0 1900 0 1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_67
timestamp 1607319584
transform -1 0 1980 0 1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_52
timestamp 1607319584
transform -1 0 2020 0 1 2505
box -2 -3 42 103
use BUFX4  BUFX4_54
timestamp 1607319584
transform 1 0 2020 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_581
timestamp 1607319584
transform 1 0 2052 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_3_0
timestamp 1607319584
transform -1 0 2084 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_3_1
timestamp 1607319584
transform -1 0 2092 0 1 2505
box -2 -3 10 103
use AOI22X1  AOI22X1_7
timestamp 1607319584
transform -1 0 2132 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_271
timestamp 1607319584
transform 1 0 2132 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_512
timestamp 1607319584
transform -1 0 2252 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_718
timestamp 1607319584
transform 1 0 2252 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_40
timestamp 1607319584
transform -1 0 2300 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_76
timestamp 1607319584
transform -1 0 2332 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_81
timestamp 1607319584
transform 1 0 2332 0 1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_9
timestamp 1607319584
transform -1 0 2404 0 1 2505
box -2 -3 42 103
use NAND3X1  NAND3X1_6
timestamp 1607319584
transform -1 0 2436 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_799
timestamp 1607319584
transform 1 0 2436 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_510
timestamp 1607319584
transform 1 0 2468 0 1 2505
box -2 -3 98 103
use AOI21X1  AOI21X1_30
timestamp 1607319584
transform 1 0 2564 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_4_0
timestamp 1607319584
transform 1 0 2596 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_4_1
timestamp 1607319584
transform 1 0 2604 0 1 2505
box -2 -3 10 103
use NOR2X1  NOR2X1_38
timestamp 1607319584
transform 1 0 2612 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_580
timestamp 1607319584
transform -1 0 2660 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_12
timestamp 1607319584
transform -1 0 2700 0 1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_22
timestamp 1607319584
transform -1 0 2740 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_223
timestamp 1607319584
transform -1 0 2764 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_3
timestamp 1607319584
transform -1 0 2796 0 1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_4
timestamp 1607319584
transform 1 0 2796 0 1 2505
box -2 -3 42 103
use INVX1  INVX1_348
timestamp 1607319584
transform 1 0 2836 0 1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_502
timestamp 1607319584
transform -1 0 2948 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_222
timestamp 1607319584
transform 1 0 2948 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_44
timestamp 1607319584
transform -1 0 3004 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_52
timestamp 1607319584
transform 1 0 3004 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_476
timestamp 1607319584
transform -1 0 3052 0 1 2505
box -2 -3 18 103
use FILL  FILL_25_5_0
timestamp 1607319584
transform -1 0 3060 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_5_1
timestamp 1607319584
transform -1 0 3068 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_504
timestamp 1607319584
transform -1 0 3164 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_224
timestamp 1607319584
transform 1 0 3164 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_46
timestamp 1607319584
transform -1 0 3220 0 1 2505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_31
timestamp 1607319584
transform -1 0 3292 0 1 2505
box -2 -3 74 103
use NOR2X1  NOR2X1_28
timestamp 1607319584
transform -1 0 3316 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1607319584
transform -1 0 3348 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_494
timestamp 1607319584
transform 1 0 3348 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_579
timestamp 1607319584
transform -1 0 3468 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_844
timestamp 1607319584
transform 1 0 3468 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_1618
timestamp 1607319584
transform -1 0 3524 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_273
timestamp 1607319584
transform 1 0 3524 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_6_0
timestamp 1607319584
transform 1 0 3620 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_6_1
timestamp 1607319584
transform 1 0 3628 0 1 2505
box -2 -3 10 103
use INVX1  INVX1_19
timestamp 1607319584
transform 1 0 3636 0 1 2505
box -2 -3 18 103
use AOI22X1  AOI22X1_1
timestamp 1607319584
transform -1 0 3692 0 1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_804
timestamp 1607319584
transform 1 0 3692 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_813
timestamp 1607319584
transform -1 0 3756 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_215
timestamp 1607319584
transform 1 0 3756 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_65
timestamp 1607319584
transform 1 0 3780 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1607319584
transform -1 0 3836 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_28
timestamp 1607319584
transform 1 0 3836 0 1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_385
timestamp 1607319584
transform -1 0 3948 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_216
timestamp 1607319584
transform 1 0 3948 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_281
timestamp 1607319584
transform -1 0 4068 0 1 2505
box -2 -3 98 103
use BUFX4  BUFX4_223
timestamp 1607319584
transform -1 0 4100 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_7_0
timestamp 1607319584
transform -1 0 4108 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_7_1
timestamp 1607319584
transform -1 0 4116 0 1 2505
box -2 -3 10 103
use MUX2X1  MUX2X1_320
timestamp 1607319584
transform -1 0 4164 0 1 2505
box -2 -3 50 103
use AOI21X1  AOI21X1_105
timestamp 1607319584
transform 1 0 4164 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_131
timestamp 1607319584
transform -1 0 4220 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_815
timestamp 1607319584
transform 1 0 4220 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_670
timestamp 1607319584
transform -1 0 4340 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_230
timestamp 1607319584
transform 1 0 4340 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_232
timestamp 1607319584
transform -1 0 4404 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_28
timestamp 1607319584
transform -1 0 4436 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_372
timestamp 1607319584
transform 1 0 4436 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_507
timestamp 1607319584
transform -1 0 4556 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_373
timestamp 1607319584
transform 1 0 4556 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_25
timestamp 1607319584
transform 1 0 4580 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1607319584
transform -1 0 4636 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_8_0
timestamp 1607319584
transform -1 0 4644 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_8_1
timestamp 1607319584
transform -1 0 4652 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_491
timestamp 1607319584
transform -1 0 4748 0 1 2505
box -2 -3 98 103
use BUFX4  BUFX4_11
timestamp 1607319584
transform 1 0 4748 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_21
timestamp 1607319584
transform 1 0 4780 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1607319584
transform -1 0 4836 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_156
timestamp 1607319584
transform 1 0 4836 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_219
timestamp 1607319584
transform 1 0 4852 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_29
timestamp 1607319584
transform -1 0 4916 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_828
timestamp 1607319584
transform -1 0 5012 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_506
timestamp 1607319584
transform 1 0 5012 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_304
timestamp 1607319584
transform 1 0 5108 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_40
timestamp 1607319584
transform 1 0 5132 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_324
timestamp 1607319584
transform -1 0 5180 0 1 2505
box -2 -3 26 103
use FILL  FILL_26_1
timestamp 1607319584
transform 1 0 5180 0 1 2505
box -2 -3 10 103
use FILL  FILL_26_2
timestamp 1607319584
transform 1 0 5188 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_801
timestamp 1607319584
transform 1 0 4 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_123
timestamp 1607319584
transform 1 0 100 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_98
timestamp 1607319584
transform -1 0 156 0 -1 2705
box -2 -3 34 103
use BUFX2  BUFX2_7
timestamp 1607319584
transform -1 0 180 0 -1 2705
box -2 -3 26 103
use MUX2X1  MUX2X1_6
timestamp 1607319584
transform -1 0 228 0 -1 2705
box -2 -3 50 103
use AOI21X1  AOI21X1_58
timestamp 1607319584
transform 1 0 228 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_59
timestamp 1607319584
transform 1 0 260 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_75
timestamp 1607319584
transform -1 0 316 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_217
timestamp 1607319584
transform 1 0 316 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_176
timestamp 1607319584
transform -1 0 372 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_642
timestamp 1607319584
transform 1 0 372 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_101
timestamp 1607319584
transform 1 0 468 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_410
timestamp 1607319584
transform 1 0 484 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_85
timestamp 1607319584
transform -1 0 540 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_0_0
timestamp 1607319584
transform -1 0 548 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_0_1
timestamp 1607319584
transform -1 0 556 0 -1 2705
box -2 -3 10 103
use NAND2X1  NAND2X1_88
timestamp 1607319584
transform -1 0 580 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1031
timestamp 1607319584
transform -1 0 676 0 -1 2705
box -2 -3 98 103
use MUX2X1  MUX2X1_7
timestamp 1607319584
transform -1 0 724 0 -1 2705
box -2 -3 50 103
use INVX1  INVX1_421
timestamp 1607319584
transform -1 0 740 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_647
timestamp 1607319584
transform -1 0 836 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_415
timestamp 1607319584
transform 1 0 836 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_165
timestamp 1607319584
transform -1 0 884 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_643
timestamp 1607319584
transform -1 0 980 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_411
timestamp 1607319584
transform 1 0 980 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_86
timestamp 1607319584
transform -1 0 1036 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_1_0
timestamp 1607319584
transform 1 0 1036 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_1_1
timestamp 1607319584
transform 1 0 1044 0 -1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_175
timestamp 1607319584
transform 1 0 1052 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_216
timestamp 1607319584
transform -1 0 1108 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_990
timestamp 1607319584
transform 1 0 1108 0 -1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_319
timestamp 1607319584
transform -1 0 1228 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_894
timestamp 1607319584
transform -1 0 1260 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_388
timestamp 1607319584
transform 1 0 1260 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_213
timestamp 1607319584
transform 1 0 1356 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_68
timestamp 1607319584
transform 1 0 1372 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_6
timestamp 1607319584
transform 1 0 1404 0 -1 2705
box -2 -3 18 103
use OAI22X1  OAI22X1_1
timestamp 1607319584
transform 1 0 1420 0 -1 2705
box -2 -3 42 103
use INVX1  INVX1_8
timestamp 1607319584
transform -1 0 1476 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_122
timestamp 1607319584
transform -1 0 1500 0 -1 2705
box -2 -3 26 103
use MUX2X1  MUX2X1_76
timestamp 1607319584
transform -1 0 1548 0 -1 2705
box -2 -3 50 103
use NAND2X1  NAND2X1_90
timestamp 1607319584
transform -1 0 1572 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_2_0
timestamp 1607319584
transform 1 0 1572 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_2_1
timestamp 1607319584
transform 1 0 1580 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_396
timestamp 1607319584
transform 1 0 1588 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1001
timestamp 1607319584
transform 1 0 1684 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_78
timestamp 1607319584
transform 1 0 1716 0 -1 2705
box -2 -3 50 103
use INVX1  INVX1_470
timestamp 1607319584
transform 1 0 1764 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_1258
timestamp 1607319584
transform 1 0 1780 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_400
timestamp 1607319584
transform 1 0 1812 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_10
timestamp 1607319584
transform 1 0 1908 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_8
timestamp 1607319584
transform -1 0 1964 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_321
timestamp 1607319584
transform 1 0 1964 0 -1 2705
box -2 -3 50 103
use AOI21X1  AOI21X1_2
timestamp 1607319584
transform 1 0 2012 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_4
timestamp 1607319584
transform -1 0 2068 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_3_0
timestamp 1607319584
transform -1 0 2076 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_3_1
timestamp 1607319584
transform -1 0 2084 0 -1 2705
box -2 -3 10 103
use NAND2X1  NAND2X1_297
timestamp 1607319584
transform -1 0 2108 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_394
timestamp 1607319584
transform -1 0 2204 0 -1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_14
timestamp 1607319584
transform -1 0 2228 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_15
timestamp 1607319584
transform 1 0 2228 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_16
timestamp 1607319584
transform -1 0 2276 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_17
timestamp 1607319584
transform 1 0 2276 0 -1 2705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_94
timestamp 1607319584
transform -1 0 2372 0 -1 2705
box -2 -3 74 103
use OAI21X1  OAI21X1_105
timestamp 1607319584
transform 1 0 2372 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_106
timestamp 1607319584
transform -1 0 2436 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_417
timestamp 1607319584
transform 1 0 2436 0 -1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_47
timestamp 1607319584
transform -1 0 2556 0 -1 2705
box -2 -3 26 103
use BUFX4  BUFX4_47
timestamp 1607319584
transform -1 0 2588 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_4_0
timestamp 1607319584
transform 1 0 2588 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_4_1
timestamp 1607319584
transform 1 0 2596 0 -1 2705
box -2 -3 10 103
use BUFX4  BUFX4_46
timestamp 1607319584
transform 1 0 2604 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_45
timestamp 1607319584
transform -1 0 2668 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_44
timestamp 1607319584
transform 1 0 2668 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_407
timestamp 1607319584
transform 1 0 2700 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_441
timestamp 1607319584
transform 1 0 2732 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_812
timestamp 1607319584
transform -1 0 2860 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_810
timestamp 1607319584
transform 1 0 2860 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_198
timestamp 1607319584
transform 1 0 2892 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_27
timestamp 1607319584
transform -1 0 2940 0 -1 2705
box -2 -3 18 103
use BUFX4  BUFX4_111
timestamp 1607319584
transform -1 0 2972 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_387
timestamp 1607319584
transform 1 0 2972 0 -1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_845
timestamp 1607319584
transform 1 0 3068 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_5_0
timestamp 1607319584
transform 1 0 3092 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_5_1
timestamp 1607319584
transform 1 0 3100 0 -1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_196
timestamp 1607319584
transform 1 0 3108 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_41
timestamp 1607319584
transform -1 0 3172 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_488
timestamp 1607319584
transform 1 0 3172 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_475
timestamp 1607319584
transform 1 0 3268 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_216
timestamp 1607319584
transform 1 0 3284 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1607319584
transform -1 0 3340 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_802
timestamp 1607319584
transform -1 0 3372 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1619
timestamp 1607319584
transform -1 0 3404 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_274
timestamp 1607319584
transform 1 0 3404 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_78
timestamp 1607319584
transform 1 0 3500 0 -1 2705
box -2 -3 18 103
use BUFX4  BUFX4_304
timestamp 1607319584
transform -1 0 3548 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_57
timestamp 1607319584
transform -1 0 3596 0 -1 2705
box -2 -3 50 103
use FILL  FILL_26_6_0
timestamp 1607319584
transform 1 0 3596 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_6_1
timestamp 1607319584
transform 1 0 3604 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_866
timestamp 1607319584
transform 1 0 3612 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_55
timestamp 1607319584
transform -1 0 3692 0 -1 2705
box -2 -3 50 103
use NAND2X1  NAND2X1_290
timestamp 1607319584
transform 1 0 3692 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_225
timestamp 1607319584
transform 1 0 3716 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_3
timestamp 1607319584
transform 1 0 3740 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_1
timestamp 1607319584
transform -1 0 3796 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_393
timestamp 1607319584
transform -1 0 3892 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_361
timestamp 1607319584
transform -1 0 3916 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_287
timestamp 1607319584
transform -1 0 3948 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_282
timestamp 1607319584
transform -1 0 4044 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_360
timestamp 1607319584
transform 1 0 4044 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_286
timestamp 1607319584
transform -1 0 4100 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_331
timestamp 1607319584
transform -1 0 4132 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_7_0
timestamp 1607319584
transform -1 0 4140 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_7_1
timestamp 1607319584
transform -1 0 4148 0 -1 2705
box -2 -3 10 103
use NAND3X1  NAND3X1_5
timestamp 1607319584
transform -1 0 4180 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_191
timestamp 1607319584
transform 1 0 4180 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_248
timestamp 1607319584
transform 1 0 4212 0 -1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_93
timestamp 1607319584
transform -1 0 4316 0 -1 2705
box -2 -3 74 103
use NOR2X1  NOR2X1_334
timestamp 1607319584
transform 1 0 4316 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_264
timestamp 1607319584
transform -1 0 4372 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_161
timestamp 1607319584
transform -1 0 4404 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_226
timestamp 1607319584
transform 1 0 4404 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_35
timestamp 1607319584
transform 1 0 4436 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_213
timestamp 1607319584
transform -1 0 4492 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_163
timestamp 1607319584
transform -1 0 4524 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_283
timestamp 1607319584
transform -1 0 4540 0 -1 2705
box -2 -3 18 103
use BUFX4  BUFX4_162
timestamp 1607319584
transform -1 0 4572 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_331
timestamp 1607319584
transform -1 0 4596 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_252
timestamp 1607319584
transform 1 0 4596 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_8_0
timestamp 1607319584
transform -1 0 4628 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_8_1
timestamp 1607319584
transform -1 0 4636 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_803
timestamp 1607319584
transform -1 0 4668 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_214
timestamp 1607319584
transform 1 0 4668 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_297
timestamp 1607319584
transform -1 0 4788 0 -1 2705
box -2 -3 98 103
use BUFX4  BUFX4_164
timestamp 1607319584
transform 1 0 4788 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_499
timestamp 1607319584
transform -1 0 4916 0 -1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_464
timestamp 1607319584
transform 1 0 4916 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_824
timestamp 1607319584
transform 1 0 4940 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_826
timestamp 1607319584
transform 1 0 4964 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_1449
timestamp 1607319584
transform -1 0 5020 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_830
timestamp 1607319584
transform 1 0 5020 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1607319584
transform -1 0 5068 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_251
timestamp 1607319584
transform 1 0 5068 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_333
timestamp 1607319584
transform 1 0 5092 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_263
timestamp 1607319584
transform -1 0 5148 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_410
timestamp 1607319584
transform -1 0 5164 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_775
timestamp 1607319584
transform -1 0 5188 0 -1 2705
box -2 -3 26 103
use FILL  FILL_27_1
timestamp 1607319584
transform -1 0 5196 0 -1 2705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_88
timestamp 1607319584
transform 1 0 4 0 1 2705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_100
timestamp 1607319584
transform 1 0 76 0 1 2705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_650
timestamp 1607319584
transform 1 0 148 0 1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_74
timestamp 1607319584
transform -1 0 268 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_651
timestamp 1607319584
transform 1 0 268 0 1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_314
timestamp 1607319584
transform -1 0 388 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_645
timestamp 1607319584
transform 1 0 388 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_293
timestamp 1607319584
transform 1 0 484 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_413
timestamp 1607319584
transform 1 0 500 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_0_0
timestamp 1607319584
transform 1 0 532 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_0_1
timestamp 1607319584
transform 1 0 540 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_1081
timestamp 1607319584
transform 1 0 548 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_521
timestamp 1607319584
transform 1 0 580 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_653
timestamp 1607319584
transform -1 0 700 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_655
timestamp 1607319584
transform 1 0 700 0 1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_659
timestamp 1607319584
transform -1 0 820 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_63
timestamp 1607319584
transform 1 0 820 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_79
timestamp 1607319584
transform 1 0 852 0 1 2705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_72
timestamp 1607319584
transform 1 0 876 0 1 2705
box -2 -3 74 103
use BUFX4  BUFX4_88
timestamp 1607319584
transform 1 0 948 0 1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_33
timestamp 1607319584
transform 1 0 980 0 1 2705
box -2 -3 74 103
use FILL  FILL_27_1_0
timestamp 1607319584
transform 1 0 1052 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_1_1
timestamp 1607319584
transform 1 0 1060 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_730
timestamp 1607319584
transform 1 0 1068 0 1 2705
box -2 -3 98 103
use AOI21X1  AOI21X1_66
timestamp 1607319584
transform 1 0 1164 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_84
timestamp 1607319584
transform 1 0 1196 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_102
timestamp 1607319584
transform 1 0 1220 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_546
timestamp 1607319584
transform -1 0 1276 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_106
timestamp 1607319584
transform -1 0 1292 0 1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_722
timestamp 1607319584
transform -1 0 1388 0 1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_9
timestamp 1607319584
transform -1 0 1412 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_408
timestamp 1607319584
transform -1 0 1444 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_104
timestamp 1607319584
transform 1 0 1444 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_548
timestamp 1607319584
transform -1 0 1500 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_234
timestamp 1607319584
transform -1 0 1516 0 1 2705
box -2 -3 18 103
use FILL  FILL_27_2_0
timestamp 1607319584
transform -1 0 1524 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_2_1
timestamp 1607319584
transform -1 0 1532 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_724
timestamp 1607319584
transform -1 0 1628 0 1 2705
box -2 -3 98 103
use AOI21X1  AOI21X1_4
timestamp 1607319584
transform 1 0 1628 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1607319584
transform -1 0 1684 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_435
timestamp 1607319584
transform -1 0 1708 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_86
timestamp 1607319584
transform -1 0 1740 0 1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_157
timestamp 1607319584
transform 1 0 1740 0 1 2705
box -2 -3 50 103
use NAND2X1  NAND2X1_712
timestamp 1607319584
transform -1 0 1812 0 1 2705
box -2 -3 26 103
use MUX2X1  MUX2X1_159
timestamp 1607319584
transform 1 0 1812 0 1 2705
box -2 -3 50 103
use AOI21X1  AOI21X1_67
timestamp 1607319584
transform 1 0 1860 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_731
timestamp 1607319584
transform 1 0 1892 0 1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_85
timestamp 1607319584
transform -1 0 2012 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_388
timestamp 1607319584
transform -1 0 2036 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_84
timestamp 1607319584
transform 1 0 2036 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_3_0
timestamp 1607319584
transform 1 0 2068 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_3_1
timestamp 1607319584
transform 1 0 2076 0 1 2705
box -2 -3 10 103
use MUX2X1  MUX2X1_124
timestamp 1607319584
transform 1 0 2084 0 1 2705
box -2 -3 50 103
use OAI21X1  OAI21X1_958
timestamp 1607319584
transform -1 0 2164 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_1
timestamp 1607319584
transform -1 0 2180 0 1 2705
box -2 -3 18 103
use INVX1  INVX1_170
timestamp 1607319584
transform -1 0 2196 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_547
timestamp 1607319584
transform 1 0 2196 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_103
timestamp 1607319584
transform -1 0 2252 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_723
timestamp 1607319584
transform -1 0 2348 0 1 2705
box -2 -3 98 103
use MUX2X1  MUX2X1_126
timestamp 1607319584
transform 1 0 2348 0 1 2705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_276
timestamp 1607319584
transform 1 0 2396 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_206
timestamp 1607319584
transform 1 0 2492 0 1 2705
box -2 -3 18 103
use BUFX4  BUFX4_22
timestamp 1607319584
transform -1 0 2540 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_26
timestamp 1607319584
transform 1 0 2540 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_811
timestamp 1607319584
transform 1 0 2556 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_4_0
timestamp 1607319584
transform 1 0 2588 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_4_1
timestamp 1607319584
transform 1 0 2596 0 1 2705
box -2 -3 10 103
use BUFX4  BUFX4_70
timestamp 1607319584
transform 1 0 2604 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_71
timestamp 1607319584
transform 1 0 2636 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_409
timestamp 1607319584
transform 1 0 2668 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_90
timestamp 1607319584
transform 1 0 2764 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_89
timestamp 1607319584
transform -1 0 2828 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_224
timestamp 1607319584
transform -1 0 2852 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_74
timestamp 1607319584
transform 1 0 2852 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1607319584
transform 1 0 2884 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_401
timestamp 1607319584
transform -1 0 3012 0 1 2705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_4
timestamp 1607319584
transform -1 0 3084 0 1 2705
box -2 -3 74 103
use NAND2X1  NAND2X1_107
timestamp 1607319584
transform -1 0 3108 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_5_0
timestamp 1607319584
transform 1 0 3108 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_5_1
timestamp 1607319584
transform 1 0 3116 0 1 2705
box -2 -3 10 103
use NAND2X1  NAND2X1_8
timestamp 1607319584
transform 1 0 3124 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_67
timestamp 1607319584
transform -1 0 3180 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_149
timestamp 1607319584
transform 1 0 3180 0 1 2705
box -2 -3 18 103
use BUFX4  BUFX4_59
timestamp 1607319584
transform -1 0 3228 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_69
timestamp 1607319584
transform -1 0 3260 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_58
timestamp 1607319584
transform 1 0 3260 0 1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_75
timestamp 1607319584
transform 1 0 3292 0 1 2705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_89
timestamp 1607319584
transform 1 0 3364 0 1 2705
box -2 -3 74 103
use BUFX4  BUFX4_326
timestamp 1607319584
transform -1 0 3468 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_327
timestamp 1607319584
transform -1 0 3500 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1607319584
transform -1 0 3532 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_329
timestamp 1607319584
transform 1 0 3532 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_20
timestamp 1607319584
transform -1 0 3596 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_6_0
timestamp 1607319584
transform 1 0 3596 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_6_1
timestamp 1607319584
transform 1 0 3604 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_1057
timestamp 1607319584
transform 1 0 3612 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_496
timestamp 1607319584
transform 1 0 3644 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_21
timestamp 1607319584
transform 1 0 3668 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_328
timestamp 1607319584
transform 1 0 3700 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_269
timestamp 1607319584
transform -1 0 3828 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1610
timestamp 1607319584
transform -1 0 3860 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1611
timestamp 1607319584
transform -1 0 3892 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_865
timestamp 1607319584
transform 1 0 3892 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_289
timestamp 1607319584
transform 1 0 3924 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_1604
timestamp 1607319584
transform 1 0 3948 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1605
timestamp 1607319584
transform -1 0 4012 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_266
timestamp 1607319584
transform -1 0 4108 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_7_0
timestamp 1607319584
transform 1 0 4108 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_7_1
timestamp 1607319584
transform 1 0 4116 0 1 2705
box -2 -3 10 103
use MUX2X1  MUX2X1_51
timestamp 1607319584
transform 1 0 4124 0 1 2705
box -2 -3 50 103
use MUX2X1  MUX2X1_50
timestamp 1607319584
transform -1 0 4220 0 1 2705
box -2 -3 50 103
use OAI21X1  OAI21X1_859
timestamp 1607319584
transform 1 0 4220 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_282
timestamp 1607319584
transform 1 0 4252 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_170
timestamp 1607319584
transform -1 0 4372 0 1 2705
box -2 -3 98 103
use BUFX4  BUFX4_333
timestamp 1607319584
transform -1 0 4404 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_332
timestamp 1607319584
transform 1 0 4404 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_485
timestamp 1607319584
transform 1 0 4436 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_832
timestamp 1607319584
transform -1 0 4564 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_206
timestamp 1607319584
transform -1 0 4596 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_254
timestamp 1607319584
transform 1 0 4596 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_8_0
timestamp 1607319584
transform -1 0 4628 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_8_1
timestamp 1607319584
transform -1 0 4636 0 1 2705
box -2 -3 10 103
use MUX2X1  MUX2X1_98
timestamp 1607319584
transform -1 0 4684 0 1 2705
box -2 -3 50 103
use NOR2X1  NOR2X1_370
timestamp 1607319584
transform -1 0 4708 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_294
timestamp 1607319584
transform -1 0 4740 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1607319584
transform -1 0 4836 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_1028
timestamp 1607319584
transform 1 0 4836 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_330
timestamp 1607319584
transform -1 0 4900 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_923
timestamp 1607319584
transform 1 0 4900 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_335
timestamp 1607319584
transform -1 0 4964 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_1451
timestamp 1607319584
transform 1 0 4964 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_161
timestamp 1607319584
transform 1 0 4996 0 1 2705
box -2 -3 98 103
use BUFX4  BUFX4_334
timestamp 1607319584
transform -1 0 5124 0 1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_63
timestamp 1607319584
transform 1 0 5124 0 1 2705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_809
timestamp 1607319584
transform -1 0 100 0 -1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_4
timestamp 1607319584
transform 1 0 100 0 -1 2905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_769
timestamp 1607319584
transform 1 0 148 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_802
timestamp 1607319584
transform 1 0 244 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_608
timestamp 1607319584
transform 1 0 340 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_135
timestamp 1607319584
transform -1 0 396 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_113
timestamp 1607319584
transform 1 0 396 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_775
timestamp 1607319584
transform 1 0 420 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_429
timestamp 1607319584
transform 1 0 516 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_0_0
timestamp 1607319584
transform 1 0 532 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_0_1
timestamp 1607319584
transform 1 0 540 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_803
timestamp 1607319584
transform 1 0 548 0 -1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_77
timestamp 1607319584
transform 1 0 644 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_175
timestamp 1607319584
transform 1 0 668 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_609
timestamp 1607319584
transform 1 0 684 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_136
timestamp 1607319584
transform -1 0 740 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1217
timestamp 1607319584
transform -1 0 772 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_452
timestamp 1607319584
transform 1 0 772 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_766
timestamp 1607319584
transform -1 0 900 0 -1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_177
timestamp 1607319584
transform 1 0 900 0 -1 2905
box -2 -3 50 103
use AOI22X1  AOI22X1_37
timestamp 1607319584
transform -1 0 988 0 -1 2905
box -2 -3 42 103
use BUFX4  BUFX4_361
timestamp 1607319584
transform -1 0 1020 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_270
timestamp 1607319584
transform -1 0 1068 0 -1 2905
box -2 -3 50 103
use FILL  FILL_28_1_0
timestamp 1607319584
transform 1 0 1068 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_1_1
timestamp 1607319584
transform 1 0 1076 0 -1 2905
box -2 -3 10 103
use MUX2X1  MUX2X1_268
timestamp 1607319584
transform 1 0 1084 0 -1 2905
box -2 -3 50 103
use BUFX4  BUFX4_362
timestamp 1607319584
transform -1 0 1164 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1150
timestamp 1607319584
transform -1 0 1196 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_408
timestamp 1607319584
transform 1 0 1196 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_88
timestamp 1607319584
transform 1 0 1292 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1607319584
transform -1 0 1356 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_411
timestamp 1607319584
transform 1 0 1356 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_94
timestamp 1607319584
transform 1 0 1452 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1607319584
transform -1 0 1516 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_367
timestamp 1607319584
transform -1 0 1540 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_938
timestamp 1607319584
transform 1 0 1540 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_2_0
timestamp 1607319584
transform 1 0 1572 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_2_1
timestamp 1607319584
transform 1 0 1580 0 -1 2905
box -2 -3 10 103
use MUX2X1  MUX2X1_77
timestamp 1607319584
transform 1 0 1588 0 -1 2905
box -2 -3 50 103
use MUX2X1  MUX2X1_318
timestamp 1607319584
transform 1 0 1636 0 -1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_103
timestamp 1607319584
transform 1 0 1684 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1607319584
transform -1 0 1748 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_416
timestamp 1607319584
transform -1 0 1844 0 -1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_350
timestamp 1607319584
transform 1 0 1844 0 -1 2905
box -2 -3 50 103
use BUFX4  BUFX4_174
timestamp 1607319584
transform 1 0 1892 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1260
timestamp 1607319584
transform -1 0 1956 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_319
timestamp 1607319584
transform -1 0 2004 0 -1 2905
box -2 -3 50 103
use BUFX4  BUFX4_25
timestamp 1607319584
transform -1 0 2036 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_873
timestamp 1607319584
transform 1 0 2036 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_3_0
timestamp 1607319584
transform -1 0 2076 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_3_1
timestamp 1607319584
transform -1 0 2084 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_85
timestamp 1607319584
transform -1 0 2100 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_66
timestamp 1607319584
transform 1 0 2100 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1607319584
transform -1 0 2156 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_386
timestamp 1607319584
transform -1 0 2252 0 -1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_61
timestamp 1607319584
transform -1 0 2300 0 -1 2905
box -2 -3 50 103
use INVX1  INVX1_362
timestamp 1607319584
transform 1 0 2300 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_726
timestamp 1607319584
transform -1 0 2412 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_550
timestamp 1607319584
transform 1 0 2412 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_106
timestamp 1607319584
transform -1 0 2468 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_847
timestamp 1607319584
transform -1 0 2492 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1621
timestamp 1607319584
transform -1 0 2524 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_125
timestamp 1607319584
transform 1 0 2524 0 -1 2905
box -2 -3 50 103
use FILL  FILL_28_4_0
timestamp 1607319584
transform -1 0 2580 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_4_1
timestamp 1607319584
transform -1 0 2588 0 -1 2905
box -2 -3 10 103
use MUX2X1  MUX2X1_153
timestamp 1607319584
transform -1 0 2636 0 -1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_960
timestamp 1607319584
transform -1 0 2668 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_172
timestamp 1607319584
transform -1 0 2684 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_755
timestamp 1607319584
transform -1 0 2780 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_563
timestamp 1607319584
transform 1 0 2780 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1607319584
transform -1 0 2836 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_154
timestamp 1607319584
transform 1 0 2836 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_153
timestamp 1607319584
transform -1 0 2900 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_177
timestamp 1607319584
transform 1 0 2900 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_111
timestamp 1607319584
transform -1 0 2980 0 -1 2905
box -2 -3 50 103
use MUX2X1  MUX2X1_109
timestamp 1607319584
transform -1 0 3028 0 -1 2905
box -2 -3 50 103
use INVX1  INVX1_426
timestamp 1607319584
transform -1 0 3044 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_551
timestamp 1607319584
transform 1 0 3044 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_17
timestamp 1607319584
transform 1 0 3076 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_5_0
timestamp 1607319584
transform -1 0 3100 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_5_1
timestamp 1607319584
transform -1 0 3108 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_727
timestamp 1607319584
transform -1 0 3204 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_937
timestamp 1607319584
transform 1 0 3204 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_56
timestamp 1607319584
transform 1 0 3236 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_240
timestamp 1607319584
transform 1 0 3268 0 -1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_807
timestamp 1607319584
transform -1 0 3340 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_366
timestamp 1607319584
transform 1 0 3340 0 -1 2905
box -2 -3 26 103
use MUX2X1  MUX2X1_239
timestamp 1607319584
transform 1 0 3364 0 -1 2905
box -2 -3 50 103
use MUX2X1  MUX2X1_201
timestamp 1607319584
transform -1 0 3460 0 -1 2905
box -2 -3 50 103
use NOR2X1  NOR2X1_5
timestamp 1607319584
transform 1 0 3460 0 -1 2905
box -2 -3 26 103
use BUFX4  BUFX4_97
timestamp 1607319584
transform -1 0 3516 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_152
timestamp 1607319584
transform 1 0 3516 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_808
timestamp 1607319584
transform -1 0 3572 0 -1 2905
box -2 -3 26 103
use INVX8  INVX8_5
timestamp 1607319584
transform 1 0 3572 0 -1 2905
box -2 -3 42 103
use FILL  FILL_28_6_0
timestamp 1607319584
transform 1 0 3612 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_6_1
timestamp 1607319584
transform 1 0 3620 0 -1 2905
box -2 -3 10 103
use MUX2X1  MUX2X1_199
timestamp 1607319584
transform 1 0 3628 0 -1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_1058
timestamp 1607319584
transform -1 0 3708 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_200
timestamp 1607319584
transform -1 0 3740 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_236
timestamp 1607319584
transform 1 0 3740 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_259
timestamp 1607319584
transform -1 0 3804 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_215
timestamp 1607319584
transform -1 0 3836 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_224
timestamp 1607319584
transform 1 0 3836 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_23
timestamp 1607319584
transform 1 0 3868 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_806
timestamp 1607319584
transform 1 0 3900 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1112
timestamp 1607319584
transform 1 0 3924 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_147
timestamp 1607319584
transform -1 0 4004 0 -1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_791
timestamp 1607319584
transform 1 0 4004 0 -1 2905
box -2 -3 26 103
use MUX2X1  MUX2X1_145
timestamp 1607319584
transform -1 0 4076 0 -1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_827
timestamp 1607319584
transform 1 0 4076 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_7_0
timestamp 1607319584
transform -1 0 4116 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_7_1
timestamp 1607319584
transform -1 0 4124 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_985
timestamp 1607319584
transform -1 0 4156 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_137
timestamp 1607319584
transform 1 0 4156 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_197
timestamp 1607319584
transform -1 0 4196 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_986
timestamp 1607319584
transform -1 0 4228 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_813
timestamp 1607319584
transform 1 0 4228 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_610
timestamp 1607319584
transform -1 0 4284 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_239
timestamp 1607319584
transform 1 0 4284 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_804
timestamp 1607319584
transform -1 0 4396 0 -1 2905
box -2 -3 98 103
use BUFX4  BUFX4_180
timestamp 1607319584
transform -1 0 4428 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1027
timestamp 1607319584
transform 1 0 4428 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_176
timestamp 1607319584
transform 1 0 4460 0 -1 2905
box -2 -3 50 103
use MUX2X1  MUX2X1_49
timestamp 1607319584
transform 1 0 4508 0 -1 2905
box -2 -3 50 103
use MUX2X1  MUX2X1_99
timestamp 1607319584
transform -1 0 4604 0 -1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_821
timestamp 1607319584
transform 1 0 4604 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_8_0
timestamp 1607319584
transform -1 0 4636 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_8_1
timestamp 1607319584
transform -1 0 4644 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_1446
timestamp 1607319584
transform -1 0 4676 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_198
timestamp 1607319584
transform -1 0 4692 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_1444
timestamp 1607319584
transform 1 0 4692 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_819
timestamp 1607319584
transform -1 0 4748 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_326
timestamp 1607319584
transform -1 0 4764 0 -1 2905
box -2 -3 18 103
use BUFX4  BUFX4_27
timestamp 1607319584
transform -1 0 4796 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_858
timestamp 1607319584
transform 1 0 4796 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_171
timestamp 1607319584
transform 1 0 4828 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_135
timestamp 1607319584
transform -1 0 4940 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_163
timestamp 1607319584
transform -1 0 5036 0 -1 2905
box -2 -3 98 103
use INVX1  INVX1_70
timestamp 1607319584
transform -1 0 5052 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_1442
timestamp 1607319584
transform 1 0 5052 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1607319584
transform -1 0 5180 0 -1 2905
box -2 -3 98 103
use FILL  FILL_29_1
timestamp 1607319584
transform -1 0 5188 0 -1 2905
box -2 -3 10 103
use FILL  FILL_29_2
timestamp 1607319584
transform -1 0 5196 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_794
timestamp 1607319584
transform -1 0 100 0 1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_115
timestamp 1607319584
transform 1 0 100 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_91
timestamp 1607319584
transform -1 0 156 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_125
timestamp 1607319584
transform 1 0 156 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_99
timestamp 1607319584
transform -1 0 212 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_450
timestamp 1607319584
transform -1 0 244 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_774
timestamp 1607319584
transform 1 0 244 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_111
timestamp 1607319584
transform 1 0 340 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_580
timestamp 1607319584
transform 1 0 356 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_579
timestamp 1607319584
transform -1 0 420 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_3
timestamp 1607319584
transform -1 0 468 0 1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_582
timestamp 1607319584
transform 1 0 468 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_581
timestamp 1607319584
transform -1 0 532 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_0_0
timestamp 1607319584
transform -1 0 540 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_0_1
timestamp 1607319584
transform -1 0 548 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_899
timestamp 1607319584
transform -1 0 580 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_451
timestamp 1607319584
transform 1 0 580 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_130
timestamp 1607319584
transform -1 0 644 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_61
timestamp 1607319584
transform -1 0 676 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_269
timestamp 1607319584
transform 1 0 676 0 1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_1152
timestamp 1607319584
transform 1 0 724 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_963
timestamp 1607319584
transform -1 0 788 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_597
timestamp 1607319584
transform 1 0 788 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_453
timestamp 1607319584
transform 1 0 812 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_449
timestamp 1607319584
transform 1 0 844 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_80
timestamp 1607319584
transform -1 0 924 0 1 2905
box -2 -3 50 103
use NOR2X1  NOR2X1_108
timestamp 1607319584
transform 1 0 924 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_86
timestamp 1607319584
transform -1 0 980 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_104
timestamp 1607319584
transform -1 0 1012 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_128
timestamp 1607319584
transform 1 0 1012 0 1 2905
box -2 -3 50 103
use FILL  FILL_29_1_0
timestamp 1607319584
transform 1 0 1060 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_1_1
timestamp 1607319584
transform 1 0 1068 0 1 2905
box -2 -3 10 103
use BUFX4  BUFX4_363
timestamp 1607319584
transform 1 0 1076 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_70
timestamp 1607319584
transform 1 0 1108 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_88
timestamp 1607319584
transform -1 0 1164 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_595
timestamp 1607319584
transform -1 0 1188 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_734
timestamp 1607319584
transform -1 0 1284 0 1 2905
box -2 -3 98 103
use BUFX4  BUFX4_356
timestamp 1607319584
transform 1 0 1284 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_84
timestamp 1607319584
transform 1 0 1316 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1607319584
transform 1 0 1348 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_406
timestamp 1607319584
transform 1 0 1380 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_342
timestamp 1607319584
transform 1 0 1476 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_410
timestamp 1607319584
transform 1 0 1492 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_2_0
timestamp 1607319584
transform 1 0 1588 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_2_1
timestamp 1607319584
transform 1 0 1596 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_874
timestamp 1607319584
transform 1 0 1604 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_298
timestamp 1607319584
transform 1 0 1636 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_91
timestamp 1607319584
transform -1 0 1692 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_92
timestamp 1607319584
transform -1 0 1724 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_209
timestamp 1607319584
transform 1 0 1724 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_193
timestamp 1607319584
transform -1 0 1788 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_168
timestamp 1607319584
transform 1 0 1788 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_167
timestamp 1607319584
transform 1 0 1820 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_448
timestamp 1607319584
transform 1 0 1852 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_714
timestamp 1607319584
transform -1 0 1972 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_185
timestamp 1607319584
transform -1 0 2004 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_85
timestamp 1607319584
transform 1 0 2004 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_107
timestamp 1607319584
transform -1 0 2060 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_3_0
timestamp 1607319584
transform 1 0 2060 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_3_1
timestamp 1607319584
transform 1 0 2068 0 1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_765
timestamp 1607319584
transform 1 0 2076 0 1 2905
box -2 -3 98 103
use MUX2X1  MUX2X1_222
timestamp 1607319584
transform 1 0 2172 0 1 2905
box -2 -3 50 103
use MUX2X1  MUX2X1_221
timestamp 1607319584
transform 1 0 2220 0 1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_19
timestamp 1607319584
transform -1 0 2292 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_528
timestamp 1607319584
transform -1 0 2316 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1088
timestamp 1607319584
transform -1 0 2348 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_757
timestamp 1607319584
transform 1 0 2348 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_300
timestamp 1607319584
transform 1 0 2444 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_565
timestamp 1607319584
transform 1 0 2460 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_63
timestamp 1607319584
transform 1 0 2492 0 1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_121
timestamp 1607319584
transform -1 0 2564 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_222
timestamp 1607319584
transform -1 0 2588 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_4_0
timestamp 1607319584
transform 1 0 2588 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_4_1
timestamp 1607319584
transform 1 0 2596 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_994
timestamp 1607319584
transform 1 0 2604 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_151
timestamp 1607319584
transform -1 0 2684 0 1 2905
box -2 -3 50 103
use OAI21X1  OAI21X1_1216
timestamp 1607319584
transform -1 0 2716 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_317
timestamp 1607319584
transform -1 0 2764 0 1 2905
box -2 -3 50 103
use NAND2X1  NAND2X1_123
timestamp 1607319584
transform 1 0 2764 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_567
timestamp 1607319584
transform -1 0 2820 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_428
timestamp 1607319584
transform -1 0 2836 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_759
timestamp 1607319584
transform -1 0 2932 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_665
timestamp 1607319584
transform -1 0 2956 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1215
timestamp 1607319584
transform -1 0 2988 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_427
timestamp 1607319584
transform -1 0 3004 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_743
timestamp 1607319584
transform -1 0 3100 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_5_0
timestamp 1607319584
transform 1 0 3100 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_5_1
timestamp 1607319584
transform 1 0 3108 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_559
timestamp 1607319584
transform 1 0 3116 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_115
timestamp 1607319584
transform -1 0 3172 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_390
timestamp 1607319584
transform 1 0 3172 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_105
timestamp 1607319584
transform 1 0 3196 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_83
timestamp 1607319584
transform -1 0 3252 0 1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_238
timestamp 1607319584
transform 1 0 3252 0 1 2905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_763
timestamp 1607319584
transform 1 0 3300 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_395
timestamp 1607319584
transform -1 0 3492 0 1 2905
box -2 -3 98 103
use AOI21X1  AOI21X1_3
timestamp 1607319584
transform -1 0 3524 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_1375
timestamp 1607319584
transform 1 0 3524 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1607319584
transform 1 0 3556 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_6_0
timestamp 1607319584
transform 1 0 3652 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_6_1
timestamp 1607319584
transform 1 0 3660 0 1 2905
box -2 -3 10 103
use INVX1  INVX1_387
timestamp 1607319584
transform 1 0 3668 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_497
timestamp 1607319584
transform -1 0 3708 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1175
timestamp 1607319584
transform 1 0 3708 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_206
timestamp 1607319584
transform -1 0 3772 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_848
timestamp 1607319584
transform 1 0 3772 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1622
timestamp 1607319584
transform -1 0 3828 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_270
timestamp 1607319584
transform -1 0 3844 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_277
timestamp 1607319584
transform 1 0 3844 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_805
timestamp 1607319584
transform -1 0 3964 0 1 2905
box -2 -3 26 103
use MUX2X1  MUX2X1_287
timestamp 1607319584
transform 1 0 3964 0 1 2905
box -2 -3 50 103
use BUFX4  BUFX4_262
timestamp 1607319584
transform -1 0 4044 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_253
timestamp 1607319584
transform -1 0 4076 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_204
timestamp 1607319584
transform -1 0 4108 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_555
timestamp 1607319584
transform 1 0 4108 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_7_0
timestamp 1607319584
transform 1 0 4132 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_7_1
timestamp 1607319584
transform 1 0 4140 0 1 2905
box -2 -3 10 103
use BUFX4  BUFX4_222
timestamp 1607319584
transform 1 0 4148 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_419
timestamp 1607319584
transform 1 0 4180 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_418
timestamp 1607319584
transform 1 0 4204 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_238
timestamp 1607319584
transform -1 0 4260 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_278
timestamp 1607319584
transform 1 0 4260 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_336
timestamp 1607319584
transform 1 0 4292 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_266
timestamp 1607319584
transform -1 0 4348 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_172
timestamp 1607319584
transform -1 0 4444 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_71
timestamp 1607319584
transform -1 0 4460 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_162
timestamp 1607319584
transform -1 0 4556 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_825
timestamp 1607319584
transform 1 0 4556 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_1450
timestamp 1607319584
transform -1 0 4612 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_463
timestamp 1607319584
transform -1 0 4636 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_8_0
timestamp 1607319584
transform -1 0 4644 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_8_1
timestamp 1607319584
transform -1 0 4652 0 1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_205
timestamp 1607319584
transform -1 0 4684 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_250
timestamp 1607319584
transform 1 0 4684 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1607319584
transform -1 0 4804 0 1 2905
box -2 -3 98 103
use BUFX4  BUFX4_390
timestamp 1607319584
transform -1 0 4836 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_265
timestamp 1607319584
transform 1 0 4836 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_243
timestamp 1607319584
transform 1 0 4868 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_335
timestamp 1607319584
transform -1 0 4924 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_351
timestamp 1607319584
transform -1 0 4948 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_281
timestamp 1607319584
transform 1 0 4948 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1607319584
transform -1 0 5068 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_817
timestamp 1607319584
transform -1 0 5092 0 1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_61
timestamp 1607319584
transform -1 0 5164 0 1 2905
box -2 -3 74 103
use AOI21X1  AOI21X1_256
timestamp 1607319584
transform 1 0 5164 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_793
timestamp 1607319584
transform -1 0 100 0 -1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_324
timestamp 1607319584
transform -1 0 124 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_114
timestamp 1607319584
transform 1 0 4 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_90
timestamp 1607319584
transform -1 0 60 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_601
timestamp 1607319584
transform -1 0 92 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_898
timestamp 1607319584
transform 1 0 92 0 1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_2
timestamp 1607319584
transform -1 0 172 0 -1 3105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_785
timestamp 1607319584
transform -1 0 268 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_110
timestamp 1607319584
transform -1 0 140 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_786
timestamp 1607319584
transform -1 0 236 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_112
timestamp 1607319584
transform 1 0 268 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_89
timestamp 1607319584
transform -1 0 324 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_777
timestamp 1607319584
transform 1 0 236 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_570
timestamp 1607319584
transform 1 0 324 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_569
timestamp 1607319584
transform -1 0 388 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_585
timestamp 1607319584
transform -1 0 420 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_586
timestamp 1607319584
transform 1 0 332 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_107
timestamp 1607319584
transform -1 0 396 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_325
timestamp 1607319584
transform -1 0 420 0 1 3105
box -2 -3 26 103
use MUX2X1  MUX2X1_1
timestamp 1607319584
transform 1 0 420 0 -1 3105
box -2 -3 50 103
use BUFX4  BUFX4_108
timestamp 1607319584
transform 1 0 468 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_0_0
timestamp 1607319584
transform 1 0 500 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_0_1
timestamp 1607319584
transform 1 0 508 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_596
timestamp 1607319584
transform 1 0 420 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_595
timestamp 1607319584
transform -1 0 484 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_98
timestamp 1607319584
transform -1 0 508 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_78
timestamp 1607319584
transform -1 0 540 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_750
timestamp 1607319584
transform 1 0 516 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_0_0
timestamp 1607319584
transform -1 0 548 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_0_1
timestamp 1607319584
transform -1 0 556 0 1 3105
box -2 -3 10 103
use BUFX4  BUFX4_106
timestamp 1607319584
transform -1 0 588 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_758
timestamp 1607319584
transform 1 0 588 0 1 3105
box -2 -3 98 103
use INVX1  INVX1_365
timestamp 1607319584
transform 1 0 612 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_596
timestamp 1607319584
transform -1 0 652 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1151
timestamp 1607319584
transform -1 0 684 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_122
timestamp 1607319584
transform -1 0 708 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_364
timestamp 1607319584
transform 1 0 708 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_566
timestamp 1607319584
transform -1 0 716 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_363
timestamp 1607319584
transform -1 0 740 0 -1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_742
timestamp 1607319584
transform -1 0 836 0 -1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_394
timestamp 1607319584
transform -1 0 740 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_668
timestamp 1607319584
transform -1 0 764 0 1 3105
box -2 -3 26 103
use MUX2X1  MUX2X1_79
timestamp 1607319584
transform -1 0 812 0 1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_558
timestamp 1607319584
transform -1 0 868 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_81
timestamp 1607319584
transform 1 0 868 0 -1 3105
box -2 -3 50 103
use NAND2X1  NAND2X1_114
timestamp 1607319584
transform 1 0 812 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_105
timestamp 1607319584
transform 1 0 836 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_359
timestamp 1607319584
transform 1 0 868 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_599
timestamp 1607319584
transform -1 0 924 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1153
timestamp 1607319584
transform -1 0 948 0 -1 3105
box -2 -3 34 103
use AOI22X1  AOI22X1_17
timestamp 1607319584
transform -1 0 988 0 -1 3105
box -2 -3 42 103
use MUX2X1  MUX2X1_271
timestamp 1607319584
transform 1 0 988 0 -1 3105
box -2 -3 50 103
use BUFX4  BUFX4_360
timestamp 1607319584
transform -1 0 956 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_402
timestamp 1607319584
transform 1 0 956 0 1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_125
timestamp 1607319584
transform 1 0 1036 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_1_0
timestamp 1607319584
transform -1 0 1068 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_1_1
timestamp 1607319584
transform -1 0 1076 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_149
timestamp 1607319584
transform -1 0 1100 0 -1 3105
box -2 -3 26 103
use BUFX4  BUFX4_358
timestamp 1607319584
transform 1 0 1100 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_1_0
timestamp 1607319584
transform -1 0 1060 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_1_1
timestamp 1607319584
transform -1 0 1068 0 1 3105
box -2 -3 10 103
use BUFX4  BUFX4_396
timestamp 1607319584
transform -1 0 1100 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_80
timestamp 1607319584
transform 1 0 1100 0 1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_129
timestamp 1607319584
transform -1 0 1180 0 -1 3105
box -2 -3 50 103
use AOI22X1  AOI22X1_77
timestamp 1607319584
transform -1 0 1220 0 -1 3105
box -2 -3 42 103
use OAI21X1  OAI21X1_76
timestamp 1607319584
transform 1 0 1132 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_75
timestamp 1607319584
transform -1 0 1196 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_79
timestamp 1607319584
transform -1 0 1228 0 1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_369
timestamp 1607319584
transform 1 0 1220 0 -1 3105
box -2 -3 50 103
use BUFX4  BUFX4_357
timestamp 1607319584
transform 1 0 1268 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_111
timestamp 1607319584
transform 1 0 1300 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_77
timestamp 1607319584
transform 1 0 1228 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_78
timestamp 1607319584
transform -1 0 1292 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_403
timestamp 1607319584
transform 1 0 1292 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_1022
timestamp 1607319584
transform -1 0 1356 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_957
timestamp 1607319584
transform 1 0 1356 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_86
timestamp 1607319584
transform -1 0 1412 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_457
timestamp 1607319584
transform -1 0 1436 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_732
timestamp 1607319584
transform -1 0 1484 0 1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_68
timestamp 1607319584
transform -1 0 1468 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_150
timestamp 1607319584
transform 1 0 1468 0 -1 3105
box -2 -3 18 103
use INVX1  INVX1_86
timestamp 1607319584
transform 1 0 1484 0 -1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_749
timestamp 1607319584
transform 1 0 1500 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_214
timestamp 1607319584
transform 1 0 1484 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_574
timestamp 1607319584
transform -1 0 1524 0 1 3105
box -2 -3 26 103
use FILL  FILL_30_2_0
timestamp 1607319584
transform 1 0 1596 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_2_1
timestamp 1607319584
transform 1 0 1604 0 -1 3105
box -2 -3 10 103
use AOI21X1  AOI21X1_77
timestamp 1607319584
transform 1 0 1612 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1002
timestamp 1607319584
transform 1 0 1524 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_2_0
timestamp 1607319584
transform -1 0 1564 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_2_1
timestamp 1607319584
transform -1 0 1572 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_436
timestamp 1607319584
transform -1 0 1596 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_95
timestamp 1607319584
transform -1 0 1628 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_97
timestamp 1607319584
transform 1 0 1644 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1085
timestamp 1607319584
transform 1 0 1668 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1130
timestamp 1607319584
transform 1 0 1700 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_316
timestamp 1607319584
transform 1 0 1628 0 1 3105
box -2 -3 50 103
use NAND2X1  NAND2X1_525
timestamp 1607319584
transform -1 0 1700 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1214
timestamp 1607319584
transform -1 0 1732 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_355
timestamp 1607319584
transform 1 0 1732 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_365
timestamp 1607319584
transform 1 0 1764 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_255
timestamp 1607319584
transform -1 0 1844 0 -1 3105
box -2 -3 50 103
use BUFX4  BUFX4_364
timestamp 1607319584
transform 1 0 1732 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_398
timestamp 1607319584
transform -1 0 1860 0 1 3105
box -2 -3 98 103
use MUX2X1  MUX2X1_253
timestamp 1607319584
transform -1 0 1892 0 -1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_1129
timestamp 1607319584
transform -1 0 1924 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_573
timestamp 1607319584
transform 1 0 1860 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_8
timestamp 1607319584
transform 1 0 1884 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_6
timestamp 1607319584
transform -1 0 1940 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_527
timestamp 1607319584
transform -1 0 1948 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_472
timestamp 1607319584
transform -1 0 1964 0 -1 3105
box -2 -3 18 103
use BUFX4  BUFX4_100
timestamp 1607319584
transform -1 0 1996 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_220
timestamp 1607319584
transform 1 0 1996 0 -1 3105
box -2 -3 50 103
use BUFX4  BUFX4_309
timestamp 1607319584
transform -1 0 1972 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_733
timestamp 1607319584
transform 1 0 1972 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_1087
timestamp 1607319584
transform -1 0 2076 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_3_0
timestamp 1607319584
transform -1 0 2084 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_3_1
timestamp 1607319584
transform -1 0 2092 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_1086
timestamp 1607319584
transform -1 0 2124 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_18
timestamp 1607319584
transform -1 0 2148 0 -1 3105
box -2 -3 26 103
use FILL  FILL_31_3_0
timestamp 1607319584
transform 1 0 2068 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_3_1
timestamp 1607319584
transform 1 0 2076 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_526
timestamp 1607319584
transform 1 0 2084 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_87
timestamp 1607319584
transform 1 0 2108 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_298
timestamp 1607319584
transform -1 0 2164 0 -1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_725
timestamp 1607319584
transform -1 0 2260 0 -1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_69
timestamp 1607319584
transform -1 0 2164 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_109
timestamp 1607319584
transform -1 0 2188 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_87
timestamp 1607319584
transform -1 0 2220 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_767
timestamp 1607319584
transform 1 0 2220 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_549
timestamp 1607319584
transform 1 0 2260 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_666
timestamp 1607319584
transform -1 0 2316 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_284
timestamp 1607319584
transform 1 0 2316 0 -1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_111
timestamp 1607319584
transform -1 0 2340 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_428
timestamp 1607319584
transform 1 0 2412 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_555
timestamp 1607319584
transform -1 0 2372 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_171
timestamp 1607319584
transform -1 0 2388 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_739
timestamp 1607319584
transform -1 0 2484 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_363
timestamp 1607319584
transform 1 0 2436 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_289
timestamp 1607319584
transform -1 0 2492 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_105
timestamp 1607319584
transform -1 0 2516 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_959
timestamp 1607319584
transform 1 0 2516 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_303
timestamp 1607319584
transform -1 0 2532 0 1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_86
timestamp 1607319584
transform 1 0 2564 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_79
timestamp 1607319584
transform 1 0 2532 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_389
timestamp 1607319584
transform 1 0 2572 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_99
timestamp 1607319584
transform -1 0 2572 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_85
timestamp 1607319584
transform -1 0 2644 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_4_1
timestamp 1607319584
transform -1 0 2612 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_4_0
timestamp 1607319584
transform -1 0 2604 0 1 3105
box -2 -3 10 103
use FILL  FILL_30_4_1
timestamp 1607319584
transform -1 0 2612 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_4_0
timestamp 1607319584
transform -1 0 2604 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_751
timestamp 1607319584
transform -1 0 2708 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_747
timestamp 1607319584
transform -1 0 2804 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_407
timestamp 1607319584
transform -1 0 2740 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_95
timestamp 1607319584
transform 1 0 2804 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_75
timestamp 1607319584
transform -1 0 2860 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1607319584
transform -1 0 2764 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_82
timestamp 1607319584
transform 1 0 2764 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_81
timestamp 1607319584
transform 1 0 2796 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_405
timestamp 1607319584
transform 1 0 2828 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_98
timestamp 1607319584
transform 1 0 2860 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1607319584
transform 1 0 2892 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_413
timestamp 1607319584
transform 1 0 2924 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_278
timestamp 1607319584
transform 1 0 2924 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_505
timestamp 1607319584
transform -1 0 3044 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_358
timestamp 1607319584
transform -1 0 2964 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_565
timestamp 1607319584
transform 1 0 2964 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1066
timestamp 1607319584
transform 1 0 2988 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1612
timestamp 1607319584
transform 1 0 3020 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_642
timestamp 1607319584
transform 1 0 3044 0 -1 3105
box -2 -3 26 103
use MUX2X1  MUX2X1_205
timestamp 1607319584
transform -1 0 3116 0 -1 3105
box -2 -3 50 103
use FILL  FILL_30_5_0
timestamp 1607319584
transform 1 0 3116 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_5_1
timestamp 1607319584
transform 1 0 3124 0 -1 3105
box -2 -3 10 103
use MUX2X1  MUX2X1_207
timestamp 1607319584
transform 1 0 3132 0 -1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_1613
timestamp 1607319584
transform -1 0 3084 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_5_0
timestamp 1607319584
transform -1 0 3092 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_5_1
timestamp 1607319584
transform -1 0 3100 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_270
timestamp 1607319584
transform -1 0 3196 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1607319584
transform 1 0 3180 0 -1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_850
timestamp 1607319584
transform 1 0 3196 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1624
timestamp 1607319584
transform -1 0 3252 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_323
timestamp 1607319584
transform 1 0 3276 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_1374
timestamp 1607319584
transform 1 0 3292 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_803
timestamp 1607319584
transform 1 0 3324 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_279
timestamp 1607319584
transform 1 0 3252 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_399
timestamp 1607319584
transform -1 0 3444 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_398
timestamp 1607319584
transform 1 0 3348 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_1111
timestamp 1607319584
transform 1 0 3364 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1607319584
transform -1 0 3420 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_5
timestamp 1607319584
transform -1 0 3452 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_9
timestamp 1607319584
transform 1 0 3444 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1065
timestamp 1607319584
transform -1 0 3500 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_7
timestamp 1607319584
transform -1 0 3532 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_10
timestamp 1607319584
transform 1 0 3532 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_504
timestamp 1607319584
transform 1 0 3452 0 1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_397
timestamp 1607319584
transform -1 0 3572 0 1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_290
timestamp 1607319584
transform 1 0 3572 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_269
timestamp 1607319584
transform 1 0 3588 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_69
timestamp 1607319584
transform -1 0 3588 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_364
timestamp 1607319584
transform -1 0 3644 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_6_1
timestamp 1607319584
transform -1 0 3620 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_6_0
timestamp 1607319584
transform -1 0 3612 0 1 3105
box -2 -3 10 103
use INVX1  INVX1_277
timestamp 1607319584
transform -1 0 3636 0 -1 3105
box -2 -3 18 103
use FILL  FILL_30_6_1
timestamp 1607319584
transform -1 0 3620 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_6_0
timestamp 1607319584
transform -1 0 3612 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_389
timestamp 1607319584
transform -1 0 3732 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_301
timestamp 1607319584
transform -1 0 3828 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_285
timestamp 1607319584
transform -1 0 3740 0 1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_634
timestamp 1607319584
transform 1 0 3740 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_374
timestamp 1607319584
transform 1 0 3828 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1614
timestamp 1607319584
transform 1 0 3764 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1615
timestamp 1607319584
transform -1 0 3828 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_271
timestamp 1607319584
transform -1 0 3924 0 1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_298
timestamp 1607319584
transform -1 0 3884 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_99
timestamp 1607319584
transform 1 0 3884 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_324
timestamp 1607319584
transform 1 0 3916 0 -1 3105
box -2 -3 18 103
use MUX2X1  MUX2X1_288
timestamp 1607319584
transform 1 0 3932 0 -1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_1606
timestamp 1607319584
transform 1 0 3924 0 1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_146
timestamp 1607319584
transform -1 0 4028 0 -1 3105
box -2 -3 50 103
use OAI21X1  OAI21X1_987
timestamp 1607319584
transform 1 0 4028 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1607
timestamp 1607319584
transform -1 0 3988 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_267
timestamp 1607319584
transform -1 0 4084 0 1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_420
timestamp 1607319584
transform 1 0 4060 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_804
timestamp 1607319584
transform 1 0 4084 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_7_0
timestamp 1607319584
transform 1 0 4108 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_7_1
timestamp 1607319584
transform 1 0 4116 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_156
timestamp 1607319584
transform 1 0 4124 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_7_0
timestamp 1607319584
transform 1 0 4084 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_7_1
timestamp 1607319584
transform 1 0 4092 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_173
timestamp 1607319584
transform 1 0 4100 0 1 3105
box -2 -3 98 103
use MUX2X1  MUX2X1_243
timestamp 1607319584
transform -1 0 4268 0 -1 3105
box -2 -3 50 103
use AOI21X1  AOI21X1_258
timestamp 1607319584
transform 1 0 4196 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_326
timestamp 1607319584
transform 1 0 4228 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_556
timestamp 1607319584
transform 1 0 4268 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1113
timestamp 1607319584
transform 1 0 4292 0 -1 3105
box -2 -3 34 103
use MUX2X1  MUX2X1_241
timestamp 1607319584
transform 1 0 4324 0 -1 3105
box -2 -3 50 103
use MUX2X1  MUX2X1_195
timestamp 1607319584
transform -1 0 4300 0 1 3105
box -2 -3 50 103
use CLKBUF1  CLKBUF1_12
timestamp 1607319584
transform -1 0 4372 0 1 3105
box -2 -3 74 103
use AOI21X1  AOI21X1_102
timestamp 1607319584
transform 1 0 4372 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_128
timestamp 1607319584
transform -1 0 4428 0 -1 3105
box -2 -3 26 103
use BUFX4  BUFX4_216
timestamp 1607319584
transform 1 0 4428 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_812
timestamp 1607319584
transform 1 0 4372 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_1114
timestamp 1607319584
transform -1 0 4492 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_557
timestamp 1607319584
transform 1 0 4492 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1416
timestamp 1607319584
transform 1 0 4516 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1415
timestamp 1607319584
transform -1 0 4580 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_280
timestamp 1607319584
transform 1 0 4468 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_857
timestamp 1607319584
transform -1 0 4524 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_242
timestamp 1607319584
transform -1 0 4556 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1431
timestamp 1607319584
transform -1 0 4612 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1432
timestamp 1607319584
transform -1 0 4644 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_8_0
timestamp 1607319584
transform -1 0 4652 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1607319584
transform -1 0 4652 0 1 3105
box -2 -3 98 103
use FILL  FILL_30_8_1
timestamp 1607319584
transform -1 0 4660 0 -1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_328
timestamp 1607319584
transform -1 0 4684 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_260
timestamp 1607319584
transform -1 0 4716 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_158
timestamp 1607319584
transform -1 0 4812 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_8_0
timestamp 1607319584
transform 1 0 4652 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_8_1
timestamp 1607319584
transform 1 0 4660 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_248
timestamp 1607319584
transform 1 0 4668 0 1 3105
box -2 -3 26 103
use MUX2X1  MUX2X1_193
timestamp 1607319584
transform 1 0 4692 0 1 3105
box -2 -3 50 103
use NAND2X1  NAND2X1_852
timestamp 1607319584
transform -1 0 4764 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1435
timestamp 1607319584
transform 1 0 4812 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1436
timestamp 1607319584
transform -1 0 4876 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1626
timestamp 1607319584
transform -1 0 4796 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_18
timestamp 1607319584
transform -1 0 4812 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_289
timestamp 1607319584
transform -1 0 4908 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1607319584
transform -1 0 4972 0 -1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_1050
timestamp 1607319584
transform 1 0 4908 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_249
timestamp 1607319584
transform 1 0 4940 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_829
timestamp 1607319584
transform -1 0 5004 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_199
timestamp 1607319584
transform -1 0 5020 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_820
timestamp 1607319584
transform 1 0 5020 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1445
timestamp 1607319584
transform -1 0 5076 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_1452
timestamp 1607319584
transform -1 0 4996 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_164
timestamp 1607319584
transform -1 0 5092 0 1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_816
timestamp 1607319584
transform 1 0 5076 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_1441
timestamp 1607319584
transform -1 0 5132 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_42
timestamp 1607319584
transform -1 0 5148 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_820
timestamp 1607319584
transform -1 0 5180 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1607319584
transform -1 0 5188 0 1 3105
box -2 -3 98 103
use FILL  FILL_31_1
timestamp 1607319584
transform -1 0 5188 0 -1 3105
box -2 -3 10 103
use FILL  FILL_31_2
timestamp 1607319584
transform -1 0 5196 0 -1 3105
box -2 -3 10 103
use FILL  FILL_32_1
timestamp 1607319584
transform 1 0 5188 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_810
timestamp 1607319584
transform -1 0 100 0 -1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_128
timestamp 1607319584
transform -1 0 124 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_778
timestamp 1607319584
transform 1 0 124 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_588
timestamp 1607319584
transform 1 0 220 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_587
timestamp 1607319584
transform -1 0 284 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_109
timestamp 1607319584
transform 1 0 284 0 -1 3305
box -2 -3 18 103
use AOI21X1  AOI21X1_95
timestamp 1607319584
transform -1 0 332 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_897
timestamp 1607319584
transform 1 0 332 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_323
timestamp 1607319584
transform -1 0 388 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_782
timestamp 1607319584
transform 1 0 388 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_783
timestamp 1607319584
transform 1 0 484 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_0_0
timestamp 1607319584
transform 1 0 580 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_0_1
timestamp 1607319584
transform 1 0 588 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_598
timestamp 1607319584
transform 1 0 596 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_597
timestamp 1607319584
transform -1 0 660 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_101
timestamp 1607319584
transform 1 0 660 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_127
timestamp 1607319584
transform -1 0 716 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_592
timestamp 1607319584
transform 1 0 716 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_780
timestamp 1607319584
transform 1 0 748 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_591
timestamp 1607319584
transform -1 0 876 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1154
timestamp 1607319584
transform -1 0 908 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_84
timestamp 1607319584
transform 1 0 908 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_148
timestamp 1607319584
transform -1 0 972 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_458
timestamp 1607319584
transform -1 0 1004 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_1_0
timestamp 1607319584
transform 1 0 1004 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_1_1
timestamp 1607319584
transform 1 0 1012 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_404
timestamp 1607319584
transform 1 0 1020 0 -1 3305
box -2 -3 98 103
use BUFX4  BUFX4_110
timestamp 1607319584
transform -1 0 1148 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_425
timestamp 1607319584
transform -1 0 1180 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_1
timestamp 1607319584
transform -1 0 1204 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_169
timestamp 1607319584
transform 1 0 1204 0 -1 3305
box -2 -3 18 103
use MUX2X1  MUX2X1_174
timestamp 1607319584
transform -1 0 1268 0 -1 3305
box -2 -3 50 103
use BUFX4  BUFX4_249
timestamp 1607319584
transform -1 0 1300 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_120
timestamp 1607319584
transform -1 0 1324 0 -1 3305
box -2 -3 26 103
use MUX2X1  MUX2X1_172
timestamp 1607319584
transform -1 0 1372 0 -1 3305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_414
timestamp 1607319584
transform 1 0 1372 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_100
timestamp 1607319584
transform 1 0 1468 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_99
timestamp 1607319584
transform -1 0 1532 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_2_0
timestamp 1607319584
transform -1 0 1540 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_2_1
timestamp 1607319584
transform -1 0 1548 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_412
timestamp 1607319584
transform -1 0 1644 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_96
timestamp 1607319584
transform -1 0 1676 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_176
timestamp 1607319584
transform -1 0 1708 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_471
timestamp 1607319584
transform 1 0 1708 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1259
timestamp 1607319584
transform 1 0 1724 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_11
timestamp 1607319584
transform 1 0 1756 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_70
timestamp 1607319584
transform -1 0 1812 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_390
timestamp 1607319584
transform 1 0 1812 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_341
timestamp 1607319584
transform 1 0 1908 0 -1 3305
box -2 -3 18 103
use BUFX4  BUFX4_369
timestamp 1607319584
transform -1 0 1956 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_440
timestamp 1607319584
transform -1 0 2052 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_152
timestamp 1607319584
transform 1 0 2052 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_3_0
timestamp 1607319584
transform -1 0 2092 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_3_1
timestamp 1607319584
transform -1 0 2100 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_151
timestamp 1607319584
transform -1 0 2132 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_371
timestamp 1607319584
transform 1 0 2132 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_374
timestamp 1607319584
transform 1 0 2164 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_425
timestamp 1607319584
transform 1 0 2196 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_122
timestamp 1607319584
transform 1 0 2292 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_121
timestamp 1607319584
transform -1 0 2356 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_408
timestamp 1607319584
transform 1 0 2356 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1196
timestamp 1607319584
transform 1 0 2372 0 -1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_302
timestamp 1607319584
transform -1 0 2452 0 -1 3305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_415
timestamp 1607319584
transform 1 0 2452 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_102
timestamp 1607319584
transform 1 0 2548 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_4_0
timestamp 1607319584
transform -1 0 2588 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_4_1
timestamp 1607319584
transform -1 0 2596 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_101
timestamp 1607319584
transform -1 0 2628 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_643
timestamp 1607319584
transform -1 0 2652 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_406
timestamp 1607319584
transform 1 0 2652 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1194
timestamp 1607319584
transform 1 0 2668 0 -1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_301
timestamp 1607319584
transform -1 0 2748 0 -1 3305
box -2 -3 50 103
use INVX1  INVX1_25
timestamp 1607319584
transform 1 0 2748 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1193
timestamp 1607319584
transform -1 0 2796 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_71
timestamp 1607319584
transform 1 0 2796 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1607319584
transform -1 0 2852 0 -1 3305
box -2 -3 26 103
use MUX2X1  MUX2X1_249
timestamp 1607319584
transform -1 0 2900 0 -1 3305
box -2 -3 50 103
use MUX2X1  MUX2X1_247
timestamp 1607319584
transform -1 0 2948 0 -1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_1122
timestamp 1607319584
transform -1 0 2980 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1121
timestamp 1607319584
transform -1 0 3012 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_359
timestamp 1607319584
transform -1 0 3036 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_333
timestamp 1607319584
transform -1 0 3052 0 -1 3305
box -2 -3 18 103
use BUFX4  BUFX4_57
timestamp 1607319584
transform -1 0 3084 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_5_0
timestamp 1607319584
transform 1 0 3084 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_5_1
timestamp 1607319584
transform 1 0 3092 0 -1 3305
box -2 -3 10 103
use AOI21X1  AOI21X1_292
timestamp 1607319584
transform 1 0 3100 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_366
timestamp 1607319584
transform -1 0 3156 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_287
timestamp 1607319584
transform 1 0 3156 0 -1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_635
timestamp 1607319584
transform -1 0 3276 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1607319584
transform 1 0 3276 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1370
timestamp 1607319584
transform -1 0 3404 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_67
timestamp 1607319584
transform 1 0 3404 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1186
timestamp 1607319584
transform 1 0 3420 0 -1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_297
timestamp 1607319584
transform -1 0 3500 0 -1 3305
box -2 -3 50 103
use MUX2X1  MUX2X1_295
timestamp 1607319584
transform -1 0 3548 0 -1 3305
box -2 -3 50 103
use MUX2X1  MUX2X1_336
timestamp 1607319584
transform 1 0 3548 0 -1 3305
box -2 -3 50 103
use NAND2X1  NAND2X1_498
timestamp 1607319584
transform 1 0 3596 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_6_0
timestamp 1607319584
transform -1 0 3628 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_6_1
timestamp 1607319584
transform -1 0 3636 0 -1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_358
timestamp 1607319584
transform -1 0 3660 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_77
timestamp 1607319584
transform 1 0 3660 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1185
timestamp 1607319584
transform -1 0 3708 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_397
timestamp 1607319584
transform -1 0 3724 0 -1 3305
box -2 -3 18 103
use BUFX4  BUFX4_345
timestamp 1607319584
transform 1 0 3724 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1637
timestamp 1607319584
transform 1 0 3756 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1636
timestamp 1607319584
transform 1 0 3788 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_306
timestamp 1607319584
transform 1 0 3820 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_80
timestamp 1607319584
transform 1 0 3916 0 -1 3305
box -2 -3 18 103
use MUX2X1  MUX2X1_56
timestamp 1607319584
transform -1 0 3980 0 -1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_1176
timestamp 1607319584
transform 1 0 3980 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1607319584
transform 1 0 4012 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_7_0
timestamp 1607319584
transform -1 0 4116 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_7_1
timestamp 1607319584
transform -1 0 4124 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_1371
timestamp 1607319584
transform -1 0 4156 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_489
timestamp 1607319584
transform 1 0 4156 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1051
timestamp 1607319584
transform -1 0 4212 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_337
timestamp 1607319584
transform 1 0 4212 0 -1 3305
box -2 -3 26 103
use MUX2X1  MUX2X1_194
timestamp 1607319584
transform 1 0 4236 0 -1 3305
box -2 -3 50 103
use INVX1  INVX1_325
timestamp 1607319584
transform 1 0 4284 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1607319584
transform -1 0 4396 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1453
timestamp 1607319584
transform 1 0 4396 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_828
timestamp 1607319584
transform -1 0 4452 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_263
timestamp 1607319584
transform -1 0 4468 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_165
timestamp 1607319584
transform -1 0 4564 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_69
timestamp 1607319584
transform -1 0 4580 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1411
timestamp 1607319584
transform 1 0 4580 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1412
timestamp 1607319584
transform -1 0 4644 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_8_0
timestamp 1607319584
transform -1 0 4652 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_8_1
timestamp 1607319584
transform -1 0 4660 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1607319584
transform -1 0 4756 0 -1 3305
box -2 -3 98 103
use BUFX4  BUFX4_228
timestamp 1607319584
transform -1 0 4788 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_240
timestamp 1607319584
transform -1 0 4820 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_828
timestamp 1607319584
transform 1 0 4820 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_829
timestamp 1607319584
transform 1 0 4852 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_827
timestamp 1607319584
transform 1 0 4876 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_255
timestamp 1607319584
transform 1 0 4900 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_323
timestamp 1607319584
transform -1 0 4956 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_153
timestamp 1607319584
transform -1 0 5052 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1607319584
transform 1 0 5052 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_134
timestamp 1607319584
transform 1 0 5148 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1443
timestamp 1607319584
transform 1 0 5164 0 -1 3305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_74
timestamp 1607319584
transform 1 0 4 0 1 3305
box -2 -3 74 103
use NOR2X1  NOR2X1_126
timestamp 1607319584
transform 1 0 76 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_100
timestamp 1607319584
transform -1 0 132 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_770
timestamp 1607319584
transform 1 0 132 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_572
timestamp 1607319584
transform 1 0 228 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_571
timestamp 1607319584
transform -1 0 292 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_798
timestamp 1607319584
transform 1 0 292 0 1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_119
timestamp 1607319584
transform -1 0 412 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_773
timestamp 1607319584
transform 1 0 412 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_578
timestamp 1607319584
transform 1 0 508 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_0_0
timestamp 1607319584
transform -1 0 548 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_0_1
timestamp 1607319584
transform -1 0 556 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_577
timestamp 1607319584
transform -1 0 588 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_811
timestamp 1607319584
transform 1 0 588 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_599
timestamp 1607319584
transform 1 0 684 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_600
timestamp 1607319584
transform -1 0 748 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_784
timestamp 1607319584
transform -1 0 844 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_600
timestamp 1607319584
transform -1 0 868 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_764
timestamp 1607319584
transform 1 0 868 0 1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_106
timestamp 1607319584
transform -1 0 988 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_715
timestamp 1607319584
transform 1 0 988 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_1_0
timestamp 1607319584
transform 1 0 1084 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_1_1
timestamp 1607319584
transform 1 0 1092 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_534
timestamp 1607319584
transform 1 0 1100 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_533
timestamp 1607319584
transform 1 0 1132 0 1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_173
timestamp 1607319584
transform 1 0 1164 0 1 3305
box -2 -3 50 103
use NAND2X1  NAND2X1_459
timestamp 1607319584
transform -1 0 1236 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1024
timestamp 1607319584
transform -1 0 1268 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_236
timestamp 1607319584
transform -1 0 1284 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_564
timestamp 1607319584
transform 1 0 1284 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_756
timestamp 1607319584
transform -1 0 1412 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_387
timestamp 1607319584
transform -1 0 1436 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1021
timestamp 1607319584
transform -1 0 1468 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_418
timestamp 1607319584
transform -1 0 1500 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_538
timestamp 1607319584
transform 1 0 1500 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_537
timestamp 1607319584
transform 1 0 1532 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_2_0
timestamp 1607319584
transform 1 0 1564 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_2_1
timestamp 1607319584
transform 1 0 1572 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_717
timestamp 1607319584
transform 1 0 1580 0 1 3305
box -2 -3 98 103
use BUFX4  BUFX4_196
timestamp 1607319584
transform 1 0 1676 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_664
timestamp 1607319584
transform -1 0 1732 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_713
timestamp 1607319584
transform 1 0 1732 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_135
timestamp 1607319584
transform 1 0 1756 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_136
timestamp 1607319584
transform -1 0 1820 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_432
timestamp 1607319584
transform -1 0 1916 0 1 3305
box -2 -3 98 103
use MUX2X1  MUX2X1_308
timestamp 1607319584
transform -1 0 1964 0 1 3305
box -2 -3 50 103
use OAI21X1  OAI21X1_156
timestamp 1607319584
transform 1 0 1964 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_155
timestamp 1607319584
transform -1 0 2028 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1203
timestamp 1607319584
transform 1 0 2028 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_299
timestamp 1607319584
transform -1 0 2076 0 1 3305
box -2 -3 18 103
use FILL  FILL_33_3_0
timestamp 1607319584
transform -1 0 2084 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_3_1
timestamp 1607319584
transform -1 0 2092 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_741
timestamp 1607319584
transform -1 0 2188 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_557
timestamp 1607319584
transform 1 0 2188 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_113
timestamp 1607319584
transform -1 0 2244 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_175
timestamp 1607319584
transform -1 0 2276 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_165
timestamp 1607319584
transform 1 0 2276 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_166
timestamp 1607319584
transform -1 0 2340 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_447
timestamp 1607319584
transform 1 0 2340 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_645
timestamp 1607319584
transform -1 0 2460 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_422
timestamp 1607319584
transform 1 0 2460 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_134
timestamp 1607319584
transform 1 0 2492 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_133
timestamp 1607319584
transform 1 0 2524 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1195
timestamp 1607319584
transform 1 0 2556 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_4_0
timestamp 1607319584
transform 1 0 2588 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_4_1
timestamp 1607319584
transform 1 0 2596 0 1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_644
timestamp 1607319584
transform 1 0 2604 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_431
timestamp 1607319584
transform -1 0 2724 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_268
timestamp 1607319584
transform 1 0 2724 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1609
timestamp 1607319584
transform 1 0 2820 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1608
timestamp 1607319584
transform -1 0 2884 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_427
timestamp 1607319584
transform -1 0 2908 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_993
timestamp 1607319584
transform -1 0 2940 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_566
timestamp 1607319584
transform -1 0 2964 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_334
timestamp 1607319584
transform -1 0 2980 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_278
timestamp 1607319584
transform -1 0 3076 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1623
timestamp 1607319584
transform 1 0 3076 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_5_0
timestamp 1607319584
transform -1 0 3116 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_5_1
timestamp 1607319584
transform -1 0 3124 0 1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_849
timestamp 1607319584
transform -1 0 3148 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_405
timestamp 1607319584
transform -1 0 3164 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_391
timestamp 1607319584
transform -1 0 3260 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1596
timestamp 1607319584
transform 1 0 3260 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1597
timestamp 1607319584
transform -1 0 3324 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_262
timestamp 1607319584
transform -1 0 3420 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_283
timestamp 1607319584
transform -1 0 3516 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_623
timestamp 1607319584
transform -1 0 3540 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1595
timestamp 1607319584
transform 1 0 3540 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1594
timestamp 1607319584
transform 1 0 3572 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_6_0
timestamp 1607319584
transform 1 0 3604 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_6_1
timestamp 1607319584
transform 1 0 3612 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_261
timestamp 1607319584
transform 1 0 3620 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_805
timestamp 1607319584
transform 1 0 3716 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_348
timestamp 1607319584
transform 1 0 3748 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1598
timestamp 1607319584
transform 1 0 3780 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1599
timestamp 1607319584
transform -1 0 3844 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_263
timestamp 1607319584
transform -1 0 3940 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_868
timestamp 1607319584
transform -1 0 3972 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_166
timestamp 1607319584
transform 1 0 3972 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_624
timestamp 1607319584
transform -1 0 4028 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_420
timestamp 1607319584
transform 1 0 4028 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_217
timestamp 1607319584
transform -1 0 4084 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_457
timestamp 1607319584
transform 1 0 4084 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_7_0
timestamp 1607319584
transform 1 0 4116 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_7_1
timestamp 1607319584
transform 1 0 4124 0 1 3305
box -2 -3 10 103
use INVX1  INVX1_131
timestamp 1607319584
transform 1 0 4132 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_1602
timestamp 1607319584
transform 1 0 4148 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1603
timestamp 1607319584
transform -1 0 4212 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_244
timestamp 1607319584
transform -1 0 4236 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_267
timestamp 1607319584
transform -1 0 4268 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_265
timestamp 1607319584
transform 1 0 4268 0 1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_332
timestamp 1607319584
transform -1 0 4388 0 1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_322
timestamp 1607319584
transform -1 0 4412 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1420
timestamp 1607319584
transform -1 0 4444 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1607319584
transform -1 0 4540 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_1427
timestamp 1607319584
transform -1 0 4572 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1428
timestamp 1607319584
transform -1 0 4604 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1115
timestamp 1607319584
transform 1 0 4604 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_8_0
timestamp 1607319584
transform -1 0 4644 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_8_1
timestamp 1607319584
transform -1 0 4652 0 1 3305
box -2 -3 10 103
use BUFX4  BUFX4_221
timestamp 1607319584
transform -1 0 4684 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_186
timestamp 1607319584
transform -1 0 4716 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_250
timestamp 1607319584
transform -1 0 4748 0 1 3305
box -2 -3 34 103
use MUX2X1  MUX2X1_97
timestamp 1607319584
transform 1 0 4748 0 1 3305
box -2 -3 50 103
use BUFX4  BUFX4_245
timestamp 1607319584
transform -1 0 4828 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_247
timestamp 1607319584
transform 1 0 4828 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_244
timestamp 1607319584
transform 1 0 4852 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1425
timestamp 1607319584
transform 1 0 4884 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_488
timestamp 1607319584
transform 1 0 4916 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_1426
timestamp 1607319584
transform -1 0 4972 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1454
timestamp 1607319584
transform -1 0 5004 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1607319584
transform -1 0 5100 0 1 3305
box -2 -3 98 103
use INVX1  INVX1_262
timestamp 1607319584
transform -1 0 5116 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_922
timestamp 1607319584
transform -1 0 5148 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_822
timestamp 1607319584
transform 1 0 5148 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_327
timestamp 1607319584
transform -1 0 5188 0 1 3305
box -2 -3 18 103
use FILL  FILL_34_1
timestamp 1607319584
transform 1 0 5188 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_772
timestamp 1607319584
transform -1 0 100 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_576
timestamp 1607319584
transform -1 0 132 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_575
timestamp 1607319584
transform -1 0 164 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_594
timestamp 1607319584
transform 1 0 164 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_593
timestamp 1607319584
transform -1 0 228 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_237
timestamp 1607319584
transform 1 0 228 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_530
timestamp 1607319584
transform -1 0 268 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_787
timestamp 1607319584
transform 1 0 268 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_602
timestamp 1607319584
transform 1 0 364 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_129
timestamp 1607319584
transform -1 0 420 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1089
timestamp 1607319584
transform -1 0 452 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_301
timestamp 1607319584
transform -1 0 468 0 -1 3505
box -2 -3 18 103
use MUX2X1  MUX2X1_223
timestamp 1607319584
transform -1 0 516 0 -1 3505
box -2 -3 50 103
use FILL  FILL_34_0_0
timestamp 1607319584
transform -1 0 524 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_0_1
timestamp 1607319584
transform -1 0 532 0 -1 3505
box -2 -3 10 103
use MUX2X1  MUX2X1_127
timestamp 1607319584
transform -1 0 580 0 -1 3505
box -2 -3 50 103
use INVX1  INVX1_3
timestamp 1607319584
transform 1 0 580 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_126
timestamp 1607319584
transform -1 0 620 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_127
timestamp 1607319584
transform -1 0 644 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1025
timestamp 1607319584
transform 1 0 644 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_737
timestamp 1607319584
transform 1 0 676 0 -1 3505
box -2 -3 26 103
use MUX2X1  MUX2X1_175
timestamp 1607319584
transform -1 0 748 0 -1 3505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_748
timestamp 1607319584
transform 1 0 748 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_461
timestamp 1607319584
transform -1 0 868 0 -1 3505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_29
timestamp 1607319584
transform 1 0 868 0 -1 3505
box -2 -3 74 103
use NAND2X1  NAND2X1_458
timestamp 1607319584
transform -1 0 964 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1023
timestamp 1607319584
transform -1 0 996 0 -1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_367
timestamp 1607319584
transform -1 0 1044 0 -1 3505
box -2 -3 50 103
use FILL  FILL_34_1_0
timestamp 1607319584
transform 1 0 1044 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_1_1
timestamp 1607319584
transform 1 0 1052 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_542
timestamp 1607319584
transform 1 0 1060 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_541
timestamp 1607319584
transform -1 0 1124 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_429
timestamp 1607319584
transform 1 0 1124 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_735
timestamp 1607319584
transform 1 0 1156 0 -1 3505
box -2 -3 98 103
use AOI21X1  AOI21X1_71
timestamp 1607319584
transform 1 0 1252 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_89
timestamp 1607319584
transform 1 0 1284 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_893
timestamp 1607319584
transform 1 0 1308 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_92
timestamp 1607319584
transform 1 0 1340 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_81
timestamp 1607319584
transform -1 0 1388 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_663
timestamp 1607319584
transform -1 0 1412 0 -1 3505
box -2 -3 26 103
use BUFX4  BUFX4_295
timestamp 1607319584
transform 1 0 1412 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_82
timestamp 1607319584
transform 1 0 1444 0 -1 3505
box -2 -3 26 103
use BUFX4  BUFX4_267
timestamp 1607319584
transform -1 0 1500 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_187
timestamp 1607319584
transform 1 0 1500 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_181
timestamp 1607319584
transform -1 0 1564 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_2_0
timestamp 1607319584
transform -1 0 1572 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_2_1
timestamp 1607319584
transform -1 0 1580 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1213
timestamp 1607319584
transform -1 0 1612 0 -1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_254
timestamp 1607319584
transform 1 0 1612 0 -1 3505
box -2 -3 50 103
use OAI21X1  OAI21X1_1132
timestamp 1607319584
transform -1 0 1692 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_344
timestamp 1607319584
transform -1 0 1708 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_1204
timestamp 1607319584
transform -1 0 1740 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_442
timestamp 1607319584
transform 1 0 1740 0 -1 3505
box -2 -3 98 103
use MUX2X1  MUX2X1_309
timestamp 1607319584
transform 1 0 1836 0 -1 3505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_438
timestamp 1607319584
transform -1 0 1980 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_300
timestamp 1607319584
transform 1 0 1980 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_148
timestamp 1607319584
transform 1 0 2004 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_147
timestamp 1607319584
transform -1 0 2068 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_3_0
timestamp 1607319584
transform -1 0 2076 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_3_1
timestamp 1607319584
transform -1 0 2084 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_876
timestamp 1607319584
transform -1 0 2116 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_88
timestamp 1607319584
transform -1 0 2132 0 -1 3505
box -2 -3 18 103
use MUX2X1  MUX2X1_62
timestamp 1607319584
transform -1 0 2180 0 -1 3505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_439
timestamp 1607319584
transform 1 0 2180 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_150
timestamp 1607319584
transform 1 0 2276 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1607319584
transform -1 0 2340 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_423
timestamp 1607319584
transform -1 0 2436 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_118
timestamp 1607319584
transform 1 0 2436 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_117
timestamp 1607319584
transform -1 0 2500 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_179
timestamp 1607319584
transform 1 0 2500 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_407
timestamp 1607319584
transform 1 0 2532 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_117
timestamp 1607319584
transform -1 0 2572 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_4_0
timestamp 1607319584
transform -1 0 2580 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_4_1
timestamp 1607319584
transform -1 0 2588 0 -1 3505
box -2 -3 10 103
use BUFX4  BUFX4_173
timestamp 1607319584
transform -1 0 2620 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_137
timestamp 1607319584
transform 1 0 2620 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_138
timestamp 1607319584
transform -1 0 2684 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_433
timestamp 1607319584
transform 1 0 2684 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_286
timestamp 1607319584
transform 1 0 2780 0 -1 3505
box -2 -3 98 103
use AOI21X1  AOI21X1_291
timestamp 1607319584
transform 1 0 2876 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_365
timestamp 1607319584
transform 1 0 2908 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_205
timestamp 1607319584
transform -1 0 2948 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_305
timestamp 1607319584
transform 1 0 2948 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1634
timestamp 1607319584
transform 1 0 3044 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1635
timestamp 1607319584
transform -1 0 3108 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_5_0
timestamp 1607319584
transform -1 0 3116 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_5_1
timestamp 1607319584
transform -1 0 3124 0 -1 3505
box -2 -3 10 103
use BUFX4  BUFX4_346
timestamp 1607319584
transform -1 0 3156 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_359
timestamp 1607319584
transform 1 0 3156 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_930
timestamp 1607319584
transform -1 0 3212 0 -1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_103
timestamp 1607319584
transform -1 0 3260 0 -1 3505
box -2 -3 50 103
use MUX2X1  MUX2X1_105
timestamp 1607319584
transform 1 0 3260 0 -1 3505
box -2 -3 50 103
use MUX2X1  MUX2X1_200
timestamp 1607319584
transform -1 0 3356 0 -1 3505
box -2 -3 50 103
use NOR2X1  NOR2X1_362
timestamp 1607319584
transform -1 0 3380 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_929
timestamp 1607319584
transform -1 0 3412 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_141
timestamp 1607319584
transform -1 0 3428 0 -1 3505
box -2 -3 18 103
use NOR2X1  NOR2X1_309
timestamp 1607319584
transform -1 0 3452 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1059
timestamp 1607319584
transform 1 0 3452 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_257
timestamp 1607319584
transform 1 0 3484 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_809
timestamp 1607319584
transform 1 0 3580 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_6_0
timestamp 1607319584
transform -1 0 3612 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_6_1
timestamp 1607319584
transform -1 0 3620 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1376
timestamp 1607319584
transform -1 0 3652 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_451
timestamp 1607319584
transform -1 0 3668 0 -1 3505
box -2 -3 18 103
use INVX1  INVX1_20
timestamp 1607319584
transform 1 0 3668 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1607319584
transform -1 0 3780 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1239
timestamp 1607319584
transform 1 0 3780 0 -1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_335
timestamp 1607319584
transform 1 0 3812 0 -1 3505
box -2 -3 50 103
use MUX2X1  MUX2X1_152
timestamp 1607319584
transform -1 0 3908 0 -1 3505
box -2 -3 50 103
use OAI21X1  OAI21X1_1240
timestamp 1607319584
transform 1 0 3908 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1387
timestamp 1607319584
transform 1 0 3940 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1607319584
transform -1 0 4068 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1405
timestamp 1607319584
transform -1 0 4100 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1406
timestamp 1607319584
transform -1 0 4132 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_7_0
timestamp 1607319584
transform 1 0 4132 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_7_1
timestamp 1607319584
transform 1 0 4140 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1403
timestamp 1607319584
transform 1 0 4148 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1404
timestamp 1607319584
transform -1 0 4212 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1607319584
transform -1 0 4308 0 -1 3505
box -2 -3 98 103
use MUX2X1  MUX2X1_242
timestamp 1607319584
transform 1 0 4308 0 -1 3505
box -2 -3 50 103
use BUFX4  BUFX4_389
timestamp 1607319584
transform 1 0 4356 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1419
timestamp 1607319584
transform 1 0 4388 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_867
timestamp 1607319584
transform -1 0 4452 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_291
timestamp 1607319584
transform 1 0 4452 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1607319584
transform 1 0 4476 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_175
timestamp 1607319584
transform 1 0 4572 0 -1 3505
box -2 -3 98 103
use FILL  FILL_34_8_0
timestamp 1607319584
transform -1 0 4676 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_8_1
timestamp 1607319584
transform -1 0 4684 0 -1 3505
box -2 -3 10 103
use AOI21X1  AOI21X1_269
timestamp 1607319584
transform -1 0 4716 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_823
timestamp 1607319584
transform 1 0 4716 0 -1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_295
timestamp 1607319584
transform 1 0 4740 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_371
timestamp 1607319584
transform -1 0 4796 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_298
timestamp 1607319584
transform -1 0 4892 0 -1 3505
box -2 -3 98 103
use AOI21X1  AOI21X1_259
timestamp 1607319584
transform 1 0 4892 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_327
timestamp 1607319584
transform -1 0 4948 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_157
timestamp 1607319584
transform -1 0 5044 0 -1 3505
box -2 -3 98 103
use INVX1  INVX1_41
timestamp 1607319584
transform -1 0 5060 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_159
timestamp 1607319584
transform 1 0 5060 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1447
timestamp 1607319584
transform 1 0 5156 0 -1 3505
box -2 -3 34 103
use FILL  FILL_35_1
timestamp 1607319584
transform -1 0 5196 0 -1 3505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_62
timestamp 1607319584
transform 1 0 4 0 1 3505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_781
timestamp 1607319584
transform 1 0 76 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_779
timestamp 1607319584
transform 1 0 172 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_590
timestamp 1607319584
transform 1 0 268 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_589
timestamp 1607319584
transform -1 0 332 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_392
timestamp 1607319584
transform -1 0 356 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_174
timestamp 1607319584
transform 1 0 356 0 1 3505
box -2 -3 18 103
use INVX1  INVX1_173
timestamp 1607319584
transform 1 0 372 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_961
timestamp 1607319584
transform 1 0 388 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_962
timestamp 1607319584
transform 1 0 420 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_431
timestamp 1607319584
transform 1 0 452 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_583
timestamp 1607319584
transform 1 0 484 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_427
timestamp 1607319584
transform -1 0 548 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_0_0
timestamp 1607319584
transform 1 0 548 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_0_1
timestamp 1607319584
transform 1 0 556 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_132
timestamp 1607319584
transform 1 0 564 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_605
timestamp 1607319584
transform -1 0 620 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_428
timestamp 1607319584
transform -1 0 652 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_493
timestamp 1607319584
transform 1 0 652 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_1281
timestamp 1607319584
transform 1 0 668 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_740
timestamp 1607319584
transform 1 0 700 0 1 3505
box -2 -3 98 103
use AOI21X1  AOI21X1_76
timestamp 1607319584
transform 1 0 796 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_96
timestamp 1607319584
transform -1 0 852 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_235
timestamp 1607319584
transform 1 0 852 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_556
timestamp 1607319584
transform 1 0 868 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_112
timestamp 1607319584
transform -1 0 924 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_108
timestamp 1607319584
transform -1 0 948 0 1 3505
box -2 -3 26 103
use BUFX4  BUFX4_430
timestamp 1607319584
transform 1 0 948 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1607319584
transform -1 0 1012 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_1_0
timestamp 1607319584
transform 1 0 1012 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_1_1
timestamp 1607319584
transform 1 0 1020 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_719
timestamp 1607319584
transform 1 0 1028 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_532
timestamp 1607319584
transform 1 0 1124 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_714
timestamp 1607319584
transform 1 0 1156 0 1 3505
box -2 -3 98 103
use BUFX4  BUFX4_127
timestamp 1607319584
transform 1 0 1252 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_318
timestamp 1607319584
transform -1 0 1308 0 1 3505
box -2 -3 26 103
use BUFX4  BUFX4_207
timestamp 1607319584
transform 1 0 1308 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_252
timestamp 1607319584
transform -1 0 1372 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_192
timestamp 1607319584
transform 1 0 1372 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_456
timestamp 1607319584
transform -1 0 1428 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_115
timestamp 1607319584
transform 1 0 1428 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_116
timestamp 1607319584
transform -1 0 1492 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_422
timestamp 1607319584
transform -1 0 1588 0 1 3505
box -2 -3 98 103
use FILL  FILL_35_2_0
timestamp 1607319584
transform 1 0 1588 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_2_1
timestamp 1607319584
transform 1 0 1596 0 1 3505
box -2 -3 10 103
use INVX1  INVX1_343
timestamp 1607319584
transform 1 0 1604 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_1131
timestamp 1607319584
transform -1 0 1652 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_178
timestamp 1607319584
transform -1 0 1684 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_654
timestamp 1607319584
transform 1 0 1684 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_424
timestamp 1607319584
transform -1 0 1804 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_120
timestamp 1607319584
transform 1 0 1804 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_119
timestamp 1607319584
transform -1 0 1868 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_418
timestamp 1607319584
transform 1 0 1868 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_108
timestamp 1607319584
transform 1 0 1964 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_107
timestamp 1607319584
transform -1 0 2028 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_87
timestamp 1607319584
transform 1 0 2028 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_875
timestamp 1607319584
transform 1 0 2044 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_3_0
timestamp 1607319584
transform 1 0 2076 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_3_1
timestamp 1607319584
transform 1 0 2084 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_299
timestamp 1607319584
transform 1 0 2092 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_123
timestamp 1607319584
transform -1 0 2148 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1607319584
transform -1 0 2180 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_426
timestamp 1607319584
transform -1 0 2276 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_280
timestamp 1607319584
transform 1 0 2276 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_851
timestamp 1607319584
transform 1 0 2372 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1625
timestamp 1607319584
transform -1 0 2428 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_462
timestamp 1607319584
transform 1 0 2428 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_1250
timestamp 1607319584
transform 1 0 2444 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_704
timestamp 1607319584
transform 1 0 2476 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_288
timestamp 1607319584
transform -1 0 2596 0 1 3505
box -2 -3 98 103
use FILL  FILL_35_4_0
timestamp 1607319584
transform 1 0 2596 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_4_1
timestamp 1607319584
transform 1 0 2604 0 1 3505
box -2 -3 10 103
use AOI21X1  AOI21X1_293
timestamp 1607319584
transform 1 0 2612 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_367
timestamp 1607319584
transform 1 0 2644 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_114
timestamp 1607319584
transform 1 0 2668 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_113
timestamp 1607319584
transform 1 0 2700 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_421
timestamp 1607319584
transform 1 0 2732 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_130
timestamp 1607319584
transform 1 0 2828 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_129
timestamp 1607319584
transform 1 0 2860 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_429
timestamp 1607319584
transform 1 0 2892 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_279
timestamp 1607319584
transform 1 0 2988 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_506
timestamp 1607319584
transform -1 0 3028 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1067
timestamp 1607319584
transform 1 0 3028 0 1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_206
timestamp 1607319584
transform 1 0 3060 0 1 3505
box -2 -3 50 103
use FILL  FILL_35_5_0
timestamp 1607319584
transform 1 0 3108 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_5_1
timestamp 1607319584
transform 1 0 3116 0 1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1592
timestamp 1607319584
transform 1 0 3124 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_260
timestamp 1607319584
transform -1 0 3252 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_142
timestamp 1607319584
transform 1 0 3252 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_1593
timestamp 1607319584
transform -1 0 3300 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_280
timestamp 1607319584
transform -1 0 3332 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_80
timestamp 1607319584
transform 1 0 3332 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_288
timestamp 1607319584
transform -1 0 3396 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_554
timestamp 1607319584
transform -1 0 3420 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1620
timestamp 1607319584
transform 1 0 3420 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_846
timestamp 1607319584
transform -1 0 3476 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_856
timestamp 1607319584
transform 1 0 3476 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1630
timestamp 1607319584
transform -1 0 3532 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_271
timestamp 1607319584
transform -1 0 3548 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_293
timestamp 1607319584
transform -1 0 3644 0 1 3505
box -2 -3 98 103
use FILL  FILL_35_6_0
timestamp 1607319584
transform 1 0 3644 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_6_1
timestamp 1607319584
transform 1 0 3652 0 1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_1587
timestamp 1607319584
transform 1 0 3660 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1586
timestamp 1607319584
transform -1 0 3724 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_347
timestamp 1607319584
transform -1 0 3756 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_692
timestamp 1607319584
transform 1 0 3756 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_195
timestamp 1607319584
transform -1 0 3796 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1607319584
transform -1 0 3892 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_1372
timestamp 1607319584
transform 1 0 3892 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1373
timestamp 1607319584
transform -1 0 3956 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_259
timestamp 1607319584
transform -1 0 3972 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_693
timestamp 1607319584
transform -1 0 3996 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1607319584
transform -1 0 4092 0 1 3505
box -2 -3 98 103
use BUFX4  BUFX4_466
timestamp 1607319584
transform 1 0 4092 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_7_0
timestamp 1607319584
transform 1 0 4124 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_7_1
timestamp 1607319584
transform 1 0 4132 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_802
timestamp 1607319584
transform 1 0 4140 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1369
timestamp 1607319584
transform -1 0 4196 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_825
timestamp 1607319584
transform 1 0 4196 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1607319584
transform -1 0 4244 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1607319584
transform -1 0 4340 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_831
timestamp 1607319584
transform 1 0 4340 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1456
timestamp 1607319584
transform -1 0 4396 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_455
timestamp 1607319584
transform -1 0 4412 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_168
timestamp 1607319584
transform -1 0 4508 0 1 3505
box -2 -3 98 103
use NOR2X1  NOR2X1_321
timestamp 1607319584
transform -1 0 4532 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1417
timestamp 1607319584
transform 1 0 4532 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1418
timestamp 1607319584
transform -1 0 4596 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_261
timestamp 1607319584
transform 1 0 4596 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_1049
timestamp 1607319584
transform 1 0 4612 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_8_0
timestamp 1607319584
transform 1 0 4644 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_8_1
timestamp 1607319584
transform 1 0 4652 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_627
timestamp 1607319584
transform 1 0 4660 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_339
timestamp 1607319584
transform 1 0 4684 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1179
timestamp 1607319584
transform -1 0 4740 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1448
timestamp 1607319584
transform -1 0 4772 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_454
timestamp 1607319584
transform -1 0 4788 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_152
timestamp 1607319584
transform -1 0 4884 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_830
timestamp 1607319584
transform 1 0 4884 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_1455
timestamp 1607319584
transform -1 0 4940 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_391
timestamp 1607319584
transform -1 0 4956 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_167
timestamp 1607319584
transform -1 0 5052 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_350
timestamp 1607319584
transform -1 0 5076 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_261
timestamp 1607319584
transform 1 0 5076 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_329
timestamp 1607319584
transform -1 0 5132 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_390
timestamp 1607319584
transform -1 0 5148 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_818
timestamp 1607319584
transform -1 0 5172 0 1 3505
box -2 -3 26 103
use FILL  FILL_36_1
timestamp 1607319584
transform 1 0 5172 0 1 3505
box -2 -3 10 103
use FILL  FILL_36_2
timestamp 1607319584
transform 1 0 5180 0 1 3505
box -2 -3 10 103
use FILL  FILL_36_3
timestamp 1607319584
transform 1 0 5188 0 1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_116
timestamp 1607319584
transform 1 0 4 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_92
timestamp 1607319584
transform -1 0 60 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_771
timestamp 1607319584
transform 1 0 60 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_574
timestamp 1607319584
transform 1 0 156 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_573
timestamp 1607319584
transform -1 0 220 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_93
timestamp 1607319584
transform 1 0 220 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_117
timestamp 1607319584
transform -1 0 276 0 -1 3705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_26
timestamp 1607319584
transform 1 0 276 0 -1 3705
box -2 -3 74 103
use NOR2X1  NOR2X1_121
timestamp 1607319584
transform 1 0 348 0 -1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_393
timestamp 1607319584
transform -1 0 396 0 -1 3705
box -2 -3 26 103
use MUX2X1  MUX2X1_372
timestamp 1607319584
transform -1 0 444 0 -1 3705
box -2 -3 50 103
use BUFX4  BUFX4_298
timestamp 1607319584
transform -1 0 476 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_584
timestamp 1607319584
transform 1 0 476 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_0_0
timestamp 1607319584
transform 1 0 508 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_0_1
timestamp 1607319584
transform 1 0 516 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_790
timestamp 1607319584
transform 1 0 524 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_366
timestamp 1607319584
transform 1 0 620 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_1282
timestamp 1607319584
transform 1 0 636 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_462
timestamp 1607319584
transform -1 0 692 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1026
timestamp 1607319584
transform -1 0 724 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_728
timestamp 1607319584
transform 1 0 724 0 -1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_96
timestamp 1607319584
transform -1 0 852 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_490
timestamp 1607319584
transform 1 0 852 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_552
timestamp 1607319584
transform 1 0 868 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_84
timestamp 1607319584
transform -1 0 948 0 -1 3705
box -2 -3 50 103
use MUX2X1  MUX2X1_82
timestamp 1607319584
transform -1 0 996 0 -1 3705
box -2 -3 50 103
use BUFX4  BUFX4_372
timestamp 1607319584
transform -1 0 1028 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_91
timestamp 1607319584
transform -1 0 1052 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_1_0
timestamp 1607319584
transform -1 0 1060 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_1_1
timestamp 1607319584
transform -1 0 1068 0 -1 3705
box -2 -3 10 103
use BUFX4  BUFX4_296
timestamp 1607319584
transform -1 0 1100 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_965
timestamp 1607319584
transform 1 0 1100 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_531
timestamp 1607319584
transform -1 0 1164 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_535
timestamp 1607319584
transform 1 0 1164 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_536
timestamp 1607319584
transform -1 0 1228 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_716
timestamp 1607319584
transform 1 0 1228 0 -1 3705
box -2 -3 98 103
use BUFX4  BUFX4_379
timestamp 1607319584
transform -1 0 1356 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_428
timestamp 1607319584
transform 1 0 1356 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_128
timestamp 1607319584
transform 1 0 1452 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1218
timestamp 1607319584
transform -1 0 1516 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_131
timestamp 1607319584
transform 1 0 1516 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_2_0
timestamp 1607319584
transform -1 0 1556 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_2_1
timestamp 1607319584
transform -1 0 1564 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_132
timestamp 1607319584
transform -1 0 1596 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_575
timestamp 1607319584
transform 1 0 1596 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_430
timestamp 1607319584
transform -1 0 1716 0 -1 3705
box -2 -3 98 103
use BUFX4  BUFX4_150
timestamp 1607319584
transform -1 0 1748 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_307
timestamp 1607319584
transform 1 0 1748 0 -1 3705
box -2 -3 50 103
use MUX2X1  MUX2X1_130
timestamp 1607319584
transform -1 0 1844 0 -1 3705
box -2 -3 50 103
use MUX2X1  MUX2X1_132
timestamp 1607319584
transform 1 0 1844 0 -1 3705
box -2 -3 50 103
use MUX2X1  MUX2X1_40
timestamp 1607319584
transform 1 0 1892 0 -1 3705
box -2 -3 50 103
use MUX2X1  MUX2X1_42
timestamp 1607319584
transform 1 0 1940 0 -1 3705
box -2 -3 50 103
use OAI21X1  OAI21X1_846
timestamp 1607319584
transform -1 0 2020 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_58
timestamp 1607319584
transform -1 0 2036 0 -1 3705
box -2 -3 18 103
use FILL  FILL_36_3_0
timestamp 1607319584
transform -1 0 2044 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_3_1
timestamp 1607319584
transform -1 0 2052 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_721
timestamp 1607319584
transform -1 0 2148 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_545
timestamp 1607319584
transform 1 0 2148 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_101
timestamp 1607319584
transform -1 0 2204 0 -1 3705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_77
timestamp 1607319584
transform -1 0 2276 0 -1 3705
box -2 -3 74 103
use MUX2X1  MUX2X1_345
timestamp 1607319584
transform -1 0 2324 0 -1 3705
box -2 -3 50 103
use MUX2X1  MUX2X1_343
timestamp 1607319584
transform -1 0 2372 0 -1 3705
box -2 -3 50 103
use OAI21X1  OAI21X1_139
timestamp 1607319584
transform 1 0 2372 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_753
timestamp 1607319584
transform 1 0 2404 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_60
timestamp 1607319584
transform 1 0 2500 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_561
timestamp 1607319584
transform -1 0 2548 0 -1 3705
box -2 -3 34 103
use INVX4  INVX4_3
timestamp 1607319584
transform -1 0 2572 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_4_0
timestamp 1607319584
transform -1 0 2580 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_4_1
timestamp 1607319584
transform -1 0 2588 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1249
timestamp 1607319584
transform -1 0 2620 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_394
timestamp 1607319584
transform -1 0 2652 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_461
timestamp 1607319584
transform -1 0 2668 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_264
timestamp 1607319584
transform -1 0 2764 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_1600
timestamp 1607319584
transform -1 0 2796 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1601
timestamp 1607319584
transform -1 0 2828 0 -1 3705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_48
timestamp 1607319584
transform -1 0 2900 0 -1 3705
box -2 -3 74 103
use OAI21X1  OAI21X1_1642
timestamp 1607319584
transform 1 0 2900 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1643
timestamp 1607319584
transform -1 0 2964 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_309
timestamp 1607319584
transform 1 0 2964 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_272
timestamp 1607319584
transform 1 0 3060 0 -1 3705
box -2 -3 18 103
use AOI21X1  AOI21X1_253
timestamp 1607319584
transform 1 0 3076 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_5_0
timestamp 1607319584
transform -1 0 3116 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_5_1
timestamp 1607319584
transform -1 0 3124 0 -1 3705
box -2 -3 10 103
use NOR2X1  NOR2X1_318
timestamp 1607319584
transform -1 0 3148 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_275
timestamp 1607319584
transform 1 0 3148 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_1060
timestamp 1607319584
transform 1 0 3244 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_499
timestamp 1607319584
transform 1 0 3276 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1607319584
transform 1 0 3300 0 -1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_252
timestamp 1607319584
transform 1 0 3396 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_317
timestamp 1607319584
transform 1 0 3428 0 -1 3705
box -2 -3 26 103
use MUX2X1  MUX2X1_104
timestamp 1607319584
transform 1 0 3452 0 -1 3705
box -2 -3 50 103
use OAI21X1  OAI21X1_1591
timestamp 1607319584
transform 1 0 3500 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1590
timestamp 1607319584
transform -1 0 3564 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_369
timestamp 1607319584
transform 1 0 3564 0 -1 3705
box -2 -3 26 103
use BUFX4  BUFX4_373
timestamp 1607319584
transform 1 0 3588 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_6_0
timestamp 1607319584
transform 1 0 3620 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_6_1
timestamp 1607319584
transform 1 0 3628 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1658
timestamp 1607319584
transform 1 0 3636 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1659
timestamp 1607319584
transform -1 0 3700 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_317
timestamp 1607319584
transform -1 0 3796 0 -1 3705
box -2 -3 98 103
use NOR2X1  NOR2X1_319
timestamp 1607319584
transform 1 0 3796 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_254
timestamp 1607319584
transform -1 0 3852 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_399
timestamp 1607319584
transform -1 0 3884 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_279
timestamp 1607319584
transform 1 0 3884 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_311
timestamp 1607319584
transform 1 0 3916 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1408
timestamp 1607319584
transform 1 0 3940 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1407
timestamp 1607319584
transform -1 0 4004 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_286
timestamp 1607319584
transform 1 0 4004 0 -1 3705
box -2 -3 50 103
use OAI21X1  OAI21X1_1388
timestamp 1607319584
transform -1 0 4084 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_7_0
timestamp 1607319584
transform -1 0 4092 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_7_1
timestamp 1607319584
transform -1 0 4100 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1607319584
transform -1 0 4196 0 -1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_243
timestamp 1607319584
transform 1 0 4196 0 -1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_312
timestamp 1607319584
transform 1 0 4220 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_247
timestamp 1607319584
transform -1 0 4276 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1607319584
transform -1 0 4372 0 -1 3705
box -2 -3 98 103
use BUFX4  BUFX4_397
timestamp 1607319584
transform 1 0 4372 0 -1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_339
timestamp 1607319584
transform 1 0 4404 0 -1 3705
box -2 -3 50 103
use NAND2X1  NAND2X1_853
timestamp 1607319584
transform 1 0 4452 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1627
timestamp 1607319584
transform -1 0 4508 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_79
timestamp 1607319584
transform -1 0 4524 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_290
timestamp 1607319584
transform -1 0 4620 0 -1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_558
timestamp 1607319584
transform 1 0 4620 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_8_0
timestamp 1607319584
transform 1 0 4644 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_8_1
timestamp 1607319584
transform 1 0 4652 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1242
timestamp 1607319584
transform 1 0 4660 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_695
timestamp 1607319584
transform -1 0 4716 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_174
timestamp 1607319584
transform -1 0 4812 0 -1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_349
timestamp 1607319584
transform 1 0 4812 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_921
timestamp 1607319584
transform -1 0 4868 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_330
timestamp 1607319584
transform -1 0 4892 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_262
timestamp 1607319584
transform -1 0 4924 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_160
timestamp 1607319584
transform -1 0 5020 0 -1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_257
timestamp 1607319584
transform 1 0 5020 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_325
timestamp 1607319584
transform 1 0 5052 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1178
timestamp 1607319584
transform 1 0 5076 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_626
timestamp 1607319584
transform 1 0 5108 0 -1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_340
timestamp 1607319584
transform 1 0 5132 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_270
timestamp 1607319584
transform -1 0 5188 0 -1 3705
box -2 -3 34 103
use FILL  FILL_37_1
timestamp 1607319584
transform -1 0 5196 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_795
timestamp 1607319584
transform -1 0 100 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_788
timestamp 1607319584
transform 1 0 100 0 1 3705
box -2 -3 98 103
use INVX1  INVX1_238
timestamp 1607319584
transform 1 0 196 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_796
timestamp 1607319584
transform 1 0 212 0 1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_97
timestamp 1607319584
transform 1 0 308 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_531
timestamp 1607319584
transform -1 0 364 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1090
timestamp 1607319584
transform -1 0 396 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_603
timestamp 1607319584
transform 1 0 396 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_130
timestamp 1607319584
transform -1 0 452 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_776
timestamp 1607319584
transform 1 0 452 0 1 3705
box -2 -3 98 103
use FILL  FILL_37_0_0
timestamp 1607319584
transform 1 0 548 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_0_1
timestamp 1607319584
transform 1 0 556 0 1 3705
box -2 -3 10 103
use INVX1  INVX1_494
timestamp 1607319584
transform 1 0 564 0 1 3705
box -2 -3 18 103
use CLKBUF1  CLKBUF1_92
timestamp 1607319584
transform -1 0 652 0 1 3705
box -2 -3 74 103
use NAND2X1  NAND2X1_738
timestamp 1607319584
transform -1 0 676 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_607
timestamp 1607319584
transform 1 0 676 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_134
timestamp 1607319584
transform -1 0 732 0 1 3705
box -2 -3 26 103
use MUX2X1  MUX2X1_83
timestamp 1607319584
transform -1 0 780 0 1 3705
box -2 -3 50 103
use NOR2X1  NOR2X1_120
timestamp 1607319584
transform -1 0 804 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_799
timestamp 1607319584
transform 1 0 804 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_654
timestamp 1607319584
transform 1 0 900 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_152
timestamp 1607319584
transform -1 0 956 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_901
timestamp 1607319584
transform -1 0 988 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1278
timestamp 1607319584
transform 1 0 988 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_902
timestamp 1607319584
transform 1 0 1020 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_1_0
timestamp 1607319584
transform -1 0 1060 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_1_1
timestamp 1607319584
transform -1 0 1068 0 1 3705
box -2 -3 10 103
use NAND2X1  NAND2X1_328
timestamp 1607319584
transform -1 0 1092 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1149
timestamp 1607319584
transform 1 0 1092 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_396
timestamp 1607319584
transform -1 0 1148 0 1 3705
box -2 -3 26 103
use BUFX4  BUFX4_116
timestamp 1607319584
transform -1 0 1180 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_707
timestamp 1607319584
transform -1 0 1276 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_594
timestamp 1607319584
transform 1 0 1276 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_539
timestamp 1607319584
transform 1 0 1300 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_540
timestamp 1607319584
transform -1 0 1364 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_718
timestamp 1607319584
transform -1 0 1460 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_669
timestamp 1607319584
transform -1 0 1484 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_791
timestamp 1607319584
transform 1 0 1484 0 1 3705
box -2 -3 98 103
use FILL  FILL_37_2_0
timestamp 1607319584
transform 1 0 1580 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_2_1
timestamp 1607319584
transform 1 0 1588 0 1 3705
box -2 -3 10 103
use INVX1  INVX1_430
timestamp 1607319584
transform 1 0 1596 0 1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_606
timestamp 1607319584
transform 1 0 1612 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_133
timestamp 1607319584
transform -1 0 1668 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_576
timestamp 1607319584
transform -1 0 1692 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_437
timestamp 1607319584
transform -1 0 1716 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_416
timestamp 1607319584
transform 1 0 1716 0 1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_127
timestamp 1607319584
transform -1 0 1764 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_397
timestamp 1607319584
transform -1 0 1788 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_966
timestamp 1607319584
transform -1 0 1820 0 1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_261
timestamp 1607319584
transform -1 0 1868 0 1 3705
box -2 -3 50 103
use OAI21X1  OAI21X1_125
timestamp 1607319584
transform 1 0 1868 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_126
timestamp 1607319584
transform -1 0 1932 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_427
timestamp 1607319584
transform 1 0 1932 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_268
timestamp 1607319584
transform 1 0 2028 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_653
timestamp 1607319584
transform 1 0 2052 0 1 3705
box -2 -3 26 103
use FILL  FILL_37_3_0
timestamp 1607319584
transform 1 0 2076 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_3_1
timestamp 1607319584
transform 1 0 2084 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_729
timestamp 1607319584
transform 1 0 2092 0 1 3705
box -2 -3 98 103
use NOR2X1  NOR2X1_83
timestamp 1607319584
transform 1 0 2188 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_65
timestamp 1607319584
transform -1 0 2244 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_368
timestamp 1607319584
transform -1 0 2268 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_178
timestamp 1607319584
transform -1 0 2284 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_851
timestamp 1607319584
transform -1 0 2380 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_655
timestamp 1607319584
transform 1 0 2380 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_153
timestamp 1607319584
transform -1 0 2436 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_140
timestamp 1607319584
transform -1 0 2468 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_434
timestamp 1607319584
transform -1 0 2564 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_703
timestamp 1607319584
transform 1 0 2564 0 1 3705
box -2 -3 26 103
use FILL  FILL_37_4_0
timestamp 1607319584
transform 1 0 2588 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_4_1
timestamp 1607319584
transform 1 0 2596 0 1 3705
box -2 -3 10 103
use INVX8  INVX8_2
timestamp 1607319584
transform 1 0 2604 0 1 3705
box -2 -3 42 103
use OAI21X1  OAI21X1_1617
timestamp 1607319584
transform 1 0 2644 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1616
timestamp 1607319584
transform -1 0 2708 0 1 3705
box -2 -3 34 103
use MUX2X1  MUX2X1_117
timestamp 1607319584
transform -1 0 2756 0 1 3705
box -2 -3 50 103
use CLKBUF1  CLKBUF1_49
timestamp 1607319584
transform -1 0 2828 0 1 3705
box -2 -3 74 103
use BUFX4  BUFX4_79
timestamp 1607319584
transform -1 0 2860 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_93
timestamp 1607319584
transform -1 0 2884 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_73
timestamp 1607319584
transform -1 0 2916 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_745
timestamp 1607319584
transform -1 0 3012 0 1 3705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_39
timestamp 1607319584
transform 1 0 3012 0 1 3705
box -2 -3 74 103
use FILL  FILL_37_5_0
timestamp 1607319584
transform 1 0 3084 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_5_1
timestamp 1607319584
transform 1 0 3092 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1607319584
transform 1 0 3100 0 1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_251
timestamp 1607319584
transform 1 0 3196 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_316
timestamp 1607319584
transform -1 0 3252 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1607319584
transform 1 0 3252 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_485
timestamp 1607319584
transform -1 0 3372 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_855
timestamp 1607319584
transform -1 0 3404 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_368
timestamp 1607319584
transform -1 0 3428 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_259
timestamp 1607319584
transform -1 0 3524 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_843
timestamp 1607319584
transform 1 0 3524 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1589
timestamp 1607319584
transform 1 0 3548 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_114
timestamp 1607319584
transform -1 0 3612 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_6_0
timestamp 1607319584
transform 1 0 3612 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_6_1
timestamp 1607319584
transform 1 0 3620 0 1 3705
box -2 -3 10 103
use INVX2  INVX2_10
timestamp 1607319584
transform 1 0 3628 0 1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_842
timestamp 1607319584
transform -1 0 3668 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_861
timestamp 1607319584
transform 1 0 3668 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_860
timestamp 1607319584
transform 1 0 3692 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1047
timestamp 1607319584
transform -1 0 3748 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1607319584
transform -1 0 3844 0 1 3705
box -2 -3 98 103
use AOI21X1  AOI21X1_203
timestamp 1607319584
transform -1 0 3876 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_240
timestamp 1607319584
transform 1 0 3876 0 1 3705
box -2 -3 26 103
use BUFX4  BUFX4_151
timestamp 1607319584
transform 1 0 3900 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_292
timestamp 1607319584
transform 1 0 3932 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1607319584
transform 1 0 3956 0 1 3705
box -2 -3 98 103
use BUFX4  BUFX4_112
timestamp 1607319584
transform 1 0 4052 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_246
timestamp 1607319584
transform 1 0 4084 0 1 3705
box -2 -3 26 103
use FILL  FILL_37_7_0
timestamp 1607319584
transform 1 0 4108 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_7_1
timestamp 1607319584
transform 1 0 4116 0 1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1398
timestamp 1607319584
transform 1 0 4124 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1607319584
transform -1 0 4252 0 1 3705
box -2 -3 98 103
use MUX2X1  MUX2X1_291
timestamp 1607319584
transform 1 0 4252 0 1 3705
box -2 -3 50 103
use OAI21X1  OAI21X1_1052
timestamp 1607319584
transform -1 0 4332 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1243
timestamp 1607319584
transform 1 0 4332 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_696
timestamp 1607319584
transform -1 0 4388 0 1 3705
box -2 -3 26 103
use MUX2X1  MUX2X1_290
timestamp 1607319584
transform -1 0 4436 0 1 3705
box -2 -3 50 103
use NAND2X1  NAND2X1_276
timestamp 1607319584
transform 1 0 4436 0 1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1607319584
transform -1 0 4556 0 1 3705
box -2 -3 98 103
use MUX2X1  MUX2X1_289
timestamp 1607319584
transform -1 0 4604 0 1 3705
box -2 -3 50 103
use NAND2X1  NAND2X1_487
timestamp 1607319584
transform 1 0 4604 0 1 3705
box -2 -3 26 103
use FILL  FILL_37_8_0
timestamp 1607319584
transform -1 0 4636 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_8_1
timestamp 1607319584
transform -1 0 4644 0 1 3705
box -2 -3 10 103
use NOR2X1  NOR2X1_338
timestamp 1607319584
transform -1 0 4668 0 1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_268
timestamp 1607319584
transform -1 0 4700 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1177
timestamp 1607319584
transform -1 0 4732 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_625
timestamp 1607319584
transform 1 0 4732 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_389
timestamp 1607319584
transform -1 0 4772 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1607319584
transform -1 0 4868 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_155
timestamp 1607319584
transform 1 0 4868 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_1422
timestamp 1607319584
transform 1 0 4964 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1607319584
transform -1 0 5092 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_176
timestamp 1607319584
transform -1 0 5188 0 1 3705
box -2 -3 98 103
use FILL  FILL_38_1
timestamp 1607319584
transform 1 0 5188 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_797
timestamp 1607319584
transform 1 0 4 0 -1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_789
timestamp 1607319584
transform -1 0 196 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_302
timestamp 1607319584
transform 1 0 196 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_604
timestamp 1607319584
transform 1 0 212 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_131
timestamp 1607319584
transform -1 0 268 0 -1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_800
timestamp 1607319584
transform 1 0 268 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_903
timestamp 1607319584
transform 1 0 364 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_904
timestamp 1607319584
transform -1 0 428 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_116
timestamp 1607319584
transform -1 0 444 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_792
timestamp 1607319584
transform 1 0 444 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_0_0
timestamp 1607319584
transform 1 0 540 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_0_1
timestamp 1607319584
transform 1 0 548 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_738
timestamp 1607319584
transform 1 0 556 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_107
timestamp 1607319584
transform 1 0 652 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_850
timestamp 1607319584
transform 1 0 668 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_114
timestamp 1607319584
transform 1 0 764 0 -1 3905
box -2 -3 18 103
use MUX2X1  MUX2X1_180
timestamp 1607319584
transform -1 0 828 0 -1 3905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_736
timestamp 1607319584
transform 1 0 828 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_361
timestamp 1607319584
transform 1 0 924 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_177
timestamp 1607319584
transform 1 0 940 0 -1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_733
timestamp 1607319584
transform 1 0 956 0 -1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_90
timestamp 1607319584
transform 1 0 980 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_72
timestamp 1607319584
transform -1 0 1036 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_1_0
timestamp 1607319584
transform 1 0 1036 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_1_1
timestamp 1607319584
transform 1 0 1044 0 -1 3905
box -2 -3 10 103
use MUX2X1  MUX2X1_14
timestamp 1607319584
transform 1 0 1052 0 -1 3905
box -2 -3 50 103
use NOR2X1  NOR2X1_155
timestamp 1607319584
transform -1 0 1124 0 -1 3905
box -2 -3 26 103
use INVX1  INVX1_425
timestamp 1607319584
transform 1 0 1124 0 -1 3905
box -2 -3 18 103
use NOR2X1  NOR2X1_144
timestamp 1607319584
transform 1 0 1140 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_517
timestamp 1607319584
transform 1 0 1164 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_420
timestamp 1607319584
transform -1 0 1292 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_233
timestamp 1607319584
transform 1 0 1292 0 -1 3905
box -2 -3 18 103
use NOR2X1  NOR2X1_146
timestamp 1607319584
transform 1 0 1308 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_111
timestamp 1607319584
transform -1 0 1364 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_112
timestamp 1607319584
transform -1 0 1396 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_264
timestamp 1607319584
transform -1 0 1428 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1607319584
transform -1 0 1452 0 -1 3905
box -2 -3 26 103
use INVX1  INVX1_215
timestamp 1607319584
transform 1 0 1452 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1266
timestamp 1607319584
transform 1 0 1468 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_260
timestamp 1607319584
transform 1 0 1500 0 -1 3905
box -2 -3 50 103
use FILL  FILL_38_2_0
timestamp 1607319584
transform -1 0 1556 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_2_1
timestamp 1607319584
transform -1 0 1564 0 -1 3905
box -2 -3 10 103
use MUX2X1  MUX2X1_355
timestamp 1607319584
transform -1 0 1612 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_1003
timestamp 1607319584
transform 1 0 1612 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_158
timestamp 1607319584
transform 1 0 1644 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_1004
timestamp 1607319584
transform -1 0 1724 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_216
timestamp 1607319584
transform -1 0 1740 0 -1 3905
box -2 -3 18 103
use MUX2X1  MUX2X1_357
timestamp 1607319584
transform 1 0 1740 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_1201
timestamp 1607319584
transform 1 0 1788 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1140
timestamp 1607319584
transform -1 0 1852 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_51
timestamp 1607319584
transform -1 0 1876 0 -1 3905
box -2 -3 26 103
use MUX2X1  MUX2X1_324
timestamp 1607319584
transform 1 0 1876 0 -1 3905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_551
timestamp 1607319584
transform -1 0 2020 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_415
timestamp 1607319584
transform 1 0 2020 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_271
timestamp 1607319584
transform 1 0 2036 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_3_0
timestamp 1607319584
transform -1 0 2076 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_3_1
timestamp 1607319584
transform -1 0 2084 0 -1 3905
box -2 -3 10 103
use NAND2X1  NAND2X1_64
timestamp 1607319584
transform -1 0 2108 0 -1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_59
timestamp 1607319584
transform 1 0 2108 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_47
timestamp 1607319584
transform -1 0 2164 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_259
timestamp 1607319584
transform -1 0 2212 0 -1 3905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_419
timestamp 1607319584
transform 1 0 2212 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_110
timestamp 1607319584
transform 1 0 2308 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_109
timestamp 1607319584
transform 1 0 2340 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_151
timestamp 1607319584
transform 1 0 2372 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_939
timestamp 1607319584
transform 1 0 2388 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_213
timestamp 1607319584
transform 1 0 2420 0 -1 3905
box -2 -3 50 103
use NOR2X1  NOR2X1_156
timestamp 1607319584
transform 1 0 2468 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_125
timestamp 1607319584
transform -1 0 2524 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_344
timestamp 1607319584
transform -1 0 2572 0 -1 3905
box -2 -3 50 103
use FILL  FILL_38_4_0
timestamp 1607319584
transform -1 0 2580 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_4_1
timestamp 1607319584
transform -1 0 2588 0 -1 3905
box -2 -3 10 103
use MUX2X1  MUX2X1_41
timestamp 1607319584
transform -1 0 2636 0 -1 3905
box -2 -3 50 103
use MUX2X1  MUX2X1_110
timestamp 1607319584
transform 1 0 2636 0 -1 3905
box -2 -3 50 103
use MUX2X1  MUX2X1_116
timestamp 1607319584
transform -1 0 2732 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_847
timestamp 1607319584
transform -1 0 2764 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_269
timestamp 1607319584
transform 1 0 2764 0 -1 3905
box -2 -3 26 103
use INVX1  INVX1_280
timestamp 1607319584
transform 1 0 2788 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1068
timestamp 1607319584
transform 1 0 2804 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_59
timestamp 1607319584
transform -1 0 2852 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_737
timestamp 1607319584
transform -1 0 2948 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_553
timestamp 1607319584
transform 1 0 2948 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1251
timestamp 1607319584
transform -1 0 3012 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1110
timestamp 1607319584
transform 1 0 3012 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_553
timestamp 1607319584
transform 1 0 3044 0 -1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_859
timestamp 1607319584
transform 1 0 3068 0 -1 3905
box -2 -3 26 103
use FILL  FILL_38_5_0
timestamp 1607319584
transform 1 0 3092 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_5_1
timestamp 1607319584
transform 1 0 3100 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_299
timestamp 1607319584
transform 1 0 3108 0 -1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_372
timestamp 1607319584
transform 1 0 3204 0 -1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_360
timestamp 1607319584
transform -1 0 3252 0 -1 3905
box -2 -3 26 103
use MUX2X1  MUX2X1_47
timestamp 1607319584
transform 1 0 3252 0 -1 3905
box -2 -3 50 103
use MUX2X1  MUX2X1_48
timestamp 1607319584
transform -1 0 3348 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_931
timestamp 1607319584
transform -1 0 3380 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_636
timestamp 1607319584
transform 1 0 3380 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1187
timestamp 1607319584
transform -1 0 3436 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_296
timestamp 1607319584
transform 1 0 3436 0 -1 3905
box -2 -3 50 103
use NOR2X1  NOR2X1_376
timestamp 1607319584
transform -1 0 3508 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_300
timestamp 1607319584
transform -1 0 3540 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_258
timestamp 1607319584
transform 1 0 3540 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_6_0
timestamp 1607319584
transform -1 0 3644 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_6_1
timestamp 1607319584
transform -1 0 3652 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1588
timestamp 1607319584
transform -1 0 3684 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_454
timestamp 1607319584
transform -1 0 3716 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_191
timestamp 1607319584
transform 1 0 3716 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_1652
timestamp 1607319584
transform 1 0 3764 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1653
timestamp 1607319584
transform -1 0 3828 0 -1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_192
timestamp 1607319584
transform -1 0 3876 0 -1 3905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1607319584
transform -1 0 3972 0 -1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_314
timestamp 1607319584
transform 1 0 3972 0 -1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_249
timestamp 1607319584
transform -1 0 4028 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1607319584
transform 1 0 4028 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_7_0
timestamp 1607319584
transform 1 0 4124 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_7_1
timestamp 1607319584
transform 1 0 4132 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1397
timestamp 1607319584
transform 1 0 4140 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_348
timestamp 1607319584
transform -1 0 4196 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1393
timestamp 1607319584
transform 1 0 4196 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1394
timestamp 1607319584
transform -1 0 4260 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1607319584
transform -1 0 4356 0 -1 3905
box -2 -3 98 103
use MUX2X1  MUX2X1_46
timestamp 1607319584
transform -1 0 4404 0 -1 3905
box -2 -3 50 103
use MUX2X1  MUX2X1_337
timestamp 1607319584
transform -1 0 4452 0 -1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_853
timestamp 1607319584
transform -1 0 4484 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1347
timestamp 1607319584
transform 1 0 4484 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1348
timestamp 1607319584
transform -1 0 4548 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_399
timestamp 1607319584
transform -1 0 4564 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_295
timestamp 1607319584
transform -1 0 4660 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_8_0
timestamp 1607319584
transform -1 0 4668 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_8_1
timestamp 1607319584
transform -1 0 4676 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1632
timestamp 1607319584
transform -1 0 4708 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_264
timestamp 1607319584
transform -1 0 4724 0 -1 3905
box -2 -3 18 103
use BUFX4  BUFX4_388
timestamp 1607319584
transform 1 0 4724 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1429
timestamp 1607319584
transform 1 0 4756 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1430
timestamp 1607319584
transform -1 0 4820 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1437
timestamp 1607319584
transform 1 0 4820 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1438
timestamp 1607319584
transform -1 0 4884 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1607319584
transform -1 0 4980 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_133
timestamp 1607319584
transform -1 0 4996 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1421
timestamp 1607319584
transform -1 0 5028 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1409
timestamp 1607319584
transform 1 0 5028 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1410
timestamp 1607319584
transform -1 0 5092 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1607319584
transform -1 0 5188 0 -1 3905
box -2 -3 98 103
use FILL  FILL_39_1
timestamp 1607319584
transform -1 0 5196 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_746
timestamp 1607319584
transform 1 0 4 0 1 3905
box -2 -3 98 103
use AOI21X1  AOI21X1_74
timestamp 1607319584
transform 1 0 100 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_94
timestamp 1607319584
transform -1 0 156 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_94
timestamp 1607319584
transform 1 0 156 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_118
timestamp 1607319584
transform -1 0 212 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_856
timestamp 1607319584
transform 1 0 212 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_330
timestamp 1607319584
transform -1 0 332 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_498
timestamp 1607319584
transform 1 0 332 0 1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_660
timestamp 1607319584
transform 1 0 348 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_329
timestamp 1607319584
transform -1 0 404 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_158
timestamp 1607319584
transform -1 0 428 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_668
timestamp 1607319584
transform 1 0 428 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_166
timestamp 1607319584
transform -1 0 484 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_882
timestamp 1607319584
transform -1 0 580 0 1 3905
box -2 -3 98 103
use FILL  FILL_39_0_0
timestamp 1607319584
transform 1 0 580 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_0_1
timestamp 1607319584
transform 1 0 588 0 1 3905
box -2 -3 10 103
use NAND2X1  NAND2X1_116
timestamp 1607319584
transform 1 0 596 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_744
timestamp 1607319584
transform -1 0 716 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_554
timestamp 1607319584
transform -1 0 748 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_710
timestamp 1607319584
transform 1 0 748 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_524
timestamp 1607319584
transform 1 0 844 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_523
timestamp 1607319584
transform -1 0 908 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_858
timestamp 1607319584
transform 1 0 908 0 1 3905
box -2 -3 98 103
use MUX2X1  MUX2X1_364
timestamp 1607319584
transform -1 0 1052 0 1 3905
box -2 -3 50 103
use FILL  FILL_39_1_0
timestamp 1607319584
transform 1 0 1052 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_1_1
timestamp 1607319584
transform 1 0 1060 0 1 3905
box -2 -3 10 103
use AOI21X1  AOI21X1_118
timestamp 1607319584
transform 1 0 1068 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_148
timestamp 1607319584
transform 1 0 1100 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_525
timestamp 1607319584
transform -1 0 1156 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_320
timestamp 1607319584
transform -1 0 1180 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_518
timestamp 1607319584
transform -1 0 1212 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_895
timestamp 1607319584
transform -1 0 1244 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_63
timestamp 1607319584
transform -1 0 1268 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_293
timestamp 1607319584
transform -1 0 1300 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_294
timestamp 1607319584
transform -1 0 1332 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_536
timestamp 1607319584
transform 1 0 1332 0 1 3905
box -2 -3 98 103
use INVX1  INVX1_478
timestamp 1607319584
transform 1 0 1428 0 1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_446
timestamp 1607319584
transform 1 0 1444 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_721
timestamp 1607319584
transform -1 0 1564 0 1 3905
box -2 -3 26 103
use FILL  FILL_39_2_0
timestamp 1607319584
transform 1 0 1564 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_2_1
timestamp 1607319584
transform 1 0 1572 0 1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_163
timestamp 1607319584
transform 1 0 1580 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_164
timestamp 1607319584
transform -1 0 1644 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_160
timestamp 1607319584
transform 1 0 1644 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_159
timestamp 1607319584
transform 1 0 1676 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_438
timestamp 1607319584
transform -1 0 1732 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_297
timestamp 1607319584
transform 1 0 1732 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_652
timestamp 1607319584
transform 1 0 1764 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1202
timestamp 1607319584
transform -1 0 1820 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_585
timestamp 1607319584
transform 1 0 1820 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_651
timestamp 1607319584
transform 1 0 1844 0 1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_52
timestamp 1607319584
transform -1 0 1892 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_436
timestamp 1607319584
transform -1 0 1988 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_144
timestamp 1607319584
transform -1 0 2020 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_143
timestamp 1607319584
transform -1 0 2052 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_3_0
timestamp 1607319584
transform -1 0 2060 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_3_1
timestamp 1607319584
transform -1 0 2068 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_559
timestamp 1607319584
transform -1 0 2164 0 1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_871
timestamp 1607319584
transform 1 0 2164 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_164
timestamp 1607319584
transform 1 0 2260 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_666
timestamp 1607319584
transform -1 0 2316 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_435
timestamp 1607319584
transform 1 0 2316 0 1 3905
box -2 -3 18 103
use MUX2X1  MUX2X1_11
timestamp 1607319584
transform -1 0 2380 0 1 3905
box -2 -3 50 103
use MUX2X1  MUX2X1_13
timestamp 1607319584
transform 1 0 2380 0 1 3905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_865
timestamp 1607319584
transform -1 0 2524 0 1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_41
timestamp 1607319584
transform 1 0 2524 0 1 3905
box -2 -3 26 103
use FILL  FILL_39_4_0
timestamp 1607319584
transform -1 0 2556 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_4_1
timestamp 1607319584
transform -1 0 2564 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_272
timestamp 1607319584
transform -1 0 2660 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_940
timestamp 1607319584
transform -1 0 2692 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_152
timestamp 1607319584
transform -1 0 2708 0 1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_141
timestamp 1607319584
transform -1 0 2740 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1607319584
transform -1 0 2772 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_848
timestamp 1607319584
transform 1 0 2772 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_145
timestamp 1607319584
transform 1 0 2804 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_507
timestamp 1607319584
transform -1 0 2860 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_146
timestamp 1607319584
transform 1 0 2860 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_437
timestamp 1607319584
transform 1 0 2892 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_109
timestamp 1607319584
transform -1 0 3012 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_170
timestamp 1607319584
transform -1 0 3044 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_705
timestamp 1607319584
transform 1 0 3044 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1633
timestamp 1607319584
transform -1 0 3100 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_5_0
timestamp 1607319584
transform -1 0 3108 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_5_1
timestamp 1607319584
transform -1 0 3116 0 1 3905
box -2 -3 10 103
use INVX1  INVX1_463
timestamp 1607319584
transform -1 0 3132 0 1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_296
timestamp 1607319584
transform -1 0 3228 0 1 3905
box -2 -3 98 103
use AOI21X1  AOI21X1_296
timestamp 1607319584
transform -1 0 3260 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_322
timestamp 1607319584
transform -1 0 3276 0 1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1607319584
transform -1 0 3372 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_278
timestamp 1607319584
transform -1 0 3396 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1366
timestamp 1607319584
transform 1 0 3396 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_799
timestamp 1607319584
transform -1 0 3452 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_291
timestamp 1607319584
transform 1 0 3452 0 1 3905
box -2 -3 98 103
use INVX1  INVX1_143
timestamp 1607319584
transform 1 0 3548 0 1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1628
timestamp 1607319584
transform 1 0 3564 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_854
timestamp 1607319584
transform -1 0 3620 0 1 3905
box -2 -3 26 103
use FILL  FILL_39_6_0
timestamp 1607319584
transform 1 0 3620 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_6_1
timestamp 1607319584
transform 1 0 3628 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_313
timestamp 1607319584
transform 1 0 3636 0 1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_303
timestamp 1607319584
transform -1 0 3828 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_242
timestamp 1607319584
transform 1 0 3828 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1607319584
transform -1 0 3948 0 1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_305
timestamp 1607319584
transform 1 0 3948 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_244
timestamp 1607319584
transform -1 0 4004 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_314
timestamp 1607319584
transform -1 0 4100 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_347
timestamp 1607319584
transform 1 0 4100 0 1 3905
box -2 -3 26 103
use FILL  FILL_39_7_0
timestamp 1607319584
transform 1 0 4124 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_7_1
timestamp 1607319584
transform 1 0 4132 0 1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_826
timestamp 1607319584
transform 1 0 4140 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_622
timestamp 1607319584
transform -1 0 4196 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_245
timestamp 1607319584
transform 1 0 4196 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_919
timestamp 1607319584
transform 1 0 4220 0 1 3905
box -2 -3 34 103
use MUX2X1  MUX2X1_95
timestamp 1607319584
transform 1 0 4252 0 1 3905
box -2 -3 50 103
use OAI21X1  OAI21X1_920
timestamp 1607319584
transform -1 0 4332 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_306
timestamp 1607319584
transform 1 0 4332 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_245
timestamp 1607319584
transform -1 0 4388 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_299
timestamp 1607319584
transform -1 0 4412 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_814
timestamp 1607319584
transform 1 0 4412 0 1 3905
box -2 -3 26 103
use MUX2X1  MUX2X1_338
timestamp 1607319584
transform -1 0 4484 0 1 3905
box -2 -3 50 103
use BUFX4  BUFX4_463
timestamp 1607319584
transform 1 0 4484 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_297
timestamp 1607319584
transform -1 0 4540 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_854
timestamp 1607319584
transform 1 0 4540 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_277
timestamp 1607319584
transform -1 0 4596 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1241
timestamp 1607319584
transform -1 0 4628 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_8_0
timestamp 1607319584
transform 1 0 4628 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_8_1
timestamp 1607319584
transform 1 0 4636 0 1 3905
box -2 -3 10 103
use NAND2X1  NAND2X1_490
timestamp 1607319584
transform 1 0 4644 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_858
timestamp 1607319584
transform 1 0 4668 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_795
timestamp 1607319584
transform 1 0 4692 0 1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1362
timestamp 1607319584
transform -1 0 4748 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_66
timestamp 1607319584
transform -1 0 4764 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_855
timestamp 1607319584
transform 1 0 4764 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1607319584
transform 1 0 4788 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1433
timestamp 1607319584
transform 1 0 4884 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1434
timestamp 1607319584
transform 1 0 4916 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1607319584
transform -1 0 5044 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_1414
timestamp 1607319584
transform 1 0 5044 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1413
timestamp 1607319584
transform -1 0 5108 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_453
timestamp 1607319584
transform -1 0 5124 0 1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1423
timestamp 1607319584
transform 1 0 5124 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1424
timestamp 1607319584
transform -1 0 5188 0 1 3905
box -2 -3 34 103
use FILL  FILL_40_1
timestamp 1607319584
transform 1 0 5188 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_752
timestamp 1607319584
transform 1 0 4 0 -1 4105
box -2 -3 98 103
use AOI21X1  AOI21X1_80
timestamp 1607319584
transform 1 0 100 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_100
timestamp 1607319584
transform -1 0 156 0 -1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_866
timestamp 1607319584
transform 1 0 156 0 -1 4105
box -2 -3 98 103
use INVX1  INVX1_115
timestamp 1607319584
transform 1 0 252 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_661
timestamp 1607319584
transform 1 0 268 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1607319584
transform -1 0 324 0 -1 4105
box -2 -3 26 103
use MUX2X1  MUX2X1_370
timestamp 1607319584
transform 1 0 324 0 -1 4105
box -2 -3 50 103
use MUX2X1  MUX2X1_371
timestamp 1607319584
transform 1 0 372 0 -1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_1288
timestamp 1607319584
transform -1 0 452 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_170
timestamp 1607319584
transform -1 0 476 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_734
timestamp 1607319584
transform -1 0 500 0 -1 4105
box -2 -3 26 103
use INVX1  INVX1_500
timestamp 1607319584
transform -1 0 516 0 -1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_172
timestamp 1607319584
transform -1 0 540 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_0_0
timestamp 1607319584
transform -1 0 548 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_0_1
timestamp 1607319584
transform -1 0 556 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1279
timestamp 1607319584
transform -1 0 588 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_560
timestamp 1607319584
transform 1 0 588 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_491
timestamp 1607319584
transform -1 0 636 0 -1 4105
box -2 -3 18 103
use MUX2X1  MUX2X1_365
timestamp 1607319584
transform 1 0 636 0 -1 4105
box -2 -3 50 103
use BUFX4  BUFX4_299
timestamp 1607319584
transform -1 0 716 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_110
timestamp 1607319584
transform -1 0 740 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_156
timestamp 1607319584
transform -1 0 764 0 -1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_852
timestamp 1607319584
transform 1 0 764 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_656
timestamp 1607319584
transform -1 0 892 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_154
timestamp 1607319584
transform -1 0 916 0 -1 4105
box -2 -3 26 103
use MUX2X1  MUX2X1_276
timestamp 1607319584
transform 1 0 916 0 -1 4105
box -2 -3 50 103
use MUX2X1  MUX2X1_366
timestamp 1607319584
transform -1 0 1012 0 -1 4105
box -2 -3 50 103
use FILL  FILL_40_1_0
timestamp 1607319584
transform 1 0 1012 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_1_1
timestamp 1607319584
transform 1 0 1020 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_711
timestamp 1607319584
transform 1 0 1028 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_526
timestamp 1607319584
transform -1 0 1156 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_118
timestamp 1607319584
transform 1 0 1156 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_845
timestamp 1607319584
transform 1 0 1188 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_105
timestamp 1607319584
transform 1 0 1220 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_270
timestamp 1607319584
transform -1 0 1268 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_550
timestamp 1607319584
transform 1 0 1268 0 -1 4105
box -2 -3 98 103
use INVX1  INVX1_351
timestamp 1607319584
transform 1 0 1364 0 -1 4105
box -2 -3 18 103
use NOR2X1  NOR2X1_102
timestamp 1607319584
transform 1 0 1380 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1139
timestamp 1607319584
transform 1 0 1404 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_297
timestamp 1607319584
transform 1 0 1436 0 -1 4105
box -2 -3 18 103
use MUX2X1  MUX2X1_164
timestamp 1607319584
transform 1 0 1452 0 -1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_1012
timestamp 1607319584
transform 1 0 1500 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_53
timestamp 1607319584
transform -1 0 1556 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_2_0
timestamp 1607319584
transform -1 0 1564 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_2_1
timestamp 1607319584
transform -1 0 1572 0 -1 4105
box -2 -3 10 103
use MUX2X1  MUX2X1_165
timestamp 1607319584
transform -1 0 1620 0 -1 4105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_444
timestamp 1607319584
transform 1 0 1620 0 -1 4105
box -2 -3 98 103
use MUX2X1  MUX2X1_69
timestamp 1607319584
transform -1 0 1764 0 -1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_1267
timestamp 1607319584
transform 1 0 1764 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_722
timestamp 1607319584
transform -1 0 1820 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1268
timestamp 1607319584
transform 1 0 1820 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_356
timestamp 1607319584
transform -1 0 1900 0 -1 4105
box -2 -3 50 103
use BUFX4  BUFX4_287
timestamp 1607319584
transform 1 0 1900 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_253
timestamp 1607319584
transform 1 0 1932 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1607319584
transform -1 0 1988 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_254
timestamp 1607319584
transform 1 0 1988 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_527
timestamp 1607319584
transform -1 0 2116 0 -1 4105
box -2 -3 98 103
use FILL  FILL_40_3_0
timestamp 1607319584
transform -1 0 2124 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_3_1
timestamp 1607319584
transform -1 0 2132 0 -1 4105
box -2 -3 10 103
use NOR2X1  NOR2X1_42
timestamp 1607319584
transform -1 0 2156 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_562
timestamp 1607319584
transform 1 0 2156 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1607319584
transform -1 0 2212 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_896
timestamp 1607319584
transform 1 0 2212 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_321
timestamp 1607319584
transform 1 0 2244 0 -1 4105
box -2 -3 26 103
use BUFX4  BUFX4_432
timestamp 1607319584
transform -1 0 2300 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_55
timestamp 1607319584
transform -1 0 2324 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1223
timestamp 1607319584
transform 1 0 2324 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_323
timestamp 1607319584
transform 1 0 2356 0 -1 4105
box -2 -3 50 103
use MUX2X1  MUX2X1_33
timestamp 1607319584
transform -1 0 2452 0 -1 4105
box -2 -3 50 103
use CLKBUF1  CLKBUF1_27
timestamp 1607319584
transform -1 0 2524 0 -1 4105
box -2 -3 74 103
use INVX1  INVX1_160
timestamp 1607319584
transform 1 0 2524 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_158
timestamp 1607319584
transform -1 0 2572 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_4_0
timestamp 1607319584
transform -1 0 2580 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_4_1
timestamp 1607319584
transform -1 0 2588 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_157
timestamp 1607319584
transform -1 0 2620 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_369
timestamp 1607319584
transform -1 0 2644 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_948
timestamp 1607319584
transform 1 0 2644 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_435
timestamp 1607319584
transform -1 0 2772 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_161
timestamp 1607319584
transform 1 0 2772 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_162
timestamp 1607319584
transform -1 0 2836 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_445
timestamp 1607319584
transform -1 0 2932 0 -1 4105
box -2 -3 98 103
use NAND2X1  NAND2X1_58
timestamp 1607319584
transform -1 0 2956 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_52
timestamp 1607319584
transform 1 0 2956 0 -1 4105
box -2 -3 26 103
use MUX2X1  MUX2X1_12
timestamp 1607319584
transform -1 0 3028 0 -1 4105
box -2 -3 50 103
use NOR2X1  NOR2X1_167
timestamp 1607319584
transform -1 0 3052 0 -1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_134
timestamp 1607319584
transform -1 0 3084 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_5_0
timestamp 1607319584
transform -1 0 3092 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_5_1
timestamp 1607319584
transform -1 0 3100 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_881
timestamp 1607319584
transform -1 0 3196 0 -1 4105
box -2 -3 98 103
use INVX1  INVX1_335
timestamp 1607319584
transform 1 0 3196 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_304
timestamp 1607319584
transform -1 0 3308 0 -1 4105
box -2 -3 98 103
use NAND2X1  NAND2X1_801
timestamp 1607319584
transform 1 0 3308 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1631
timestamp 1607319584
transform 1 0 3332 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_857
timestamp 1607319584
transform -1 0 3388 0 -1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_313
timestamp 1607319584
transform 1 0 3388 0 -1 4105
box -2 -3 26 103
use BUFX4  BUFX4_412
timestamp 1607319584
transform 1 0 3412 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_248
timestamp 1607319584
transform -1 0 3476 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_706
timestamp 1607319584
transform -1 0 3500 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1252
timestamp 1607319584
transform -1 0 3532 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_856
timestamp 1607319584
transform 1 0 3532 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1650
timestamp 1607319584
transform 1 0 3564 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_6_0
timestamp 1607319584
transform -1 0 3604 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_6_1
timestamp 1607319584
transform -1 0 3612 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1651
timestamp 1607319584
transform -1 0 3644 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_305
timestamp 1607319584
transform 1 0 3644 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_343
timestamp 1607319584
transform 1 0 3676 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_344
timestamp 1607319584
transform 1 0 3708 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_983
timestamp 1607319584
transform -1 0 3772 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_984
timestamp 1607319584
transform -1 0 3804 0 -1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_143
timestamp 1607319584
transform 1 0 3804 0 -1 4105
box -2 -3 50 103
use BUFX4  BUFX4_286
timestamp 1607319584
transform -1 0 3884 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_452
timestamp 1607319584
transform 1 0 3884 0 -1 4105
box -2 -3 18 103
use MUX2X1  MUX2X1_144
timestamp 1607319584
transform -1 0 3948 0 -1 4105
box -2 -3 50 103
use BUFX4  BUFX4_125
timestamp 1607319584
transform 1 0 3948 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1173
timestamp 1607319584
transform -1 0 4012 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_40
timestamp 1607319584
transform 1 0 4012 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_1048
timestamp 1607319584
transform -1 0 4060 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_486
timestamp 1607319584
transform 1 0 4060 0 -1 4105
box -2 -3 26 103
use MUX2X1  MUX2X1_96
timestamp 1607319584
transform 1 0 4084 0 -1 4105
box -2 -3 50 103
use FILL  FILL_40_7_0
timestamp 1607319584
transform -1 0 4140 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_7_1
timestamp 1607319584
transform -1 0 4148 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1174
timestamp 1607319584
transform -1 0 4180 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1367
timestamp 1607319584
transform 1 0 4180 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_800
timestamp 1607319584
transform -1 0 4236 0 -1 4105
box -2 -3 26 103
use INVX1  INVX1_386
timestamp 1607319584
transform -1 0 4252 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_1401
timestamp 1607319584
transform 1 0 4252 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1402
timestamp 1607319584
transform -1 0 4316 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_132
timestamp 1607319584
transform 1 0 4316 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1607319584
transform -1 0 4428 0 -1 4105
box -2 -3 98 103
use NAND2X1  NAND2X1_815
timestamp 1607319584
transform 1 0 4428 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_995
timestamp 1607319584
transform -1 0 4484 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_65
timestamp 1607319584
transform 1 0 4484 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1607319584
transform -1 0 4596 0 -1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_301
timestamp 1607319584
transform 1 0 4596 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_8_0
timestamp 1607319584
transform -1 0 4628 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_8_1
timestamp 1607319584
transform -1 0 4636 0 -1 4105
box -2 -3 10 103
use AOI21X1  AOI21X1_240
timestamp 1607319584
transform -1 0 4668 0 -1 4105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_55
timestamp 1607319584
transform -1 0 4740 0 -1 4105
box -2 -3 74 103
use INVX1  INVX1_385
timestamp 1607319584
transform -1 0 4756 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_1629
timestamp 1607319584
transform 1 0 4756 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_207
timestamp 1607319584
transform -1 0 4804 0 -1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_292
timestamp 1607319584
transform -1 0 4900 0 -1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1607319584
transform -1 0 4996 0 -1 4105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_68
timestamp 1607319584
transform -1 0 5068 0 -1 4105
box -2 -3 74 103
use NAND2X1  NAND2X1_171
timestamp 1607319584
transform -1 0 5092 0 -1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1607319584
transform -1 0 5188 0 -1 4105
box -2 -3 98 103
use FILL  FILL_41_1
timestamp 1607319584
transform -1 0 5196 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_894
timestamp 1607319584
transform 1 0 4 0 1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_870
timestamp 1607319584
transform 1 0 100 0 1 4105
box -2 -3 98 103
use INVX1  INVX1_371
timestamp 1607319584
transform 1 0 196 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_665
timestamp 1607319584
transform 1 0 212 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_163
timestamp 1607319584
transform -1 0 268 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_744
timestamp 1607319584
transform -1 0 292 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1159
timestamp 1607319584
transform 1 0 292 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_605
timestamp 1607319584
transform -1 0 348 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1286
timestamp 1607319584
transform -1 0 380 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_606
timestamp 1607319584
transform -1 0 404 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1160
timestamp 1607319584
transform -1 0 436 0 1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_275
timestamp 1607319584
transform -1 0 484 0 1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_674
timestamp 1607319584
transform 1 0 484 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_0_0
timestamp 1607319584
transform -1 0 524 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_0_1
timestamp 1607319584
transform -1 0 532 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_888
timestamp 1607319584
transform -1 0 628 0 1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_854
timestamp 1607319584
transform 1 0 628 0 1 4105
box -2 -3 98 103
use INVX1  INVX1_370
timestamp 1607319584
transform 1 0 724 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_658
timestamp 1607319584
transform -1 0 772 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1158
timestamp 1607319584
transform 1 0 772 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_604
timestamp 1607319584
transform -1 0 828 0 1 4105
box -2 -3 26 103
use MUX2X1  MUX2X1_178
timestamp 1607319584
transform 1 0 828 0 1 4105
box -2 -3 50 103
use INVX1  INVX1_242
timestamp 1607319584
transform 1 0 876 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_1030
timestamp 1607319584
transform -1 0 924 0 1 4105
box -2 -3 34 103
use BUFX4  BUFX4_153
timestamp 1607319584
transform -1 0 956 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_327
timestamp 1607319584
transform -1 0 980 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1277
timestamp 1607319584
transform 1 0 980 0 1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_10
timestamp 1607319584
transform 1 0 1012 0 1 4105
box -2 -3 50 103
use FILL  FILL_41_1_0
timestamp 1607319584
transform 1 0 1060 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_1_1
timestamp 1607319584
transform 1 0 1068 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_708
timestamp 1607319584
transform 1 0 1076 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_520
timestamp 1607319584
transform 1 0 1172 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_267
timestamp 1607319584
transform -1 0 1228 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_519
timestamp 1607319584
transform -1 0 1260 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_446
timestamp 1607319584
transform 1 0 1260 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1011
timestamp 1607319584
transform -1 0 1316 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_166
timestamp 1607319584
transform 1 0 1316 0 1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_157
timestamp 1607319584
transform 1 0 1340 0 1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_168
timestamp 1607319584
transform 1 0 1364 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_584
timestamp 1607319584
transform 1 0 1388 0 1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_532
timestamp 1607319584
transform 1 0 1412 0 1 4105
box -2 -3 98 103
use NAND2X1  NAND2X1_447
timestamp 1607319584
transform 1 0 1508 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_260
timestamp 1607319584
transform -1 0 1564 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_2_0
timestamp 1607319584
transform 1 0 1564 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_2_1
timestamp 1607319584
transform 1 0 1572 0 1 4105
box -2 -3 10 103
use INVX1  INVX1_222
timestamp 1607319584
transform 1 0 1580 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_1010
timestamp 1607319584
transform 1 0 1596 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_445
timestamp 1607319584
transform -1 0 1652 0 1 4105
box -2 -3 26 103
use MUX2X1  MUX2X1_163
timestamp 1607319584
transform -1 0 1700 0 1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_1009
timestamp 1607319584
transform 1 0 1700 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_723
timestamp 1607319584
transform -1 0 1756 0 1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_560
timestamp 1607319584
transform -1 0 1852 0 1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_60
timestamp 1607319584
transform 1 0 1852 0 1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_48
timestamp 1607319584
transform -1 0 1908 0 1 4105
box -2 -3 34 103
use BUFX4  BUFX4_411
timestamp 1607319584
transform -1 0 1940 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_299
timestamp 1607319584
transform 1 0 1940 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_300
timestamp 1607319584
transform -1 0 2004 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_574
timestamp 1607319584
transform -1 0 2100 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_3_0
timestamp 1607319584
transform -1 0 2108 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_3_1
timestamp 1607319584
transform -1 0 2116 0 1 4105
box -2 -3 10 103
use NAND2X1  NAND2X1_258
timestamp 1607319584
transform -1 0 2140 0 1 4105
box -2 -3 26 103
use INVX1  INVX1_108
timestamp 1607319584
transform 1 0 2140 0 1 4105
box -2 -3 18 103
use INVX1  INVX1_414
timestamp 1607319584
transform -1 0 2172 0 1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_535
timestamp 1607319584
transform -1 0 2268 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_263
timestamp 1607319584
transform 1 0 2268 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_836
timestamp 1607319584
transform 1 0 2300 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_277
timestamp 1607319584
transform 1 0 2332 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_56
timestamp 1607319584
transform -1 0 2388 0 1 4105
box -2 -3 26 103
use MUX2X1  MUX2X1_32
timestamp 1607319584
transform -1 0 2436 0 1 4105
box -2 -3 50 103
use NOR2X1  NOR2X1_104
timestamp 1607319584
transform 1 0 2436 0 1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_82
timestamp 1607319584
transform -1 0 2492 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_762
timestamp 1607319584
transform -1 0 2588 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_4_0
timestamp 1607319584
transform 1 0 2588 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_4_1
timestamp 1607319584
transform 1 0 2596 0 1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1076
timestamp 1607319584
transform 1 0 2604 0 1 4105
box -2 -3 34 103
use MUX2X1  MUX2X1_212
timestamp 1607319584
transform -1 0 2684 0 1 4105
box -2 -3 50 103
use OAI21X1  OAI21X1_1075
timestamp 1607319584
transform -1 0 2716 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_269
timestamp 1607319584
transform 1 0 2716 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1607319584
transform -1 0 2772 0 1 4105
box -2 -3 26 103
use BUFX4  BUFX4_126
timestamp 1607319584
transform -1 0 2804 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_270
timestamp 1607319584
transform -1 0 2828 0 1 4105
box -2 -3 26 103
use BUFX4  BUFX4_461
timestamp 1607319584
transform -1 0 2860 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_835
timestamp 1607319584
transform -1 0 2892 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1607319584
transform -1 0 2908 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_265
timestamp 1607319584
transform 1 0 2908 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_545
timestamp 1607319584
transform -1 0 3036 0 1 4105
box -2 -3 98 103
use BUFX4  BUFX4_129
timestamp 1607319584
transform 1 0 3036 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_301
timestamp 1607319584
transform 1 0 3068 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_5_0
timestamp 1607319584
transform 1 0 3100 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_5_1
timestamp 1607319584
transform 1 0 3108 0 1 4105
box -2 -3 10 103
use NOR2X1  NOR2X1_377
timestamp 1607319584
transform 1 0 3116 0 1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_294
timestamp 1607319584
transform -1 0 3236 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_1109
timestamp 1607319584
transform 1 0 3236 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_552
timestamp 1607319584
transform 1 0 3268 0 1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1607319584
transform 1 0 3292 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_1665
timestamp 1607319584
transform 1 0 3388 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1664
timestamp 1607319584
transform 1 0 3420 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_315
timestamp 1607319584
transform -1 0 3476 0 1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_250
timestamp 1607319584
transform -1 0 3508 0 1 4105
box -2 -3 34 103
use BUFX4  BUFX4_154
timestamp 1607319584
transform 1 0 3508 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_279
timestamp 1607319584
transform 1 0 3540 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_416
timestamp 1607319584
transform -1 0 3588 0 1 4105
box -2 -3 26 103
use BUFX4  BUFX4_416
timestamp 1607319584
transform 1 0 3588 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_6_0
timestamp 1607319584
transform -1 0 3628 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_6_1
timestamp 1607319584
transform -1 0 3636 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1607319584
transform -1 0 3732 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_1400
timestamp 1607319584
transform 1 0 3732 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_417
timestamp 1607319584
transform 1 0 3764 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1399
timestamp 1607319584
transform -1 0 3820 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1355
timestamp 1607319584
transform 1 0 3820 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1607319584
transform -1 0 3948 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_1356
timestamp 1607319584
transform -1 0 3980 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_621
timestamp 1607319584
transform 1 0 3980 0 1 4105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_25
timestamp 1607319584
transform -1 0 4076 0 1 4105
box -2 -3 74 103
use FILL  FILL_41_7_0
timestamp 1607319584
transform -1 0 4084 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_7_1
timestamp 1607319584
transform -1 0 4092 0 1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1607319584
transform -1 0 4188 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_1357
timestamp 1607319584
transform -1 0 4220 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1358
timestamp 1607319584
transform -1 0 4252 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1607319584
transform -1 0 4348 0 1 4105
box -2 -3 98 103
use AOI21X1  AOI21X1_141
timestamp 1607319584
transform 1 0 4348 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_175
timestamp 1607319584
transform -1 0 4404 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_675
timestamp 1607319584
transform 1 0 4404 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1224
timestamp 1607319584
transform -1 0 4460 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_429
timestamp 1607319584
transform -1 0 4484 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_1331
timestamp 1607319584
transform 1 0 4484 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1439
timestamp 1607319584
transform 1 0 4516 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_694
timestamp 1607319584
transform 1 0 4548 0 1 4105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_895
timestamp 1607319584
transform -1 0 4668 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_8_0
timestamp 1607319584
transform -1 0 4676 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_8_1
timestamp 1607319584
transform -1 0 4684 0 1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1440
timestamp 1607319584
transform -1 0 4716 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1607319584
transform -1 0 4812 0 1 4105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_20
timestamp 1607319584
transform -1 0 4884 0 1 4105
box -2 -3 74 103
use OAI21X1  OAI21X1_1341
timestamp 1607319584
transform 1 0 4884 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1342
timestamp 1607319584
transform -1 0 4948 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1607319584
transform -1 0 5044 0 1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_673
timestamp 1607319584
transform 1 0 5044 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_436
timestamp 1607319584
transform -1 0 5092 0 1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_887
timestamp 1607319584
transform 1 0 5092 0 1 4105
box -2 -3 98 103
use FILL  FILL_42_1
timestamp 1607319584
transform 1 0 5188 0 1 4105
box -2 -3 10 103
use NOR2X1  NOR2X1_174
timestamp 1607319584
transform -1 0 28 0 -1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_140
timestamp 1607319584
transform -1 0 60 0 -1 4305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_13
timestamp 1607319584
transform -1 0 132 0 -1 4305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_874
timestamp 1607319584
transform 1 0 132 0 -1 4305
box -2 -3 98 103
use NOR2X1  NOR2X1_159
timestamp 1607319584
transform 1 0 228 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_886
timestamp 1607319584
transform 1 0 252 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_372
timestamp 1607319584
transform 1 0 348 0 -1 4305
box -2 -3 18 103
use AOI21X1  AOI21X1_122
timestamp 1607319584
transform 1 0 364 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_152
timestamp 1607319584
transform -1 0 420 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_672
timestamp 1607319584
transform 1 0 420 0 -1 4305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_54
timestamp 1607319584
transform 1 0 452 0 -1 4305
box -2 -3 74 103
use FILL  FILL_42_0_0
timestamp 1607319584
transform 1 0 524 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_0_1
timestamp 1607319584
transform 1 0 532 0 -1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_1280
timestamp 1607319584
transform 1 0 540 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_735
timestamp 1607319584
transform -1 0 596 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_768
timestamp 1607319584
transform -1 0 692 0 -1 4305
box -2 -3 98 103
use NOR2X1  NOR2X1_110
timestamp 1607319584
transform 1 0 692 0 -1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_88
timestamp 1607319584
transform -1 0 748 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_113
timestamp 1607319584
transform 1 0 748 0 -1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_603
timestamp 1607319584
transform -1 0 788 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1157
timestamp 1607319584
transform -1 0 820 0 -1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_274
timestamp 1607319584
transform 1 0 820 0 -1 4305
box -2 -3 50 103
use AOI21X1  AOI21X1_116
timestamp 1607319584
transform 1 0 868 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_145
timestamp 1607319584
transform -1 0 924 0 -1 4305
box -2 -3 26 103
use MUX2X1  MUX2X1_9
timestamp 1607319584
transform 1 0 924 0 -1 4305
box -2 -3 50 103
use INVX1  INVX1_489
timestamp 1607319584
transform 1 0 972 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_529
timestamp 1607319584
transform 1 0 988 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_530
timestamp 1607319584
transform -1 0 1052 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_1_0
timestamp 1607319584
transform 1 0 1052 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_1_1
timestamp 1607319584
transform 1 0 1060 0 -1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_713
timestamp 1607319584
transform 1 0 1068 0 -1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_100
timestamp 1607319584
transform 1 0 1164 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_99
timestamp 1607319584
transform 1 0 1188 0 -1 4305
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1607319584
transform -1 0 1228 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_515
timestamp 1607319584
transform -1 0 1260 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_521
timestamp 1607319584
transform 1 0 1260 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_46
timestamp 1607319584
transform 1 0 1292 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_58
timestamp 1607319584
transform -1 0 1348 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_558
timestamp 1607319584
transform 1 0 1348 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_224
timestamp 1607319584
transform 1 0 1444 0 -1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_576
timestamp 1607319584
transform 1 0 1460 0 -1 4305
box -2 -3 98 103
use FILL  FILL_42_2_0
timestamp 1607319584
transform 1 0 1556 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_2_1
timestamp 1607319584
transform 1 0 1564 0 -1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_304
timestamp 1607319584
transform 1 0 1572 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_303
timestamp 1607319584
transform -1 0 1636 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_301
timestamp 1607319584
transform 1 0 1636 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_302
timestamp 1607319584
transform -1 0 1700 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_575
timestamp 1607319584
transform -1 0 1796 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_413
timestamp 1607319584
transform 1 0 1796 0 -1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_444
timestamp 1607319584
transform -1 0 1836 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_530
timestamp 1607319584
transform 1 0 1836 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_94
timestamp 1607319584
transform 1 0 1932 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_258
timestamp 1607319584
transform 1 0 1948 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1607319584
transform 1 0 1980 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_48
timestamp 1607319584
transform 1 0 2012 0 -1 4305
box -2 -3 26 103
use FILL  FILL_42_3_0
timestamp 1607319584
transform 1 0 2036 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_3_1
timestamp 1607319584
transform 1 0 2044 0 -1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_754
timestamp 1607319584
transform 1 0 2052 0 -1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_67
timestamp 1607319584
transform 1 0 2148 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1138
timestamp 1607319584
transform -1 0 2204 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_352
timestamp 1607319584
transform -1 0 2220 0 -1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_66
timestamp 1607319584
transform 1 0 2220 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1137
timestamp 1607319584
transform -1 0 2276 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_262
timestamp 1607319584
transform 1 0 2276 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_278
timestamp 1607319584
transform 1 0 2308 0 -1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_131
timestamp 1607319584
transform 1 0 2340 0 -1 4305
box -2 -3 50 103
use MUX2X1  MUX2X1_228
timestamp 1607319584
transform 1 0 2388 0 -1 4305
box -2 -3 50 103
use INVX1  INVX1_288
timestamp 1607319584
transform 1 0 2436 0 -1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_443
timestamp 1607319584
transform -1 0 2548 0 -1 4305
box -2 -3 98 103
use FILL  FILL_42_4_0
timestamp 1607319584
transform 1 0 2548 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_4_1
timestamp 1607319584
transform 1 0 2556 0 -1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_549
timestamp 1607319584
transform 1 0 2564 0 -1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_515
timestamp 1607319584
transform 1 0 2660 0 -1 4305
box -2 -3 26 103
use INVX1  INVX1_287
timestamp 1607319584
transform 1 0 2684 0 -1 4305
box -2 -3 18 103
use AOI21X1  AOI21X1_81
timestamp 1607319584
transform 1 0 2700 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_103
timestamp 1607319584
transform -1 0 2756 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_761
timestamp 1607319584
transform 1 0 2756 0 -1 4305
box -2 -3 98 103
use MUX2X1  MUX2X1_31
timestamp 1607319584
transform 1 0 2852 0 -1 4305
box -2 -3 50 103
use OAI21X1  OAI21X1_946
timestamp 1607319584
transform -1 0 2932 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_158
timestamp 1607319584
transform 1 0 2932 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_259
timestamp 1607319584
transform 1 0 2948 0 -1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_115
timestamp 1607319584
transform -1 0 3028 0 -1 4305
box -2 -3 50 103
use AOI21X1  AOI21X1_299
timestamp 1607319584
transform 1 0 3028 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_375
timestamp 1607319584
transform -1 0 3084 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_169
timestamp 1607319584
transform 1 0 3084 0 -1 4305
box -2 -3 26 103
use FILL  FILL_42_5_0
timestamp 1607319584
transform -1 0 3116 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_5_1
timestamp 1607319584
transform -1 0 3124 0 -1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_1123
timestamp 1607319584
transform -1 0 3156 0 -1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_248
timestamp 1607319584
transform 1 0 3156 0 -1 4305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1607319584
transform 1 0 3204 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_450
timestamp 1607319584
transform 1 0 3300 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_1368
timestamp 1607319584
transform -1 0 3348 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1124
timestamp 1607319584
transform -1 0 3380 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_320
timestamp 1607319584
transform 1 0 3380 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1238
timestamp 1607319584
transform 1 0 3476 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_464
timestamp 1607319584
transform 1 0 3508 0 -1 4305
box -2 -3 18 103
use MUX2X1  MUX2X1_334
timestamp 1607319584
transform -1 0 3572 0 -1 4305
box -2 -3 50 103
use OAI21X1  OAI21X1_1237
timestamp 1607319584
transform -1 0 3604 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_6_0
timestamp 1607319584
transform 1 0 3604 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_6_1
timestamp 1607319584
transform 1 0 3612 0 -1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_1188
timestamp 1607319584
transform 1 0 3620 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1607319584
transform -1 0 3748 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1396
timestamp 1607319584
transform -1 0 3780 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_996
timestamp 1607319584
transform 1 0 3780 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1395
timestamp 1607319584
transform -1 0 3844 0 -1 4305
box -2 -3 34 103
use BUFX4  BUFX4_417
timestamp 1607319584
transform 1 0 3844 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_812
timestamp 1607319584
transform 1 0 3876 0 -1 4305
box -2 -3 26 103
use INVX2  INVX2_7
timestamp 1607319584
transform -1 0 3916 0 -1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_792
timestamp 1607319584
transform 1 0 3916 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_793
timestamp 1607319584
transform 1 0 3940 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_811
timestamp 1607319584
transform 1 0 3964 0 -1 4305
box -2 -3 26 103
use INVX1  INVX1_388
timestamp 1607319584
transform 1 0 3988 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_988
timestamp 1607319584
transform -1 0 4036 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_860
timestamp 1607319584
transform -1 0 4068 0 -1 4305
box -2 -3 34 103
use MUX2X1  MUX2X1_94
timestamp 1607319584
transform 1 0 4068 0 -1 4305
box -2 -3 50 103
use FILL  FILL_42_7_0
timestamp 1607319584
transform 1 0 4116 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_7_1
timestamp 1607319584
transform 1 0 4124 0 -1 4305
box -2 -3 10 103
use MUX2X1  MUX2X1_190
timestamp 1607319584
transform 1 0 4132 0 -1 4305
box -2 -3 50 103
use NAND2X1  NAND2X1_833
timestamp 1607319584
transform 1 0 4180 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_832
timestamp 1607319584
transform -1 0 4228 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_917
timestamp 1607319584
transform -1 0 4260 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_798
timestamp 1607319584
transform 1 0 4260 0 -1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_373
timestamp 1607319584
transform -1 0 4308 0 -1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_297
timestamp 1607319584
transform -1 0 4340 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_300
timestamp 1607319584
transform 1 0 4340 0 -1 4305
box -2 -3 98 103
use INVX2  INVX2_8
timestamp 1607319584
transform -1 0 4452 0 -1 4305
box -2 -3 18 103
use BUFX4  BUFX4_391
timestamp 1607319584
transform -1 0 4484 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1332
timestamp 1607319584
transform 1 0 4484 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1607319584
transform -1 0 4612 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_831
timestamp 1607319584
transform -1 0 4644 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_8_0
timestamp 1607319584
transform -1 0 4652 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_8_1
timestamp 1607319584
transform -1 0 4660 0 -1 4305
box -2 -3 10 103
use INVX1  INVX1_44
timestamp 1607319584
transform -1 0 4676 0 -1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_253
timestamp 1607319584
transform 1 0 4676 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_187
timestamp 1607319584
transform -1 0 4796 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1481
timestamp 1607319584
transform 1 0 4796 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1482
timestamp 1607319584
transform -1 0 4860 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_189
timestamp 1607319584
transform -1 0 4956 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1473
timestamp 1607319584
transform 1 0 4956 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1474
timestamp 1607319584
transform -1 0 5020 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_185
timestamp 1607319584
transform -1 0 5116 0 -1 4305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_102
timestamp 1607319584
transform 1 0 5116 0 -1 4305
box -2 -3 74 103
use FILL  FILL_43_1
timestamp 1607319584
transform -1 0 5196 0 -1 4305
box -2 -3 10 103
use NOR2X1  NOR2X1_170
timestamp 1607319584
transform -1 0 28 0 1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_136
timestamp 1607319584
transform -1 0 60 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_890
timestamp 1607319584
transform 1 0 60 0 1 4305
box -2 -3 98 103
use AOI21X1  AOI21X1_127
timestamp 1607319584
transform 1 0 156 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_743
timestamp 1607319584
transform -1 0 212 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1287
timestamp 1607319584
transform -1 0 244 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_499
timestamp 1607319584
transform 1 0 244 0 1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_1285
timestamp 1607319584
transform 1 0 260 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_741
timestamp 1607319584
transform -1 0 316 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_742
timestamp 1607319584
transform -1 0 340 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_862
timestamp 1607319584
transform 1 0 340 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_760
timestamp 1607319584
transform 1 0 436 0 1 4305
box -2 -3 98 103
use FILL  FILL_43_0_0
timestamp 1607319584
transform 1 0 532 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_0_1
timestamp 1607319584
transform 1 0 540 0 1 4305
box -2 -3 10 103
use INVX1  INVX1_492
timestamp 1607319584
transform 1 0 548 0 1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_568
timestamp 1607319584
transform 1 0 564 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_124
timestamp 1607319584
transform -1 0 620 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_648
timestamp 1607319584
transform -1 0 652 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_843
timestamp 1607319584
transform 1 0 652 0 1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_151
timestamp 1607319584
transform -1 0 772 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_642
timestamp 1607319584
transform 1 0 772 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_643
timestamp 1607319584
transform -1 0 836 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_466
timestamp 1607319584
transform -1 0 860 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_849
timestamp 1607319584
transform 1 0 860 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_543
timestamp 1607319584
transform 1 0 956 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_732
timestamp 1607319584
transform 1 0 988 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_544
timestamp 1607319584
transform -1 0 1044 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_1_0
timestamp 1607319584
transform 1 0 1044 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_1_1
timestamp 1607319584
transform 1 0 1052 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_706
timestamp 1607319584
transform 1 0 1060 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_516
timestamp 1607319584
transform 1 0 1156 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_57
timestamp 1607319584
transform 1 0 1188 0 1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_522
timestamp 1607319584
transform 1 0 1204 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_709
timestamp 1607319584
transform 1 0 1236 0 1 4305
box -2 -3 98 103
use NOR2X1  NOR2X1_101
timestamp 1607319584
transform -1 0 1356 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_564
timestamp 1607319584
transform 1 0 1356 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_279
timestamp 1607319584
transform -1 0 1484 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_280
timestamp 1607319584
transform -1 0 1516 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_2_0
timestamp 1607319584
transform -1 0 1524 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_2_1
timestamp 1607319584
transform -1 0 1532 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_544
timestamp 1607319584
transform -1 0 1628 0 1 4305
box -2 -3 98 103
use NOR2X1  NOR2X1_50
timestamp 1607319584
transform 1 0 1628 0 1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_40
timestamp 1607319584
transform -1 0 1684 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_289
timestamp 1607319584
transform 1 0 1684 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_524
timestamp 1607319584
transform 1 0 1716 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_248
timestamp 1607319584
transform 1 0 1812 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_247
timestamp 1607319584
transform -1 0 1876 0 1 4305
box -2 -3 34 103
use BUFX4  BUFX4_433
timestamp 1607319584
transform -1 0 1908 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_674
timestamp 1607319584
transform -1 0 1932 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_542
timestamp 1607319584
transform 1 0 1932 0 1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_583
timestamp 1607319584
transform -1 0 2052 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_252
timestamp 1607319584
transform 1 0 2052 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_3_0
timestamp 1607319584
transform 1 0 2084 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_3_1
timestamp 1607319584
transform 1 0 2092 0 1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_251
timestamp 1607319584
transform 1 0 2100 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_49
timestamp 1607319584
transform 1 0 2132 0 1 4305
box -2 -3 26 103
use INVX2  INVX2_2
timestamp 1607319584
transform 1 0 2156 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_582
timestamp 1607319584
transform 1 0 2172 0 1 4305
box -2 -3 26 103
use INVX1  INVX1_350
timestamp 1607319584
transform -1 0 2212 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_534
timestamp 1607319584
transform -1 0 2308 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_563
timestamp 1607319584
transform 1 0 2308 0 1 4305
box -2 -3 98 103
use MUX2X1  MUX2X1_211
timestamp 1607319584
transform 1 0 2404 0 1 4305
box -2 -3 50 103
use NAND2X1  NAND2X1_157
timestamp 1607319584
transform 1 0 2452 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1074
timestamp 1607319584
transform -1 0 2508 0 1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_45
timestamp 1607319584
transform 1 0 2508 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_57
timestamp 1607319584
transform -1 0 2564 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_516
timestamp 1607319584
transform 1 0 2564 0 1 4305
box -2 -3 26 103
use FILL  FILL_43_4_0
timestamp 1607319584
transform 1 0 2588 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_4_1
timestamp 1607319584
transform 1 0 2596 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_557
timestamp 1607319584
transform 1 0 2604 0 1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_378
timestamp 1607319584
transform 1 0 2700 0 1 4305
box -2 -3 26 103
use MUX2X1  MUX2X1_227
timestamp 1607319584
transform -1 0 2772 0 1 4305
box -2 -3 50 103
use NAND2X1  NAND2X1_162
timestamp 1607319584
transform 1 0 2772 0 1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_169
timestamp 1607319584
transform -1 0 2820 0 1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_135
timestamp 1607319584
transform -1 0 2852 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_257
timestamp 1607319584
transform 1 0 2852 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_376
timestamp 1607319584
transform 1 0 2876 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_531
timestamp 1607319584
transform -1 0 2996 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_302
timestamp 1607319584
transform 1 0 2996 0 1 4305
box -2 -3 98 103
use FILL  FILL_43_5_0
timestamp 1607319584
transform -1 0 3100 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_5_1
timestamp 1607319584
transform -1 0 3108 0 1 4305
box -2 -3 10 103
use NAND2X1  NAND2X1_567
timestamp 1607319584
transform -1 0 3132 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_671
timestamp 1607319584
transform -1 0 3164 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1096
timestamp 1607319584
transform 1 0 3164 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_308
timestamp 1607319584
transform -1 0 3212 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_885
timestamp 1607319584
transform -1 0 3308 0 1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_568
timestamp 1607319584
transform 1 0 3308 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_318
timestamp 1607319584
transform -1 0 3428 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1660
timestamp 1607319584
transform -1 0 3460 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1661
timestamp 1607319584
transform -1 0 3492 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1607319584
transform 1 0 3492 0 1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_690
timestamp 1607319584
transform 1 0 3588 0 1 4305
box -2 -3 26 103
use FILL  FILL_43_6_0
timestamp 1607319584
transform 1 0 3612 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_6_1
timestamp 1607319584
transform 1 0 3620 0 1 4305
box -2 -3 10 103
use NAND2X1  NAND2X1_691
timestamp 1607319584
transform 1 0 3628 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_637
timestamp 1607319584
transform 1 0 3652 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_319
timestamp 1607319584
transform -1 0 3772 0 1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_430
timestamp 1607319584
transform 1 0 3772 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1607319584
transform 1 0 3796 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1392
timestamp 1607319584
transform 1 0 3892 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1391
timestamp 1607319584
transform -1 0 3956 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_449
timestamp 1607319584
transform -1 0 3972 0 1 4305
box -2 -3 18 103
use BUFX4  BUFX4_167
timestamp 1607319584
transform 1 0 3972 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_421
timestamp 1607319584
transform 1 0 4004 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_283
timestamp 1607319584
transform 1 0 4028 0 1 4305
box -2 -3 26 103
use BUFX4  BUFX4_464
timestamp 1607319584
transform 1 0 4052 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1343
timestamp 1607319584
transform -1 0 4116 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_7_0
timestamp 1607319584
transform -1 0 4124 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_7_1
timestamp 1607319584
transform -1 0 4132 0 1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_1344
timestamp 1607319584
transform -1 0 4164 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1607319584
transform -1 0 4260 0 1 4305
box -2 -3 98 103
use BUFX4  BUFX4_465
timestamp 1607319584
transform 1 0 4260 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1046
timestamp 1607319584
transform -1 0 4324 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_345
timestamp 1607319584
transform 1 0 4324 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1365
timestamp 1607319584
transform -1 0 4380 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_258
timestamp 1607319584
transform -1 0 4396 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1607319584
transform -1 0 4492 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_823
timestamp 1607319584
transform -1 0 4524 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_129
timestamp 1607319584
transform -1 0 4540 0 1 4305
box -2 -3 18 103
use INVX1  INVX1_72
timestamp 1607319584
transform -1 0 4556 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_352
timestamp 1607319584
transform 1 0 4556 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_924
timestamp 1607319584
transform -1 0 4612 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_8_0
timestamp 1607319584
transform -1 0 4620 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_8_1
timestamp 1607319584
transform -1 0 4628 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_177
timestamp 1607319584
transform -1 0 4724 0 1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_1457
timestamp 1607319584
transform -1 0 4756 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1458
timestamp 1607319584
transform -1 0 4788 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1477
timestamp 1607319584
transform -1 0 4820 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1478
timestamp 1607319584
transform -1 0 4852 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1465
timestamp 1607319584
transform 1 0 4852 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1466
timestamp 1607319584
transform -1 0 4916 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_181
timestamp 1607319584
transform -1 0 5012 0 1 4305
box -2 -3 98 103
use INVX1  INVX1_37
timestamp 1607319584
transform -1 0 5028 0 1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_1329
timestamp 1607319584
transform 1 0 5028 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1330
timestamp 1607319584
transform -1 0 5092 0 1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1607319584
transform 1 0 5092 0 1 4305
box -2 -3 98 103
use FILL  FILL_44_1
timestamp 1607319584
transform 1 0 5188 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_896
timestamp 1607319584
transform 1 0 4 0 -1 4505
box -2 -3 98 103
use AOI21X1  AOI21X1_133
timestamp 1607319584
transform 1 0 100 0 -1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_165
timestamp 1607319584
transform -1 0 156 0 -1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_872
timestamp 1607319584
transform 1 0 156 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_667
timestamp 1607319584
transform 1 0 252 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_864
timestamp 1607319584
transform -1 0 380 0 -1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_154
timestamp 1607319584
transform 1 0 380 0 -1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_124
timestamp 1607319584
transform -1 0 436 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_165
timestamp 1607319584
transform -1 0 460 0 -1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_860
timestamp 1607319584
transform 1 0 460 0 -1 4505
box -2 -3 98 103
use FILL  FILL_44_0_0
timestamp 1607319584
transform 1 0 556 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_0_1
timestamp 1607319584
transform 1 0 564 0 -1 4505
box -2 -3 10 103
use OAI21X1  OAI21X1_649
timestamp 1607319584
transform 1 0 572 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_846
timestamp 1607319584
transform 1 0 604 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1029
timestamp 1607319584
transform 1 0 700 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_150
timestamp 1607319584
transform 1 0 732 0 -1 4505
box -2 -3 26 103
use INVX1  INVX1_4
timestamp 1607319584
transform -1 0 772 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_712
timestamp 1607319584
transform 1 0 772 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_528
timestamp 1607319584
transform 1 0 868 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_527
timestamp 1607319584
transform -1 0 932 0 -1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_8
timestamp 1607319584
transform 1 0 932 0 -1 4505
box -2 -3 50 103
use OAI21X1  OAI21X1_1221
timestamp 1607319584
transform 1 0 980 0 -1 4505
box -2 -3 34 103
use BUFX4  BUFX4_456
timestamp 1607319584
transform -1 0 1044 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_1_0
timestamp 1607319584
transform -1 0 1052 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_1_1
timestamp 1607319584
transform -1 0 1060 0 -1 4505
box -2 -3 10 103
use INVX8  INVX8_10
timestamp 1607319584
transform -1 0 1100 0 -1 4505
box -2 -3 42 103
use OAI21X1  OAI21X1_513
timestamp 1607319584
transform 1 0 1100 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_514
timestamp 1607319584
transform -1 0 1164 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_59
timestamp 1607319584
transform 1 0 1164 0 -1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_61
timestamp 1607319584
transform 1 0 1188 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_268
timestamp 1607319584
transform -1 0 1244 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_548
timestamp 1607319584
transform 1 0 1244 0 -1 4505
box -2 -3 98 103
use INVX1  INVX1_223
timestamp 1607319584
transform 1 0 1340 0 -1 4505
box -2 -3 18 103
use CLKBUF1  CLKBUF1_82
timestamp 1607319584
transform -1 0 1428 0 -1 4505
box -2 -3 74 103
use MUX2X1  MUX2X1_68
timestamp 1607319584
transform 1 0 1428 0 -1 4505
box -2 -3 50 103
use OAI21X1  OAI21X1_884
timestamp 1607319584
transform -1 0 1508 0 -1 4505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_57
timestamp 1607319584
transform 1 0 1508 0 -1 4505
box -2 -3 74 103
use FILL  FILL_44_2_0
timestamp 1607319584
transform 1 0 1580 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_2_1
timestamp 1607319584
transform 1 0 1588 0 -1 4505
box -2 -3 10 103
use NAND2X1  NAND2X1_65
timestamp 1607319584
transform 1 0 1596 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_290
timestamp 1607319584
transform 1 0 1620 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_569
timestamp 1607319584
transform 1 0 1652 0 -1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_49
timestamp 1607319584
transform 1 0 1748 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1265
timestamp 1607319584
transform -1 0 1804 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_480
timestamp 1607319584
transform 1 0 1804 0 -1 4505
box -2 -3 18 103
use NAND2X1  NAND2X1_720
timestamp 1607319584
transform -1 0 1844 0 -1 4505
box -2 -3 26 103
use MUX2X1  MUX2X1_322
timestamp 1607319584
transform 1 0 1844 0 -1 4505
box -2 -3 50 103
use OAI21X1  OAI21X1_1222
timestamp 1607319584
transform -1 0 1924 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_255
timestamp 1607319584
transform -1 0 1956 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_882
timestamp 1607319584
transform 1 0 1956 0 -1 4505
box -2 -3 34 103
use MUX2X1  MUX2X1_67
timestamp 1607319584
transform -1 0 2036 0 -1 4505
box -2 -3 50 103
use CLKBUF1  CLKBUF1_41
timestamp 1607319584
transform 1 0 2036 0 -1 4505
box -2 -3 74 103
use FILL  FILL_44_3_0
timestamp 1607319584
transform 1 0 2108 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_3_1
timestamp 1607319584
transform 1 0 2116 0 -1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_526
timestamp 1607319584
transform 1 0 2124 0 -1 4505
box -2 -3 98 103
use NAND2X1  NAND2X1_48
timestamp 1607319584
transform -1 0 2244 0 -1 4505
box -2 -3 26 103
use MUX2X1  MUX2X1_226
timestamp 1607319584
transform 1 0 2244 0 -1 4505
box -2 -3 50 103
use OAI21X1  OAI21X1_881
timestamp 1607319584
transform 1 0 2292 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_306
timestamp 1607319584
transform -1 0 2348 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_967
timestamp 1607319584
transform -1 0 2380 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_349
timestamp 1607319584
transform -1 0 2396 0 -1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_243
timestamp 1607319584
transform -1 0 2428 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_244
timestamp 1607319584
transform -1 0 2460 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_659
timestamp 1607319584
transform -1 0 2492 0 -1 4505
box -2 -3 34 103
use BUFX4  BUFX4_435
timestamp 1607319584
transform 1 0 2492 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_434
timestamp 1607319584
transform -1 0 2540 0 -1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_297
timestamp 1607319584
transform 1 0 2540 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_4_0
timestamp 1607319584
transform 1 0 2572 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_4_1
timestamp 1607319584
transform 1 0 2580 0 -1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_855
timestamp 1607319584
transform 1 0 2588 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1073
timestamp 1607319584
transform 1 0 2684 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_513
timestamp 1607319584
transform -1 0 2740 0 -1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_54
timestamp 1607319584
transform 1 0 2740 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_261
timestamp 1607319584
transform -1 0 2796 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_664
timestamp 1607319584
transform -1 0 2828 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_286
timestamp 1607319584
transform -1 0 2844 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_533
timestamp 1607319584
transform -1 0 2940 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1095
timestamp 1607319584
transform 1 0 2940 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_947
timestamp 1607319584
transform 1 0 2972 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_889
timestamp 1607319584
transform -1 0 3100 0 -1 4505
box -2 -3 98 103
use FILL  FILL_44_5_0
timestamp 1607319584
transform -1 0 3108 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_5_1
timestamp 1607319584
transform -1 0 3116 0 -1 4505
box -2 -3 10 103
use OAI21X1  OAI21X1_945
timestamp 1607319584
transform -1 0 3148 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_157
timestamp 1607319584
transform -1 0 3164 0 -1 4505
box -2 -3 18 103
use BUFX4  BUFX4_82
timestamp 1607319584
transform -1 0 3196 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_50
timestamp 1607319584
transform 1 0 3196 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_257
timestamp 1607319584
transform -1 0 3252 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_834
timestamp 1607319584
transform 1 0 3252 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_46
timestamp 1607319584
transform -1 0 3300 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_529
timestamp 1607319584
transform -1 0 3396 0 -1 4505
box -2 -3 98 103
use INVX1  INVX1_336
timestamp 1607319584
transform 1 0 3396 0 -1 4505
box -2 -3 18 103
use CLKBUF1  CLKBUF1_53
timestamp 1607319584
transform 1 0 3412 0 -1 4505
box -2 -3 74 103
use NAND2X1  NAND2X1_361
timestamp 1607319584
transform 1 0 3484 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_968
timestamp 1607319584
transform -1 0 3540 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1654
timestamp 1607319584
transform 1 0 3540 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1655
timestamp 1607319584
transform -1 0 3604 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_6_0
timestamp 1607319584
transform 1 0 3604 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_6_1
timestamp 1607319584
transform 1 0 3612 0 -1 4505
box -2 -3 10 103
use INVX1  INVX1_400
timestamp 1607319584
transform 1 0 3620 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_315
timestamp 1607319584
transform 1 0 3636 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1657
timestamp 1607319584
transform 1 0 3732 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_208
timestamp 1607319584
transform 1 0 3764 0 -1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_1656
timestamp 1607319584
transform -1 0 3812 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1662
timestamp 1607319584
transform 1 0 3812 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1663
timestamp 1607319584
transform -1 0 3876 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_824
timestamp 1607319584
transform -1 0 3908 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_794
timestamp 1607319584
transform -1 0 3932 0 -1 4505
box -2 -3 26 103
use INVX1  INVX1_321
timestamp 1607319584
transform -1 0 3948 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1607319584
transform -1 0 4044 0 -1 4505
box -2 -3 98 103
use MUX2X1  MUX2X1_142
timestamp 1607319584
transform 1 0 4044 0 -1 4505
box -2 -3 50 103
use BUFX4  BUFX4_460
timestamp 1607319584
transform 1 0 4092 0 -1 4505
box -2 -3 34 103
use FILL  FILL_44_7_0
timestamp 1607319584
transform 1 0 4124 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_7_1
timestamp 1607319584
transform 1 0 4132 0 -1 4505
box -2 -3 10 103
use OAI21X1  OAI21X1_1382
timestamp 1607319584
transform 1 0 4140 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1607319584
transform 1 0 4172 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1381
timestamp 1607319584
transform -1 0 4300 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1607319584
transform 1 0 4300 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1338
timestamp 1607319584
transform 1 0 4396 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1337
timestamp 1607319584
transform -1 0 4460 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1476
timestamp 1607319584
transform 1 0 4460 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1475
timestamp 1607319584
transform -1 0 4524 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_186
timestamp 1607319584
transform -1 0 4620 0 -1 4505
box -2 -3 98 103
use INVX1  INVX1_136
timestamp 1607319584
transform -1 0 4636 0 -1 4505
box -2 -3 18 103
use FILL  FILL_44_8_0
timestamp 1607319584
transform -1 0 4644 0 -1 4505
box -2 -3 10 103
use FILL  FILL_44_8_1
timestamp 1607319584
transform -1 0 4652 0 -1 4505
box -2 -3 10 103
use NAND2X1  NAND2X1_796
timestamp 1607319584
transform -1 0 4676 0 -1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1459
timestamp 1607319584
transform -1 0 4708 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1460
timestamp 1607319584
transform -1 0 4740 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1180
timestamp 1607319584
transform -1 0 4772 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_392
timestamp 1607319584
transform -1 0 4788 0 -1 4505
box -2 -3 18 103
use BUFX4  BUFX4_393
timestamp 1607319584
transform -1 0 4820 0 -1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_167
timestamp 1607319584
transform 1 0 4820 0 -1 4505
box -2 -3 26 103
use BUFX4  BUFX4_392
timestamp 1607319584
transform 1 0 4844 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1333
timestamp 1607319584
transform 1 0 4876 0 -1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1334
timestamp 1607319584
transform -1 0 4940 0 -1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1607319584
transform -1 0 5036 0 -1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_669
timestamp 1607319584
transform -1 0 5068 0 -1 4505
box -2 -3 34 103
use INVX1  INVX1_180
timestamp 1607319584
transform -1 0 5084 0 -1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_883
timestamp 1607319584
transform 1 0 5084 0 -1 4505
box -2 -3 98 103
use FILL  FILL_45_1
timestamp 1607319584
transform -1 0 5188 0 -1 4505
box -2 -3 10 103
use FILL  FILL_45_2
timestamp 1607319584
transform -1 0 5196 0 -1 4505
box -2 -3 10 103
use NOR2X1  NOR2X1_176
timestamp 1607319584
transform -1 0 28 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_142
timestamp 1607319584
transform -1 0 60 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_880
timestamp 1607319584
transform 1 0 60 0 1 4505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_878
timestamp 1607319584
transform 1 0 4 0 -1 4705
box -2 -3 98 103
use AOI21X1  AOI21X1_131
timestamp 1607319584
transform 1 0 100 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_868
timestamp 1607319584
transform 1 0 156 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_163
timestamp 1607319584
transform 1 0 132 0 -1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_838
timestamp 1607319584
transform 1 0 156 0 -1 4705
box -2 -3 98 103
use INVX1  INVX1_243
timestamp 1607319584
transform 1 0 252 0 1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_663
timestamp 1607319584
transform 1 0 268 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_161
timestamp 1607319584
transform -1 0 324 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_633
timestamp 1607319584
transform 1 0 252 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_632
timestamp 1607319584
transform -1 0 316 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_624
timestamp 1607319584
transform 1 0 324 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_625
timestamp 1607319584
transform -1 0 388 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_834
timestamp 1607319584
transform 1 0 388 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_653
timestamp 1607319584
transform 1 0 316 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_652
timestamp 1607319584
transform -1 0 380 0 -1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_129
timestamp 1607319584
transform 1 0 380 0 -1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_120
timestamp 1607319584
transform 1 0 484 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_161
timestamp 1607319584
transform -1 0 436 0 -1 4705
box -2 -3 26 103
use BUFX4  BUFX4_120
timestamp 1607319584
transform -1 0 468 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_241
timestamp 1607319584
transform 1 0 468 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_1031
timestamp 1607319584
transform 1 0 484 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_150
timestamp 1607319584
transform -1 0 540 0 1 4505
box -2 -3 26 103
use FILL  FILL_45_0_0
timestamp 1607319584
transform 1 0 540 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_0_1
timestamp 1607319584
transform 1 0 548 0 1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_833
timestamp 1607319584
transform 1 0 556 0 1 4505
box -2 -3 98 103
use NAND2X1  NAND2X1_467
timestamp 1607319584
transform -1 0 540 0 -1 4705
box -2 -3 26 103
use FILL  FILL_46_0_0
timestamp 1607319584
transform 1 0 540 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_0_1
timestamp 1607319584
transform 1 0 548 0 -1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_842
timestamp 1607319584
transform 1 0 556 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_640
timestamp 1607319584
transform -1 0 684 0 1 4505
box -2 -3 34 103
use BUFX4  BUFX4_119
timestamp 1607319584
transform 1 0 684 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_641
timestamp 1607319584
transform 1 0 652 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_369
timestamp 1607319584
transform 1 0 684 0 -1 4705
box -2 -3 18 103
use MUX2X1  MUX2X1_179
timestamp 1607319584
transform 1 0 700 0 -1 4705
box -2 -3 50 103
use NAND2X1  NAND2X1_465
timestamp 1607319584
transform -1 0 740 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_622
timestamp 1607319584
transform 1 0 740 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_623
timestamp 1607319584
transform -1 0 804 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_626
timestamp 1607319584
transform 1 0 804 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1032
timestamp 1607319584
transform 1 0 748 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_433
timestamp 1607319584
transform 1 0 780 0 -1 4705
box -2 -3 18 103
use INVX1  INVX1_305
timestamp 1607319584
transform 1 0 796 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_627
timestamp 1607319584
transform -1 0 868 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_835
timestamp 1607319584
transform 1 0 868 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_639
timestamp 1607319584
transform 1 0 812 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_638
timestamp 1607319584
transform 1 0 844 0 -1 4705
box -2 -3 34 103
use BUFX4  BUFX4_121
timestamp 1607319584
transform -1 0 908 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_841
timestamp 1607319584
transform 1 0 908 0 -1 4705
box -2 -3 98 103
use NAND2X1  NAND2X1_672
timestamp 1607319584
transform -1 0 988 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_720
timestamp 1607319584
transform -1 0 1084 0 1 4505
box -2 -3 98 103
use NAND2X1  NAND2X1_468
timestamp 1607319584
transform -1 0 1028 0 -1 4705
box -2 -3 26 103
use FILL  FILL_45_1_0
timestamp 1607319584
transform 1 0 1084 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_1_1
timestamp 1607319584
transform 1 0 1092 0 1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_705
timestamp 1607319584
transform 1 0 1100 0 1 4505
box -2 -3 98 103
use FILL  FILL_46_1_0
timestamp 1607319584
transform 1 0 1028 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_1_1
timestamp 1607319584
transform 1 0 1036 0 -1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_546
timestamp 1607319584
transform 1 0 1044 0 -1 4705
box -2 -3 98 103
use NAND2X1  NAND2X1_534
timestamp 1607319584
transform -1 0 1220 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_42
timestamp 1607319584
transform 1 0 1140 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_54
timestamp 1607319584
transform 1 0 1172 0 -1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_266
timestamp 1607319584
transform -1 0 1228 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1093
timestamp 1607319584
transform 1 0 1220 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_859
timestamp 1607319584
transform 1 0 1252 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_95
timestamp 1607319584
transform 1 0 1228 0 -1 4705
box -2 -3 18 103
use AOI21X1  AOI21X1_44
timestamp 1607319584
transform 1 0 1244 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_56
timestamp 1607319584
transform 1 0 1276 0 -1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_883
timestamp 1607319584
transform 1 0 1300 0 -1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_119
timestamp 1607319584
transform 1 0 1348 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_149
timestamp 1607319584
transform -1 0 1404 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_309
timestamp 1607319584
transform 1 0 1404 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_892
timestamp 1607319584
transform -1 0 1428 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_291
timestamp 1607319584
transform -1 0 1460 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_540
timestamp 1607319584
transform 1 0 1460 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_292
timestamp 1607319584
transform -1 0 1460 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_572
timestamp 1607319584
transform 1 0 1460 0 -1 4705
box -2 -3 98 103
use FILL  FILL_45_2_0
timestamp 1607319584
transform -1 0 1564 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_2_1
timestamp 1607319584
transform -1 0 1572 0 1 4505
box -2 -3 10 103
use INVX1  INVX1_96
timestamp 1607319584
transform -1 0 1588 0 1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_295
timestamp 1607319584
transform -1 0 1620 0 1 4505
box -2 -3 34 103
use FILL  FILL_46_2_0
timestamp 1607319584
transform 1 0 1556 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_2_1
timestamp 1607319584
transform 1 0 1564 0 -1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_296
timestamp 1607319584
transform 1 0 1572 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_272
timestamp 1607319584
transform -1 0 1636 0 -1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_36
timestamp 1607319584
transform 1 0 1620 0 1 4505
box -2 -3 34 103
use NOR2X1  NOR2X1_46
timestamp 1607319584
transform 1 0 1652 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_543
timestamp 1607319584
transform 1 0 1676 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_479
timestamp 1607319584
transform 1 0 1636 0 -1 4705
box -2 -3 18 103
use INVX1  INVX1_221
timestamp 1607319584
transform 1 0 1652 0 -1 4705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_568
timestamp 1607319584
transform 1 0 1668 0 -1 4705
box -2 -3 98 103
use AOI21X1  AOI21X1_39
timestamp 1607319584
transform -1 0 1804 0 1 4505
box -2 -3 34 103
use INVX1  INVX1_477
timestamp 1607319584
transform -1 0 1820 0 1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_528
timestamp 1607319584
transform -1 0 1916 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_288
timestamp 1607319584
transform 1 0 1764 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_287
timestamp 1607319584
transform -1 0 1828 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_256
timestamp 1607319584
transform 1 0 1916 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_520
timestamp 1607319584
transform -1 0 1924 0 -1 4705
box -2 -3 98 103
use NAND2X1  NAND2X1_535
timestamp 1607319584
transform -1 0 1972 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_307
timestamp 1607319584
transform 1 0 1972 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_875
timestamp 1607319584
transform 1 0 1996 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_239
timestamp 1607319584
transform -1 0 1956 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_240
timestamp 1607319584
transform -1 0 1988 0 -1 4705
box -2 -3 34 103
use BUFX4  BUFX4_434
timestamp 1607319584
transform -1 0 2020 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_44
timestamp 1607319584
transform 1 0 2020 0 -1 4705
box -2 -3 26 103
use FILL  FILL_45_3_0
timestamp 1607319584
transform -1 0 2100 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_3_1
timestamp 1607319584
transform -1 0 2108 0 1 4505
box -2 -3 10 103
use AOI21X1  AOI21X1_128
timestamp 1607319584
transform -1 0 2140 0 1 4505
box -2 -3 34 103
use AOI21X1  AOI21X1_34
timestamp 1607319584
transform -1 0 2076 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_3_0
timestamp 1607319584
transform -1 0 2084 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_3_1
timestamp 1607319584
transform -1 0 2092 0 -1 4705
box -2 -3 10 103
use BUFX4  BUFX4_165
timestamp 1607319584
transform -1 0 2124 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_853
timestamp 1607319584
transform 1 0 2124 0 -1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_160
timestamp 1607319584
transform 1 0 2140 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_398
timestamp 1607319584
transform -1 0 2188 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1094
timestamp 1607319584
transform -1 0 2220 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_155
timestamp 1607319584
transform -1 0 2244 0 1 4505
box -2 -3 26 103
use INVX1  INVX1_306
timestamp 1607319584
transform 1 0 2220 0 -1 4705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_522
timestamp 1607319584
transform 1 0 2244 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_657
timestamp 1607319584
transform -1 0 2268 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_48
timestamp 1607319584
transform 1 0 2268 0 -1 4705
box -2 -3 18 103
use INVX1  INVX1_93
timestamp 1607319584
transform 1 0 2284 0 -1 4705
box -2 -3 18 103
use BUFX4  BUFX4_437
timestamp 1607319584
transform 1 0 2300 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_179
timestamp 1607319584
transform 1 0 2340 0 1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_867
timestamp 1607319584
transform -1 0 2452 0 1 4505
box -2 -3 98 103
use BUFX4  BUFX4_436
timestamp 1607319584
transform 1 0 2332 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_235
timestamp 1607319584
transform 1 0 2364 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_236
timestamp 1607319584
transform -1 0 2428 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_662
timestamp 1607319584
transform 1 0 2452 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_160
timestamp 1607319584
transform -1 0 2508 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_514
timestamp 1607319584
transform 1 0 2508 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_518
timestamp 1607319584
transform -1 0 2524 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_249
timestamp 1607319584
transform 1 0 2524 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_298
timestamp 1607319584
transform 1 0 2532 0 1 4505
box -2 -3 34 103
use FILL  FILL_45_4_0
timestamp 1607319584
transform 1 0 2564 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_4_1
timestamp 1607319584
transform 1 0 2572 0 1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_573
timestamp 1607319584
transform 1 0 2580 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_250
timestamp 1607319584
transform -1 0 2588 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_4_0
timestamp 1607319584
transform 1 0 2588 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_4_1
timestamp 1607319584
transform 1 0 2596 0 -1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_525
timestamp 1607319584
transform 1 0 2604 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_294
timestamp 1607319584
transform 1 0 2676 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_293
timestamp 1607319584
transform 1 0 2708 0 1 4505
box -2 -3 34 103
use INVX1  INVX1_285
timestamp 1607319584
transform -1 0 2716 0 -1 4705
box -2 -3 18 103
use AOI21X1  AOI21X1_130
timestamp 1607319584
transform 1 0 2716 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_571
timestamp 1607319584
transform -1 0 2836 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_162
timestamp 1607319584
transform -1 0 2772 0 -1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_877
timestamp 1607319584
transform 1 0 2772 0 -1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_869
timestamp 1607319584
transform 1 0 2836 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_307
timestamp 1607319584
transform 1 0 2932 0 1 4505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_547
timestamp 1607319584
transform 1 0 2868 0 -1 4705
box -2 -3 98 103
use NAND2X1  NAND2X1_536
timestamp 1607319584
transform -1 0 2972 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_60
timestamp 1607319584
transform 1 0 2972 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_377
timestamp 1607319584
transform 1 0 2996 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_246
timestamp 1607319584
transform 1 0 3020 0 1 4505
box -2 -3 34 103
use INVX1  INVX1_159
timestamp 1607319584
transform 1 0 2964 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_267
timestamp 1607319584
transform 1 0 2980 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_833
timestamp 1607319584
transform 1 0 3012 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_241
timestamp 1607319584
transform -1 0 3100 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_255
timestamp 1607319584
transform -1 0 3068 0 -1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_245
timestamp 1607319584
transform -1 0 3084 0 1 4505
box -2 -3 34 103
use FILL  FILL_46_5_0
timestamp 1607319584
transform -1 0 3108 0 -1 4705
box -2 -3 10 103
use NAND2X1  NAND2X1_375
timestamp 1607319584
transform -1 0 3108 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_242
timestamp 1607319584
transform -1 0 3148 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_5_1
timestamp 1607319584
transform -1 0 3116 0 -1 4705
box -2 -3 10 103
use NOR2X1  NOR2X1_53
timestamp 1607319584
transform 1 0 3124 0 1 4505
box -2 -3 26 103
use FILL  FILL_45_5_1
timestamp 1607319584
transform 1 0 3116 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_5_0
timestamp 1607319584
transform 1 0 3108 0 1 4505
box -2 -3 10 103
use AOI21X1  AOI21X1_41
timestamp 1607319584
transform -1 0 3180 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_553
timestamp 1607319584
transform -1 0 3276 0 1 4505
box -2 -3 98 103
use NOR2X1  NOR2X1_55
timestamp 1607319584
transform 1 0 3148 0 -1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_43
timestamp 1607319584
transform -1 0 3204 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_537
timestamp 1607319584
transform 1 0 3204 0 -1 4705
box -2 -3 98 103
use NAND2X1  NAND2X1_256
timestamp 1607319584
transform -1 0 3300 0 1 4505
box -2 -3 26 103
use NAND2X1  NAND2X1_537
timestamp 1607319584
transform -1 0 3324 0 1 4505
box -2 -3 26 103
use AOI21X1  AOI21X1_35
timestamp 1607319584
transform 1 0 3324 0 1 4505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_11
timestamp 1607319584
transform -1 0 3372 0 -1 4705
box -2 -3 74 103
use NOR2X1  NOR2X1_45
timestamp 1607319584
transform -1 0 3380 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_539
timestamp 1607319584
transform 1 0 3380 0 1 4505
box -2 -3 98 103
use AOI21X1  AOI21X1_137
timestamp 1607319584
transform 1 0 3372 0 -1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_171
timestamp 1607319584
transform -1 0 3428 0 -1 4705
box -2 -3 26 103
use INVX1  INVX1_144
timestamp 1607319584
transform 1 0 3428 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_932
timestamp 1607319584
transform 1 0 3476 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_399
timestamp 1607319584
transform -1 0 3532 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_312
timestamp 1607319584
transform -1 0 3628 0 1 4505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_891
timestamp 1607319584
transform 1 0 3444 0 -1 4705
box -2 -3 98 103
use FILL  FILL_45_6_0
timestamp 1607319584
transform -1 0 3636 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_6_1
timestamp 1607319584
transform -1 0 3644 0 1 4505
box -2 -3 10 103
use INVX1  INVX1_68
timestamp 1607319584
transform -1 0 3556 0 -1 4705
box -2 -3 18 103
use BUFX4  BUFX4_168
timestamp 1607319584
transform 1 0 3556 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1648
timestamp 1607319584
transform -1 0 3620 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_6_0
timestamp 1607319584
transform 1 0 3620 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_6_1
timestamp 1607319584
transform 1 0 3628 0 -1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_1640
timestamp 1607319584
transform 1 0 3636 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1649
timestamp 1607319584
transform -1 0 3676 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_316
timestamp 1607319584
transform 1 0 3676 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1641
timestamp 1607319584
transform -1 0 3700 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_308
timestamp 1607319584
transform 1 0 3700 0 -1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1607319584
transform 1 0 3772 0 1 4505
box -2 -3 98 103
use INVX1  INVX1_196
timestamp 1607319584
transform -1 0 3812 0 -1 4705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1607319584
transform -1 0 3908 0 -1 4705
box -2 -3 98 103
use INVX1  INVX1_38
timestamp 1607319584
transform 1 0 3868 0 1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_1361
timestamp 1607319584
transform 1 0 3884 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1339
timestamp 1607319584
transform 1 0 3916 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1359
timestamp 1607319584
transform -1 0 3940 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1360
timestamp 1607319584
transform -1 0 3972 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1340
timestamp 1607319584
transform -1 0 3980 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1335
timestamp 1607319584
transform 1 0 3980 0 1 4505
box -2 -3 34 103
use INVX1  INVX1_193
timestamp 1607319584
transform 1 0 4012 0 1 4505
box -2 -3 18 103
use OAI21X1  OAI21X1_981
timestamp 1607319584
transform 1 0 4028 0 1 4505
box -2 -3 34 103
use BUFX4  BUFX4_468
timestamp 1607319584
transform -1 0 4004 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1377
timestamp 1607319584
transform 1 0 4004 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1378
timestamp 1607319584
transform -1 0 4068 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1389
timestamp 1607319584
transform -1 0 4116 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_260
timestamp 1607319584
transform -1 0 4084 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_1336
timestamp 1607319584
transform -1 0 4116 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_414
timestamp 1607319584
transform 1 0 4060 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1351
timestamp 1607319584
transform -1 0 4164 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_7_1
timestamp 1607319584
transform -1 0 4132 0 -1 4705
box -2 -3 10 103
use FILL  FILL_46_7_0
timestamp 1607319584
transform -1 0 4124 0 -1 4705
box -2 -3 10 103
use FILL  FILL_45_7_1
timestamp 1607319584
transform -1 0 4132 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_7_0
timestamp 1607319584
transform -1 0 4124 0 1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1607319584
transform -1 0 4228 0 1 4505
box -2 -3 98 103
use NAND2X1  NAND2X1_483
timestamp 1607319584
transform 1 0 4228 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1352
timestamp 1607319584
transform -1 0 4196 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1607319584
transform -1 0 4292 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1045
timestamp 1607319584
transform -1 0 4284 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_484
timestamp 1607319584
transform -1 0 4308 0 1 4505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_17
timestamp 1607319584
transform -1 0 4380 0 1 4505
box -2 -3 74 103
use OAI21X1  OAI21X1_1353
timestamp 1607319584
transform -1 0 4324 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1354
timestamp 1607319584
transform -1 0 4356 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_257
timestamp 1607319584
transform -1 0 4396 0 1 4505
box -2 -3 18 103
use NAND2X1  NAND2X1_697
timestamp 1607319584
transform 1 0 4396 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1244
timestamp 1607319584
transform 1 0 4420 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1349
timestamp 1607319584
transform -1 0 4388 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1350
timestamp 1607319584
transform -1 0 4420 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_456
timestamp 1607319584
transform 1 0 4420 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_1345
timestamp 1607319584
transform 1 0 4436 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_239
timestamp 1607319584
transform 1 0 4452 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1116
timestamp 1607319584
transform -1 0 4508 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_918
timestamp 1607319584
transform 1 0 4508 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_559
timestamp 1607319584
transform 1 0 4540 0 1 4505
box -2 -3 26 103
use OAI21X1  OAI21X1_1346
timestamp 1607319584
transform -1 0 4500 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_328
timestamp 1607319584
transform -1 0 4516 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_1468
timestamp 1607319584
transform 1 0 4516 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1467
timestamp 1607319584
transform -1 0 4580 0 -1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_346
timestamp 1607319584
transform 1 0 4564 0 1 4505
box -2 -3 26 103
use INVX1  INVX1_200
timestamp 1607319584
transform -1 0 4604 0 1 4505
box -2 -3 18 103
use FILL  FILL_45_8_0
timestamp 1607319584
transform -1 0 4612 0 1 4505
box -2 -3 10 103
use FILL  FILL_45_8_1
timestamp 1607319584
transform -1 0 4620 0 1 4505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_178
timestamp 1607319584
transform -1 0 4716 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1363
timestamp 1607319584
transform 1 0 4580 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1461
timestamp 1607319584
transform -1 0 4644 0 -1 4705
box -2 -3 34 103
use FILL  FILL_46_8_0
timestamp 1607319584
transform -1 0 4652 0 -1 4705
box -2 -3 10 103
use NAND2X1  NAND2X1_628
timestamp 1607319584
transform 1 0 4716 0 1 4505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_180
timestamp 1607319584
transform -1 0 4836 0 1 4505
box -2 -3 98 103
use FILL  FILL_46_8_1
timestamp 1607319584
transform -1 0 4660 0 -1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_1471
timestamp 1607319584
transform -1 0 4692 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_982
timestamp 1607319584
transform -1 0 4724 0 -1 4705
box -2 -3 34 103
use INVX1  INVX1_194
timestamp 1607319584
transform 1 0 4724 0 -1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_1364
timestamp 1607319584
transform 1 0 4740 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1464
timestamp 1607319584
transform -1 0 4868 0 1 4505
box -2 -3 34 103
use NAND2X1  NAND2X1_797
timestamp 1607319584
transform 1 0 4772 0 -1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_1463
timestamp 1607319584
transform -1 0 4828 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1480
timestamp 1607319584
transform 1 0 4828 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1485
timestamp 1607319584
transform 1 0 4868 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1486
timestamp 1607319584
transform -1 0 4932 0 1 4505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_191
timestamp 1607319584
transform -1 0 5028 0 1 4505
box -2 -3 98 103
use OAI21X1  OAI21X1_1479
timestamp 1607319584
transform -1 0 4892 0 -1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_188
timestamp 1607319584
transform -1 0 4988 0 -1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1487
timestamp 1607319584
transform 1 0 5028 0 1 4505
box -2 -3 34 103
use OAI21X1  OAI21X1_1469
timestamp 1607319584
transform 1 0 4988 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1483
timestamp 1607319584
transform 1 0 5020 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1484
timestamp 1607319584
transform 1 0 5052 0 -1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1488
timestamp 1607319584
transform -1 0 5092 0 1 4505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_84
timestamp 1607319584
transform -1 0 5164 0 1 4505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_190
timestamp 1607319584
transform -1 0 5180 0 -1 4705
box -2 -3 98 103
use NAND2X1  NAND2X1_184
timestamp 1607319584
transform -1 0 5188 0 1 4505
box -2 -3 26 103
use FILL  FILL_46_1
timestamp 1607319584
transform 1 0 5188 0 1 4505
box -2 -3 10 103
use FILL  FILL_47_1
timestamp 1607319584
transform -1 0 5188 0 -1 4705
box -2 -3 10 103
use FILL  FILL_47_2
timestamp 1607319584
transform -1 0 5196 0 -1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_840
timestamp 1607319584
transform 1 0 4 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_637
timestamp 1607319584
transform 1 0 100 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_636
timestamp 1607319584
transform -1 0 164 0 1 4705
box -2 -3 34 103
use INVX1  INVX1_497
timestamp 1607319584
transform 1 0 164 0 1 4705
box -2 -3 18 103
use OAI21X1  OAI21X1_628
timestamp 1607319584
transform 1 0 180 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_848
timestamp 1607319584
transform 1 0 212 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_647
timestamp 1607319584
transform 1 0 308 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_646
timestamp 1607319584
transform -1 0 372 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_876
timestamp 1607319584
transform 1 0 372 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_645
timestamp 1607319584
transform 1 0 468 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_644
timestamp 1607319584
transform -1 0 532 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_0_0
timestamp 1607319584
transform 1 0 532 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_0_1
timestamp 1607319584
transform 1 0 540 0 1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_634
timestamp 1607319584
transform 1 0 548 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_837
timestamp 1607319584
transform 1 0 580 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_631
timestamp 1607319584
transform 1 0 676 0 1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_168
timestamp 1607319584
transform -1 0 732 0 1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_630
timestamp 1607319584
transform -1 0 764 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_651
timestamp 1607319584
transform 1 0 764 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_650
timestamp 1607319584
transform 1 0 796 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_847
timestamp 1607319584
transform 1 0 828 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_554
timestamp 1607319584
transform 1 0 924 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_1_0
timestamp 1607319584
transform 1 0 1020 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_1_1
timestamp 1607319584
transform 1 0 1028 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_556
timestamp 1607319584
transform 1 0 1036 0 1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_172
timestamp 1607319584
transform 1 0 1132 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_138
timestamp 1607319584
transform -1 0 1188 0 1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_308
timestamp 1607319584
transform -1 0 1212 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_570
timestamp 1607319584
transform 1 0 1212 0 1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_151
timestamp 1607319584
transform -1 0 1332 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_121
timestamp 1607319584
transform -1 0 1364 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_552
timestamp 1607319584
transform 1 0 1364 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_562
timestamp 1607319584
transform 1 0 1460 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_2_0
timestamp 1607319584
transform -1 0 1564 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_2_1
timestamp 1607319584
transform -1 0 1572 0 1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_231
timestamp 1607319584
transform -1 0 1604 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_275
timestamp 1607319584
transform -1 0 1636 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_276
timestamp 1607319584
transform -1 0 1668 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_285
timestamp 1607319584
transform -1 0 1700 0 1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_673
timestamp 1607319584
transform -1 0 1724 0 1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_237
timestamp 1607319584
transform 1 0 1724 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_879
timestamp 1607319584
transform 1 0 1756 0 1 4705
box -2 -3 98 103
use AOI21X1  AOI21X1_132
timestamp 1607319584
transform 1 0 1852 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_164
timestamp 1607319584
transform -1 0 1908 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_538
timestamp 1607319584
transform 1 0 1908 0 1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_158
timestamp 1607319584
transform -1 0 2028 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_126
timestamp 1607319584
transform -1 0 2060 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_3_0
timestamp 1607319584
transform 1 0 2060 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_3_1
timestamp 1607319584
transform 1 0 2068 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_873
timestamp 1607319584
transform 1 0 2076 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_227
timestamp 1607319584
transform 1 0 2172 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_228
timestamp 1607319584
transform -1 0 2236 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_514
timestamp 1607319584
transform 1 0 2236 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_281
timestamp 1607319584
transform 1 0 2332 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_282
timestamp 1607319584
transform -1 0 2396 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_565
timestamp 1607319584
transform 1 0 2396 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_225
timestamp 1607319584
transform 1 0 2492 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1607319584
transform 1 0 2524 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_37
timestamp 1607319584
transform -1 0 2580 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_4_0
timestamp 1607319584
transform 1 0 2580 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_4_1
timestamp 1607319584
transform 1 0 2588 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_541
timestamp 1607319584
transform 1 0 2596 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_233
timestamp 1607319584
transform 1 0 2692 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_234
timestamp 1607319584
transform -1 0 2756 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_517
timestamp 1607319584
transform -1 0 2852 0 1 4705
box -2 -3 98 103
use INVX1  INVX1_45
timestamp 1607319584
transform 1 0 2852 0 1 4705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_523
timestamp 1607319584
transform 1 0 2868 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_521
timestamp 1607319584
transform 1 0 2964 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_5_0
timestamp 1607319584
transform -1 0 3068 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_5_1
timestamp 1607319584
transform -1 0 3076 0 1 4705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_555
timestamp 1607319584
transform -1 0 3172 0 1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_43
timestamp 1607319584
transform -1 0 3196 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_33
timestamp 1607319584
transform -1 0 3228 0 1 4705
box -2 -3 34 103
use AOI21X1  AOI21X1_139
timestamp 1607319584
transform 1 0 3228 0 1 4705
box -2 -3 34 103
use NOR2X1  NOR2X1_173
timestamp 1607319584
transform -1 0 3284 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_893
timestamp 1607319584
transform -1 0 3380 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1644
timestamp 1607319584
transform -1 0 3412 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1638
timestamp 1607319584
transform -1 0 3444 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1646
timestamp 1607319584
transform -1 0 3476 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1607319584
transform 1 0 3476 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1380
timestamp 1607319584
transform 1 0 3572 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_6_0
timestamp 1607319584
transform -1 0 3612 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_6_1
timestamp 1607319584
transform -1 0 3620 0 1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_1379
timestamp 1607319584
transform -1 0 3652 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1607319584
transform -1 0 3748 0 1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_307
timestamp 1607319584
transform 1 0 3748 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_246
timestamp 1607319584
transform -1 0 3804 0 1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_241
timestamp 1607319584
transform -1 0 3828 0 1 4705
box -2 -3 26 103
use OAI21X1  OAI21X1_1383
timestamp 1607319584
transform 1 0 3828 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1384
timestamp 1607319584
transform -1 0 3892 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1607319584
transform -1 0 3988 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1607319584
transform -1 0 4084 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1390
timestamp 1607319584
transform -1 0 4116 0 1 4705
box -2 -3 34 103
use FILL  FILL_47_7_0
timestamp 1607319584
transform 1 0 4116 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_7_1
timestamp 1607319584
transform 1 0 4124 0 1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_1385
timestamp 1607319584
transform 1 0 4132 0 1 4705
box -2 -3 34 103
use OAI21X1  OAI21X1_1386
timestamp 1607319584
transform -1 0 4196 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1607319584
transform -1 0 4292 0 1 4705
box -2 -3 98 103
use BUFX4  BUFX4_467
timestamp 1607319584
transform -1 0 4324 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1607319584
transform -1 0 4420 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1607319584
transform 1 0 4420 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1462
timestamp 1607319584
transform 1 0 4516 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_179
timestamp 1607319584
transform 1 0 4548 0 1 4705
box -2 -3 98 103
use FILL  FILL_47_8_0
timestamp 1607319584
transform -1 0 4652 0 1 4705
box -2 -3 10 103
use FILL  FILL_47_8_1
timestamp 1607319584
transform -1 0 4660 0 1 4705
box -2 -3 10 103
use OAI21X1  OAI21X1_1472
timestamp 1607319584
transform -1 0 4692 0 1 4705
box -2 -3 34 103
use NAND2X1  NAND2X1_415
timestamp 1607319584
transform -1 0 4716 0 1 4705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1607319584
transform -1 0 4812 0 1 4705
box -2 -3 98 103
use NOR2X1  NOR2X1_302
timestamp 1607319584
transform 1 0 4812 0 1 4705
box -2 -3 26 103
use AOI21X1  AOI21X1_241
timestamp 1607319584
transform -1 0 4868 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1607319584
transform -1 0 4964 0 1 4705
box -2 -3 98 103
use OAI21X1  OAI21X1_1470
timestamp 1607319584
transform 1 0 4964 0 1 4705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_183
timestamp 1607319584
transform -1 0 5092 0 1 4705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_192
timestamp 1607319584
transform -1 0 5188 0 1 4705
box -2 -3 98 103
use FILL  FILL_48_1
timestamp 1607319584
transform 1 0 5188 0 1 4705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_81
timestamp 1607319584
transform -1 0 76 0 -1 4905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_15
timestamp 1607319584
transform 1 0 76 0 -1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_836
timestamp 1607319584
transform -1 0 244 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_629
timestamp 1607319584
transform -1 0 276 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_845
timestamp 1607319584
transform 1 0 276 0 -1 4905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_7
timestamp 1607319584
transform 1 0 372 0 -1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_844
timestamp 1607319584
transform 1 0 444 0 -1 4905
box -2 -3 98 103
use FILL  FILL_48_0_0
timestamp 1607319584
transform -1 0 548 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_0_1
timestamp 1607319584
transform -1 0 556 0 -1 4905
box -2 -3 10 103
use OAI21X1  OAI21X1_635
timestamp 1607319584
transform -1 0 588 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_839
timestamp 1607319584
transform 1 0 588 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_670
timestamp 1607319584
transform 1 0 684 0 -1 4905
box -2 -3 34 103
use INVX1  INVX1_244
timestamp 1607319584
transform -1 0 732 0 -1 4905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_884
timestamp 1607319584
transform -1 0 828 0 -1 4905
box -2 -3 98 103
use NOR2X1  NOR2X1_147
timestamp 1607319584
transform -1 0 852 0 -1 4905
box -2 -3 26 103
use AOI21X1  AOI21X1_117
timestamp 1607319584
transform 1 0 852 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_857
timestamp 1607319584
transform 1 0 884 0 -1 4905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_95
timestamp 1607319584
transform 1 0 980 0 -1 4905
box -2 -3 74 103
use FILL  FILL_48_1_0
timestamp 1607319584
transform 1 0 1052 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_1_1
timestamp 1607319584
transform 1 0 1060 0 -1 4905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_46
timestamp 1607319584
transform 1 0 1068 0 -1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_863
timestamp 1607319584
transform 1 0 1140 0 -1 4905
box -2 -3 98 103
use AOI21X1  AOI21X1_123
timestamp 1607319584
transform 1 0 1236 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_153
timestamp 1607319584
transform 1 0 1268 0 -1 4905
box -2 -3 26 103
use BUFX4  BUFX4_18
timestamp 1607319584
transform 1 0 1292 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_861
timestamp 1607319584
transform 1 0 1324 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_516
timestamp 1607319584
transform -1 0 1516 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_232
timestamp 1607319584
transform 1 0 1516 0 -1 4905
box -2 -3 34 103
use FILL  FILL_48_2_0
timestamp 1607319584
transform 1 0 1548 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_2_1
timestamp 1607319584
transform 1 0 1556 0 -1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_567
timestamp 1607319584
transform 1 0 1564 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_286
timestamp 1607319584
transform 1 0 1660 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_519
timestamp 1607319584
transform -1 0 1788 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_238
timestamp 1607319584
transform -1 0 1820 0 -1 4905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_80
timestamp 1607319584
transform -1 0 1892 0 -1 4905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_19
timestamp 1607319584
transform 1 0 1892 0 -1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_561
timestamp 1607319584
transform 1 0 1964 0 -1 4905
box -2 -3 98 103
use FILL  FILL_48_3_0
timestamp 1607319584
transform 1 0 2060 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_3_1
timestamp 1607319584
transform 1 0 2068 0 -1 4905
box -2 -3 10 103
use OAI21X1  OAI21X1_274
timestamp 1607319584
transform 1 0 2076 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_273
timestamp 1607319584
transform -1 0 2140 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_566
timestamp 1607319584
transform 1 0 2140 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_283
timestamp 1607319584
transform -1 0 2268 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_284
timestamp 1607319584
transform -1 0 2300 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1025
timestamp 1607319584
transform -1 0 2396 0 -1 4905
box -2 -3 98 103
use BUFX2  BUFX2_1
timestamp 1607319584
transform 1 0 2396 0 -1 4905
box -2 -3 26 103
use OAI21X1  OAI21X1_226
timestamp 1607319584
transform 1 0 2420 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_513
timestamp 1607319584
transform 1 0 2452 0 -1 4905
box -2 -3 98 103
use BUFX4  BUFX4_14
timestamp 1607319584
transform 1 0 2548 0 -1 4905
box -2 -3 34 103
use FILL  FILL_48_4_0
timestamp 1607319584
transform 1 0 2580 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_4_1
timestamp 1607319584
transform 1 0 2588 0 -1 4905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_91
timestamp 1607319584
transform 1 0 2596 0 -1 4905
box -2 -3 74 103
use OAI21X1  OAI21X1_229
timestamp 1607319584
transform -1 0 2700 0 -1 4905
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1607319584
transform -1 0 2732 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_515
timestamp 1607319584
transform -1 0 2828 0 -1 4905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_1
timestamp 1607319584
transform -1 0 2900 0 -1 4905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_32
timestamp 1607319584
transform 1 0 2900 0 -1 4905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_310
timestamp 1607319584
transform 1 0 2972 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_1645
timestamp 1607319584
transform 1 0 3068 0 -1 4905
box -2 -3 34 103
use FILL  FILL_48_5_0
timestamp 1607319584
transform 1 0 3100 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_5_1
timestamp 1607319584
transform 1 0 3108 0 -1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_307
timestamp 1607319584
transform 1 0 3116 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_1639
timestamp 1607319584
transform 1 0 3212 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_311
timestamp 1607319584
transform 1 0 3244 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_1647
timestamp 1607319584
transform 1 0 3340 0 -1 4905
box -2 -3 34 103
use AOI21X1  AOI21X1_239
timestamp 1607319584
transform 1 0 3372 0 -1 4905
box -2 -3 34 103
use NOR2X1  NOR2X1_300
timestamp 1607319584
transform -1 0 3428 0 -1 4905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1607319584
transform -1 0 3524 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1607319584
transform 1 0 3524 0 -1 4905
box -2 -3 98 103
use FILL  FILL_48_6_0
timestamp 1607319584
transform 1 0 3620 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_6_1
timestamp 1607319584
transform 1 0 3628 0 -1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1607319584
transform 1 0 3636 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1607319584
transform 1 0 3732 0 -1 4905
box -2 -3 98 103
use NOR2X1  NOR2X1_304
timestamp 1607319584
transform 1 0 3828 0 -1 4905
box -2 -3 26 103
use AOI21X1  AOI21X1_243
timestamp 1607319584
transform -1 0 3884 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_182
timestamp 1607319584
transform 1 0 3884 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1607319584
transform -1 0 4076 0 -1 4905
box -2 -3 98 103
use INVX1  INVX1_130
timestamp 1607319584
transform 1 0 4076 0 -1 4905
box -2 -3 18 103
use FILL  FILL_48_7_0
timestamp 1607319584
transform 1 0 4092 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_7_1
timestamp 1607319584
transform 1 0 4100 0 -1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_184
timestamp 1607319584
transform 1 0 4108 0 -1 4905
box -2 -3 98 103
use NOR2X1  NOR2X1_303
timestamp 1607319584
transform -1 0 4228 0 -1 4905
box -2 -3 26 103
use AOI21X1  AOI21X1_242
timestamp 1607319584
transform -1 0 4260 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1607319584
transform 1 0 4260 0 -1 4905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_43
timestamp 1607319584
transform 1 0 4356 0 -1 4905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_42
timestamp 1607319584
transform -1 0 4500 0 -1 4905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_78
timestamp 1607319584
transform 1 0 4500 0 -1 4905
box -2 -3 74 103
use BUFX4  BUFX4_12
timestamp 1607319584
transform -1 0 4604 0 -1 4905
box -2 -3 34 103
use FILL  FILL_48_8_0
timestamp 1607319584
transform -1 0 4612 0 -1 4905
box -2 -3 10 103
use FILL  FILL_48_8_1
timestamp 1607319584
transform -1 0 4620 0 -1 4905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1607319584
transform -1 0 4716 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_166
timestamp 1607319584
transform 1 0 4716 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_471
timestamp 1607319584
transform 1 0 4812 0 -1 4905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_498
timestamp 1607319584
transform 1 0 4908 0 -1 4905
box -2 -3 98 103
use OAI21X1  OAI21X1_1313
timestamp 1607319584
transform -1 0 5036 0 -1 4905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1607319584
transform -1 0 5132 0 -1 4905
box -2 -3 98 103
use BUFX2  BUFX2_5
timestamp 1607319584
transform 1 0 5132 0 -1 4905
box -2 -3 26 103
use INVX1  INVX1_92
timestamp 1607319584
transform -1 0 5172 0 -1 4905
box -2 -3 18 103
use FILL  FILL_49_1
timestamp 1607319584
transform -1 0 5180 0 -1 4905
box -2 -3 10 103
use FILL  FILL_49_2
timestamp 1607319584
transform -1 0 5188 0 -1 4905
box -2 -3 10 103
use FILL  FILL_49_3
timestamp 1607319584
transform -1 0 5196 0 -1 4905
box -2 -3 10 103
<< labels >>
flabel metal6 s 536 -30 552 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1048 -30 1064 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s 5222 2848 5226 2852 3 FreeSans 24 0 0 0 a[0]
port 2 nsew
flabel metal2 s 3190 4928 3194 4932 3 FreeSans 24 90 0 0 a[1]
port 3 nsew
flabel metal3 s -26 3148 -22 3152 7 FreeSans 24 0 0 0 a[2]
port 4 nsew
flabel metal3 s -26 2348 -22 2352 7 FreeSans 24 0 0 0 a[3]
port 5 nsew
flabel metal3 s -26 2328 -22 2332 7 FreeSans 24 0 0 0 a[4]
port 6 nsew
flabel metal3 s -26 2508 -22 2512 7 FreeSans 24 0 0 0 a[5]
port 7 nsew
flabel metal3 s -26 2488 -22 2492 7 FreeSans 24 0 0 0 a[6]
port 8 nsew
flabel metal3 s 5222 2648 5226 2652 3 FreeSans 24 0 0 0 d[0]
port 9 nsew
flabel metal3 s -26 2948 -22 2952 7 FreeSans 24 0 0 0 d[1]
port 10 nsew
flabel metal3 s 5222 2748 5226 2752 3 FreeSans 24 0 0 0 d[2]
port 11 nsew
flabel metal3 s -26 2548 -22 2552 7 FreeSans 24 0 0 0 d[3]
port 12 nsew
flabel metal3 s 5222 2058 5226 2062 3 FreeSans 24 0 0 0 d[4]
port 13 nsew
flabel metal3 s 5222 2768 5226 2772 3 FreeSans 24 0 0 0 d[5]
port 14 nsew
flabel metal3 s 5222 1558 5226 1562 3 FreeSans 24 0 0 0 d[6]
port 15 nsew
flabel metal3 s -26 3548 -22 3552 7 FreeSans 24 0 0 0 d[7]
port 16 nsew
flabel metal2 s 3254 -22 3258 -18 7 FreeSans 24 270 0 0 we
port 17 nsew
flabel metal2 s 1294 4928 1298 4932 3 FreeSans 24 90 0 0 clk
port 18 nsew
flabel metal2 s 2406 4928 2410 4932 3 FreeSans 24 90 0 0 q[0]
port 19 nsew
flabel metal3 s -26 2468 -22 2472 7 FreeSans 24 0 0 0 q[1]
port 20 nsew
flabel metal2 s 2094 -22 2098 -18 7 FreeSans 24 270 0 0 q[2]
port 21 nsew
flabel metal3 s -26 2448 -22 2452 7 FreeSans 24 0 0 0 q[3]
port 22 nsew
flabel metal3 s 5222 4848 5226 4852 3 FreeSans 24 90 0 0 q[4]
port 23 nsew
flabel metal3 s -26 2368 -22 2372 7 FreeSans 24 0 0 0 q[5]
port 24 nsew
flabel metal3 s -26 2648 -22 2652 7 FreeSans 24 0 0 0 q[6]
port 25 nsew
flabel metal3 s -26 2148 -22 2152 7 FreeSans 24 0 0 0 q[7]
port 26 nsew
<< end >>
