* NGSPICE file created from ram_single.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

.subckt ram_single vdd gnd a[0] a[1] a[2] a[3] a[4] a[5] a[6] d[0] d[1] d[2] d[3]
+ d[4] d[5] d[6] d[7] we clk q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7]
XFILL_9_6_0 gnd vdd FILL
XNAND2X1_580 BUFX4_261/Y NOR2X1_38/A gnd NAND2X1_580/Y vdd NAND2X1
XNAND2X1_591 MUX2X1_4/S NAND2X1_591/B gnd NAND2X1_591/Y vdd NAND2X1
XFILL_17_5_0 gnd vdd FILL
XFILL_41_3_0 gnd vdd FILL
XFILL_42_8_1 gnd vdd FILL
XOAI21X1_382 NAND2X1_81/Y BUFX4_113/Y OAI21X1_382/C gnd OAI21X1_382/Y vdd OAI21X1
XOAI21X1_371 NOR2X1_22/B BUFX4_386/Y NAND2X1_588/B gnd OAI21X1_372/C vdd OAI21X1
XINVX1_402 INVX1_402/A gnd INVX1_402/Y vdd INVX1
XOAI21X1_360 BUFX4_377/Y NAND2X1_79/Y OAI21X1_360/C gnd OAI21X1_360/Y vdd OAI21X1
XINVX1_424 INVX1_424/A gnd INVX1_424/Y vdd INVX1
XOAI21X1_393 NOR2X1_32/B BUFX4_385/Y OAI21X1_393/C gnd OAI21X1_393/Y vdd OAI21X1
XINVX1_435 INVX1_435/A gnd INVX1_435/Y vdd INVX1
XINVX1_413 INVX1_413/A gnd INVX1_413/Y vdd INVX1
XINVX1_446 INVX1_446/A gnd INVX1_446/Y vdd INVX1
XINVX1_468 INVX1_468/A gnd INVX1_468/Y vdd INVX1
XINVX1_457 INVX1_457/A gnd INVX1_457/Y vdd INVX1
XINVX1_479 INVX1_479/A gnd INVX1_479/Y vdd INVX1
XFILL_32_3_0 gnd vdd FILL
XFILL_33_8_1 gnd vdd FILL
XOAI21X1_1612 NOR2X1_2/B BUFX4_348/Y NAND2X1_565/B gnd OAI21X1_1612/Y vdd OAI21X1
XOAI21X1_1623 INVX1_334/Y NOR2X1_358/Y NAND2X1_849/Y gnd DFFPOSX1_278/D vdd OAI21X1
XOAI21X1_1601 BUFX4_376/Y NAND2X1_842/Y OAI21X1_1600/Y gnd DFFPOSX1_264/D vdd OAI21X1
XOAI21X1_1645 NAND2X1_860/Y BUFX4_97/Y OAI21X1_1645/C gnd DFFPOSX1_310/D vdd OAI21X1
XOAI21X1_1656 BUFX4_412/Y BUFX4_344/Y NAND2X1_430/B gnd OAI21X1_1657/C vdd OAI21X1
XOAI21X1_1634 INVX4_3/A BUFX4_346/Y INVX1_17/A gnd OAI21X1_1634/Y vdd OAI21X1
XOAI21X1_1689 BUFX4_377/Y NAND2X1_871/Y OAI21X1_1689/C gnd DFFPOSX1_344/D vdd OAI21X1
XOAI21X1_1678 BUFX4_406/Y OAI21X1_5/B INVX1_146/A gnd OAI21X1_1679/C vdd OAI21X1
XOAI21X1_1667 INVX1_81/Y NOR2X1_378/Y NAND2X1_864/Y gnd OAI21X1_1667/Y vdd OAI21X1
XFILL_23_3_0 gnd vdd FILL
XFILL_24_8_1 gnd vdd FILL
XFILL_6_4_0 gnd vdd FILL
XMUX2X1_17 MUX2X1_17/A MUX2X1_15/Y BUFX4_60/Y gnd MUX2X1_17/Y vdd MUX2X1
XMUX2X1_28 MUX2X1_27/Y MUX2X1_28/B MUX2X1_42/S gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_39 MUX2X1_38/Y MUX2X1_39/B BUFX4_357/Y gnd MUX2X1_39/Y vdd MUX2X1
XFILL_15_8_1 gnd vdd FILL
XFILL_14_3_0 gnd vdd FILL
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XOAI21X1_190 BUFX4_113/Y NAND2X1_22/Y OAI21X1_190/C gnd OAI21X1_190/Y vdd OAI21X1
XDFFPOSX1_509 NOR2X1_37/A CLKBUF1_24/Y AOI21X1_29/Y gnd vdd DFFPOSX1
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XINVX1_243 INVX1_243/A gnd INVX1_243/Y vdd INVX1
XINVX1_232 INVX1_232/A gnd INVX1_232/Y vdd INVX1
XINVX1_254 INVX1_254/A gnd INVX1_254/Y vdd INVX1
XINVX1_276 INVX1_276/A gnd INVX1_276/Y vdd INVX1
XINVX1_265 INVX1_265/A gnd INVX1_265/Y vdd INVX1
XINVX1_298 INVX1_298/A gnd INVX1_298/Y vdd INVX1
XINVX1_287 INVX1_287/A gnd INVX1_287/Y vdd INVX1
XNAND2X1_21 INVX8_10/A INVX1_1/Y gnd NAND2X1_21/Y vdd NAND2X1
XNAND2X1_32 INVX8_3/A NOR2X1_21/Y gnd NAND2X1_32/Y vdd NAND2X1
XNAND2X1_43 BUFX4_447/Y NOR2X1_31/Y gnd NAND2X1_43/Y vdd NAND2X1
XNAND2X1_10 BUFX4_444/Y NOR2X1_1/Y gnd NAND2X1_10/Y vdd NAND2X1
XNAND2X1_54 BUFX4_448/Y NOR2X1_41/Y gnd NAND2X1_54/Y vdd NAND2X1
XNAND2X1_65 BUFX4_427/Y NOR2X1_51/Y gnd NAND2X1_65/Y vdd NAND2X1
XNAND2X1_76 BUFX4_428/Y NOR2X1_61/Y gnd NAND2X1_76/Y vdd NAND2X1
XNAND2X1_87 INVX8_5/A NOR2X1_71/Y gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_98 AOI22X1_9/D BUFX4_292/Y gnd BUFX4_294/A vdd NAND2X1
XFILL_35_1 gnd vdd FILL
XAOI21X1_214 BUFX4_376/Y NOR2X1_256/B NOR2X1_263/Y gnd DFFPOSX1_16/D vdd AOI21X1
XAOI21X1_225 AOI21X1_3/A NOR2X1_279/B NOR2X1_278/Y gnd DFFPOSX1_19/D vdd AOI21X1
XAOI21X1_203 AOI21X1_203/A AOI21X1_203/B BUFX4_364/Y gnd OAI21X1_827/A vdd AOI21X1
XAOI21X1_236 BUFX4_96/Y NOR2X1_289/B NOR2X1_291/Y gnd DFFPOSX1_62/D vdd AOI21X1
XAOI21X1_258 BUFX4_297/Y NOR2X1_325/B NOR2X1_326/Y gnd AOI21X1_258/Y vdd AOI21X1
XAOI21X1_247 BUFX4_125/Y NOR2X1_315/B NOR2X1_312/Y gnd AOI21X1_247/Y vdd AOI21X1
XAOI22X1_41 AOI22X1_41/A BUFX4_321/Y BUFX4_288/Y MUX2X1_198/Y gnd AOI22X1_41/Y vdd
+ AOI22X1
XAOI22X1_30 MUX2X1_141/Y BUFX4_354/Y BUFX4_155/Y AOI22X1_30/D gnd AOI22X1_30/Y vdd
+ AOI22X1
XAOI21X1_269 BUFX4_279/Y NOR2X1_338/B NOR2X1_339/Y gnd AOI21X1_269/Y vdd AOI21X1
XAOI22X1_74 AOI22X1_74/A AOI22X1_9/A NAND2X1_5/B AOI22X1_74/D gnd AOI22X1_74/Y vdd
+ AOI22X1
XAOI22X1_63 AOI22X1_63/A BUFX4_323/Y AOI22X1_6/C MUX2X1_306/Y gnd AOI22X1_63/Y vdd
+ AOI22X1
XAOI22X1_52 AOI22X1_52/A AOI22X1_7/B BUFX4_159/Y MUX2X1_252/Y gnd AOI22X1_52/Y vdd
+ AOI22X1
XOAI21X1_1431 BUFX4_151/Y BUFX4_390/Y NAND2X1_418/B gnd OAI21X1_1431/Y vdd OAI21X1
XOAI21X1_1420 BUFX4_99/Y NAND2X1_814/Y OAI21X1_1420/C gnd OAI21X1_1420/Y vdd OAI21X1
XOAI21X1_1464 NAND2X1_832/Y BUFX4_305/Y OAI21X1_1464/C gnd DFFPOSX1_180/D vdd OAI21X1
XOAI21X1_1475 BUFX4_417/Y BUFX4_393/Y NAND2X1_283/B gnd OAI21X1_1476/C vdd OAI21X1
XOAI21X1_1442 INVX1_70/Y NOR2X1_321/Y NAND2X1_817/Y gnd OAI21X1_1442/Y vdd OAI21X1
XOAI21X1_1453 INVX1_263/Y NOR2X1_331/Y NAND2X1_828/Y gnd OAI21X1_1453/Y vdd OAI21X1
XOAI21X1_1486 BUFX4_286/Y NAND2X1_833/Y OAI21X1_1485/Y gnd OAI21X1_1486/Y vdd OAI21X1
XOAI21X1_1497 NOR2X1_61/B BUFX4_94/Y INVX1_265/A gnd OAI21X1_1498/C vdd OAI21X1
XDFFPOSX1_1027 BUFX2_3/A CLKBUF1_64/Y NAND2X1_409/Y gnd vdd DFFPOSX1
XDFFPOSX1_1005 NOR2X1_224/A CLKBUF1_97/Y AOI21X1_182/Y gnd vdd DFFPOSX1
XDFFPOSX1_1016 INVX1_508/A CLKBUF1_59/Y OAI21X1_798/Y gnd vdd DFFPOSX1
XOAI22X1_3 OAI22X1_3/A INVX1_15/Y INVX1_16/Y OR2X2_1/Y gnd OAI22X1_3/Y vdd OAI22X1
XFILL_47_7_1 gnd vdd FILL
XFILL_46_2_0 gnd vdd FILL
XFILL_30_6_1 gnd vdd FILL
XDFFPOSX1_328 INVX1_465/A CLKBUF1_83/Y DFFPOSX1_328/D gnd vdd DFFPOSX1
XDFFPOSX1_306 INVX1_80/A CLKBUF1_12/Y OAI21X1_1637/Y gnd vdd DFFPOSX1
XDFFPOSX1_317 NAND2X1_499/B CLKBUF1_25/Y OAI21X1_1659/Y gnd vdd DFFPOSX1
XDFFPOSX1_339 INVX1_146/A CLKBUF1_99/Y DFFPOSX1_339/D gnd vdd DFFPOSX1
XNAND2X1_409 AOI22X1_24/Y AOI22X1_29/Y gnd NAND2X1_409/Y vdd NAND2X1
XFILL_37_2_0 gnd vdd FILL
XFILL_38_7_1 gnd vdd FILL
XBUFX4_382 BUFX4_385/A gnd INVX2_3/A vdd BUFX4
XBUFX4_360 a[2] gnd MUX2X1_48/S vdd BUFX4
XBUFX4_371 INVX8_15/Y gnd BUFX4_371/Y vdd BUFX4
XBUFX4_393 BUFX4_392/A gnd BUFX4_393/Y vdd BUFX4
XOAI21X1_915 INVX1_127/Y BUFX4_216/Y NAND2X1_343/Y gnd MUX2X1_92/B vdd OAI21X1
XFILL_20_1_0 gnd vdd FILL
XFILL_21_6_1 gnd vdd FILL
XOAI21X1_904 INVX1_116/Y BUFX4_194/Y OAI21X1_904/C gnd MUX2X1_83/A vdd OAI21X1
XOAI21X1_926 INVX1_138/Y BUFX4_238/Y NAND2X1_354/Y gnd MUX2X1_100/A vdd OAI21X1
XOAI21X1_937 INVX1_149/Y BUFX4_260/Y OAI21X1_937/C gnd MUX2X1_109/B vdd OAI21X1
XOAI21X1_948 INVX1_160/Y MUX2X1_5/S OAI21X1_948/C gnd MUX2X1_116/A vdd OAI21X1
XOAI21X1_959 INVX1_171/Y BUFX4_205/Y OAI21X1_959/C gnd MUX2X1_125/B vdd OAI21X1
XDFFPOSX1_840 INVX1_497/A CLKBUF1_81/Y OAI21X1_637/Y gnd vdd DFFPOSX1
XOAI21X1_1272 INVX1_484/Y BUFX4_237/Y NAND2X1_727/Y gnd MUX2X1_359/A vdd OAI21X1
XOAI21X1_1261 INVX1_473/Y BUFX4_215/Y NAND2X1_715/Y gnd MUX2X1_352/B vdd OAI21X1
XOAI21X1_1283 INVX1_495/Y BUFX4_259/Y NAND2X1_739/Y gnd MUX2X1_368/B vdd OAI21X1
XOAI21X1_1250 INVX1_462/Y BUFX4_193/Y NAND2X1_704/Y gnd MUX2X1_343/A vdd OAI21X1
XDFFPOSX1_851 INVX1_178/A CLKBUF1_49/Y OAI21X1_655/Y gnd vdd DFFPOSX1
XDFFPOSX1_884 INVX1_244/A CLKBUF1_15/Y OAI21X1_670/Y gnd vdd DFFPOSX1
XDFFPOSX1_873 MUX2X1_11/A CLKBUF1_19/Y AOI21X1_126/Y gnd vdd DFFPOSX1
XOAI21X1_1294 INVX1_506/Y MUX2X1_4/S NAND2X1_750/Y gnd MUX2X1_376/A vdd OAI21X1
XDFFPOSX1_862 NOR2X1_152/A CLKBUF1_7/Y AOI21X1_122/Y gnd vdd DFFPOSX1
XDFFPOSX1_895 NOR2X1_175/A CLKBUF1_20/Y AOI21X1_141/Y gnd vdd DFFPOSX1
XFILL_4_7_1 gnd vdd FILL
XFILL_28_2_0 gnd vdd FILL
XFILL_29_7_1 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 BUFX4_367/Y BUFX4_317/Y OAI21X1_19/C gnd OAI21X1_20/C vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_12_6_1 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XDFFPOSX1_103 INVX1_387/A CLKBUF1_89/Y OAI21X1_1375/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 INVX1_68/A CLKBUF1_32/Y DFFPOSX1_114/D gnd vdd DFFPOSX1
XDFFPOSX1_125 NAND2X1_486/B CLKBUF1_20/Y OAI21X1_1402/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 INVX1_453/A CLKBUF1_102/Y OAI21X1_1424/Y gnd vdd DFFPOSX1
XDFFPOSX1_169 NOR2X1_333/A CLKBUF1_24/Y AOI21X1_263/Y gnd vdd DFFPOSX1
XDFFPOSX1_158 NOR2X1_328/A CLKBUF1_61/Y AOI21X1_260/Y gnd vdd DFFPOSX1
XDFFPOSX1_147 INVX1_134/A CLKBUF1_98/Y DFFPOSX1_147/D gnd vdd DFFPOSX1
XNAND2X1_206 BUFX4_326/Y NOR2X1_228/Y gnd NAND2X1_206/Y vdd NAND2X1
XNAND2X1_217 BUFX4_205/Y NAND2X1_217/B gnd OAI21X1_805/C vdd NAND2X1
XNAND2X1_239 BUFX4_233/Y DFFPOSX1_73/Q gnd OAI21X1_823/C vdd NAND2X1
XNAND2X1_228 BUFX4_221/Y NOR2X1_13/A gnd OAI21X1_816/C vdd NAND2X1
XBUFX4_190 BUFX4_24/Y gnd BUFX4_190/Y vdd BUFX4
XNOR2X1_261 NOR2X1_261/A NOR2X1_256/B gnd NOR2X1_261/Y vdd NOR2X1
XNOR2X1_250 MUX2X1_84/S INVX4_1/Y gnd AOI22X1_1/B vdd NOR2X1
XNOR2X1_272 NOR2X1_272/A NOR2X1_265/Y gnd NOR2X1_272/Y vdd NOR2X1
XNOR2X1_294 INVX4_2/Y NOR2X1_294/B gnd INVX8_10/A vdd NOR2X1
XNOR2X1_283 NOR2X1_283/A NOR2X1_279/B gnd NOR2X1_283/Y vdd NOR2X1
XOAI21X1_701 BUFX4_146/Y BUFX4_67/Y NAND2X1_607/B gnd OAI21X1_702/C vdd OAI21X1
XOAI21X1_712 INVX1_438/Y NOR2X1_177/Y NAND2X1_181/Y gnd OAI21X1_712/Y vdd OAI21X1
XOAI21X1_723 INVX1_248/Y NOR2X1_199/Y OAI21X1_723/C gnd OAI21X1_723/Y vdd OAI21X1
XOAI21X1_767 BUFX4_302/Y OAI21X1_761/B OAI21X1_767/C gnd OAI21X1_767/Y vdd OAI21X1
XOAI21X1_734 BUFX4_455/Y BUFX4_440/Y INVX1_249/A gnd OAI21X1_735/C vdd OAI21X1
XOAI21X1_745 BUFX4_130/Y OAI21X1_757/B OAI21X1_745/C gnd OAI21X1_745/Y vdd OAI21X1
XOAI21X1_756 NOR2X1_72/B INVX2_5/A NAND2X1_680/B gnd OAI21X1_757/C vdd OAI21X1
XOAI21X1_778 BUFX4_308/Y BUFX4_438/Y INVX1_123/A gnd OAI21X1_779/C vdd OAI21X1
XOAI21X1_789 BUFX4_281/Y NAND2X1_201/Y OAI21X1_789/C gnd OAI21X1_789/Y vdd OAI21X1
XMUX2X1_201 MUX2X1_201/A MUX2X1_201/B MUX2X1_69/S gnd AOI22X1_42/A vdd MUX2X1
XMUX2X1_223 MUX2X1_223/A MUX2X1_223/B BUFX4_80/Y gnd MUX2X1_225/B vdd MUX2X1
XMUX2X1_212 MUX2X1_212/A MUX2X1_212/B BUFX4_49/Y gnd MUX2X1_213/A vdd MUX2X1
XMUX2X1_245 MUX2X1_245/A MUX2X1_245/B BUFX4_80/Y gnd MUX2X1_245/Y vdd MUX2X1
XOAI21X1_1080 INVX1_292/Y BUFX4_249/Y NAND2X1_520/Y gnd MUX2X1_215/A vdd OAI21X1
XMUX2X1_256 MUX2X1_256/A MUX2X1_256/B BUFX4_63/Y gnd MUX2X1_256/Y vdd MUX2X1
XMUX2X1_234 MUX2X1_233/Y MUX2X1_232/Y MUX2X1_69/S gnd MUX2X1_234/Y vdd MUX2X1
XOAI21X1_1091 INVX1_303/Y BUFX4_271/Y NAND2X1_532/Y gnd MUX2X1_224/B vdd OAI21X1
XDFFPOSX1_692 INVX1_232/A CLKBUF1_47/Y OAI21X1_488/Y gnd vdd DFFPOSX1
XDFFPOSX1_670 NAND2X1_591/B CLKBUF1_38/Y OAI21X1_444/Y gnd vdd DFFPOSX1
XDFFPOSX1_681 NAND2X1_265/B CLKBUF1_96/Y OAI21X1_466/Y gnd vdd DFFPOSX1
XMUX2X1_278 MUX2X1_278/A MUX2X1_278/B BUFX4_60/Y gnd MUX2X1_279/A vdd MUX2X1
XMUX2X1_267 MUX2X1_266/Y MUX2X1_267/B MUX2X1_69/S gnd MUX2X1_267/Y vdd MUX2X1
XMUX2X1_289 MUX2X1_289/A MUX2X1_289/B INVX4_1/A gnd MUX2X1_291/B vdd MUX2X1
XNAND2X1_773 BUFX4_430/Y NOR2X1_264/Y gnd NAND2X1_773/Y vdd NAND2X1
XNAND2X1_751 MUX2X1_5/S NOR2X1_227/A gnd NAND2X1_751/Y vdd NAND2X1
XNAND2X1_762 BUFX4_137/Y NOR2X1_254/Y gnd NAND2X1_762/Y vdd NAND2X1
XNAND2X1_740 BUFX4_260/Y NOR2X1_143/A gnd NAND2X1_740/Y vdd NAND2X1
XNAND2X1_784 BUFX4_449/Y NOR2X1_284/Y gnd NAND2X1_784/Y vdd NAND2X1
XNAND2X1_795 BUFX4_450/Y NOR2X1_297/Y gnd NAND2X1_795/Y vdd NAND2X1
XFILL_44_5_1 gnd vdd FILL
XFILL_43_0_0 gnd vdd FILL
XBUFX4_30 a[0] gnd BUFX4_30/Y vdd BUFX4
XBUFX4_52 BUFX4_52/A gnd BUFX4_52/Y vdd BUFX4
XBUFX4_41 BUFX4_41/A gnd BUFX4_41/Y vdd BUFX4
XBUFX4_85 BUFX4_84/A gnd BUFX4_85/Y vdd BUFX4
XBUFX4_96 INVX8_7/Y gnd BUFX4_96/Y vdd BUFX4
XBUFX4_63 BUFX4_62/A gnd BUFX4_63/Y vdd BUFX4
XBUFX4_74 a[1] gnd BUFX4_3/A vdd BUFX4
XFILL_34_0_0 gnd vdd FILL
XFILL_35_5_1 gnd vdd FILL
XFILL_1_5_1 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_26_5_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XINVX8_11 INVX8_11/A gnd INVX8_11/Y vdd INVX8
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOAI21X1_531 BUFX4_150/Y NOR2X1_91/A NAND2X1_318/B gnd OAI21X1_532/C vdd OAI21X1
XOAI21X1_520 BUFX4_299/Y NAND2X1_99/Y OAI21X1_520/C gnd OAI21X1_520/Y vdd OAI21X1
XOAI21X1_564 INVX1_236/Y NOR2X1_101/Y NAND2X1_120/Y gnd OAI21X1_564/Y vdd OAI21X1
XOAI21X1_575 NOR2X1_1/B BUFX4_107/Y INVX1_237/A gnd OAI21X1_576/C vdd OAI21X1
XOAI21X1_542 BUFX4_281/Y OAI21X1_544/B OAI21X1_542/C gnd OAI21X1_542/Y vdd OAI21X1
XOAI21X1_553 INVX1_59/Y NOR2X1_91/Y OAI21X1_553/C gnd OAI21X1_553/Y vdd OAI21X1
XOAI21X1_586 BUFX4_130/Y OAI21X1_590/B OAI21X1_586/C gnd OAI21X1_586/Y vdd OAI21X1
XOAI21X1_597 BUFX4_148/Y INVX1_3/A OAI21X1_597/C gnd OAI21X1_598/C vdd OAI21X1
XFILL_9_6_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XNAND2X1_570 BUFX4_241/Y NAND2X1_570/B gnd NAND2X1_570/Y vdd NAND2X1
XNAND2X1_581 AOI22X1_52/Y AOI22X1_53/Y gnd AOI22X1_54/D vdd NAND2X1
XNAND2X1_592 MUX2X1_8/S NAND2X1_592/B gnd NAND2X1_592/Y vdd NAND2X1
XFILL_16_0_0 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_41_3_1 gnd vdd FILL
XOAI21X1_350 BUFX4_109/Y NAND2X1_79/Y OAI21X1_350/C gnd OAI21X1_350/Y vdd OAI21X1
XOAI21X1_361 NOR2X1_22/B NOR2X1_61/A NAND2X1_261/B gnd OAI21X1_362/C vdd OAI21X1
XOAI21X1_383 BUFX4_171/Y NOR2X1_61/A INVX1_228/A gnd OAI21X1_383/Y vdd OAI21X1
XOAI21X1_372 BUFX4_102/Y NAND2X1_80/Y OAI21X1_372/C gnd OAI21X1_372/Y vdd OAI21X1
XINVX1_403 INVX1_403/A gnd INVX1_403/Y vdd INVX1
XOAI21X1_394 BUFX4_127/Y NAND2X1_82/Y OAI21X1_393/Y gnd OAI21X1_394/Y vdd OAI21X1
XINVX1_425 INVX1_425/A gnd INVX1_425/Y vdd INVX1
XINVX1_414 INVX1_414/A gnd INVX1_414/Y vdd INVX1
XINVX1_458 INVX1_458/A gnd INVX1_458/Y vdd INVX1
XINVX1_447 INVX1_447/A gnd INVX1_447/Y vdd INVX1
XINVX1_469 INVX1_469/A gnd INVX1_469/Y vdd INVX1
XINVX1_436 INVX1_436/A gnd INVX1_436/Y vdd INVX1
XFILL_32_3_1 gnd vdd FILL
XOAI21X1_1613 BUFX4_97/Y NAND2X1_843/Y OAI21X1_1612/Y gnd OAI21X1_1613/Y vdd OAI21X1
XOAI21X1_1624 INVX1_398/Y NOR2X1_358/Y NAND2X1_850/Y gnd OAI21X1_1624/Y vdd OAI21X1
XOAI21X1_1602 BUFX4_151/Y BUFX4_345/Y NAND2X1_217/B gnd OAI21X1_1602/Y vdd OAI21X1
XOAI21X1_1646 BUFX4_168/Y BUFX4_343/Y INVX1_400/A gnd OAI21X1_1647/C vdd OAI21X1
XOAI21X1_1657 BUFX4_305/Y NAND2X1_861/Y OAI21X1_1657/C gnd OAI21X1_1657/Y vdd OAI21X1
XOAI21X1_1635 NAND2X1_860/Y BUFX4_129/Y OAI21X1_1634/Y gnd DFFPOSX1_305/D vdd OAI21X1
XOAI21X1_1679 BUFX4_109/Y NAND2X1_871/Y OAI21X1_1679/C gnd DFFPOSX1_339/D vdd OAI21X1
XOAI21X1_1668 INVX1_145/Y NOR2X1_378/Y NAND2X1_865/Y gnd OAI21X1_1668/Y vdd OAI21X1
XFILL_23_3_1 gnd vdd FILL
XFILL_6_4_1 gnd vdd FILL
XMUX2X1_18 MUX2X1_18/A MUX2X1_18/B BUFX4_190/Y gnd MUX2X1_20/B vdd MUX2X1
XMUX2X1_29 MUX2X1_29/A MUX2X1_29/B BUFX4_199/Y gnd MUX2X1_29/Y vdd MUX2X1
XFILL_14_3_1 gnd vdd FILL
XAOI22X1_1 AOI22X1_1/A AOI22X1_1/B AOI22X1_1/C AOI22X1_1/D gnd NAND3X1_1/C vdd AOI22X1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XOAI21X1_191 BUFX4_147/Y BUFX4_133/Y OAI21X1_191/C gnd OAI21X1_191/Y vdd OAI21X1
XOAI21X1_180 BUFX4_98/Y NAND2X1_21/Y OAI21X1_180/C gnd OAI21X1_180/Y vdd OAI21X1
XINVX1_244 INVX1_244/A gnd INVX1_244/Y vdd INVX1
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XINVX1_233 INVX1_233/A gnd INVX1_233/Y vdd INVX1
XINVX1_222 INVX1_222/A gnd INVX1_222/Y vdd INVX1
XINVX1_266 INVX1_266/A gnd INVX1_266/Y vdd INVX1
XINVX1_255 INVX1_255/A gnd INVX1_255/Y vdd INVX1
XINVX1_277 INVX1_277/A gnd INVX1_277/Y vdd INVX1
XINVX1_299 INVX1_299/A gnd INVX1_299/Y vdd INVX1
XINVX1_288 INVX1_288/A gnd INVX1_288/Y vdd INVX1
XNAND2X1_22 INVX8_11/A INVX1_1/Y gnd NAND2X1_22/Y vdd NAND2X1
XNAND2X1_33 INVX8_4/A NOR2X1_21/Y gnd NAND2X1_33/Y vdd NAND2X1
XNAND2X1_11 BUFX4_326/Y NOR2X1_1/Y gnd NAND2X1_11/Y vdd NAND2X1
XNAND2X1_77 INVX2_3/Y INVX8_12/A gnd NAND2X1_77/Y vdd NAND2X1
XNAND2X1_44 BUFX4_329/Y NOR2X1_31/Y gnd NAND2X1_44/Y vdd NAND2X1
XNAND2X1_55 BUFX4_330/Y NOR2X1_41/Y gnd NAND2X1_55/Y vdd NAND2X1
XNAND2X1_66 INVX2_2/Y INVX4_3/Y gnd NAND2X1_66/Y vdd NAND2X1
XNAND2X1_88 INVX8_6/A NOR2X1_71/Y gnd NAND2X1_88/Y vdd NAND2X1
XNAND2X1_99 INVX8_10/A INVX1_2/Y gnd NAND2X1_99/Y vdd NAND2X1
XAOI21X1_215 BUFX4_131/Y NOR2X1_265/Y NOR2X1_266/Y gnd DFFPOSX1_41/D vdd AOI21X1
XAOI21X1_204 AOI21X1_204/A AOI21X1_204/B INVX2_6/Y gnd OAI21X1_827/B vdd AOI21X1
XAOI21X1_237 BUFX4_282/Y NOR2X1_289/B NOR2X1_292/Y gnd DFFPOSX1_63/D vdd AOI21X1
XAOI21X1_226 BUFX4_304/Y NOR2X1_279/B NOR2X1_279/Y gnd AOI21X1_226/Y vdd AOI21X1
XAOI21X1_248 BUFX4_422/Y NOR2X1_315/B NOR2X1_313/Y gnd AOI21X1_248/Y vdd AOI21X1
XAOI22X1_42 AOI22X1_42/A BUFX4_349/Y BUFX4_156/Y MUX2X1_204/Y gnd AOI22X1_42/Y vdd
+ AOI22X1
XAOI22X1_31 AOI22X1_31/A BUFX4_323/Y BUFX4_288/Y MUX2X1_150/Y gnd AOI22X1_31/Y vdd
+ AOI22X1
XAOI22X1_20 MUX2X1_93/Y BUFX4_354/Y BUFX4_155/Y MUX2X1_96/Y gnd AOI22X1_20/Y vdd AOI22X1
XAOI21X1_259 BUFX4_397/Y NOR2X1_325/B NOR2X1_327/Y gnd AOI21X1_259/Y vdd AOI21X1
XAOI22X1_75 AOI22X1_75/A BUFX4_352/Y BUFX4_157/Y MUX2X1_360/Y gnd AOI22X1_75/Y vdd
+ AOI22X1
XAOI22X1_53 AOI22X1_53/A BUFX4_320/Y INVX1_11/A AOI22X1_53/D gnd AOI22X1_53/Y vdd
+ AOI22X1
XAOI22X1_64 AOI22X1_64/A AOI22X1_9/A NAND2X1_5/B AOI22X1_64/D gnd AOI22X1_64/Y vdd
+ AOI22X1
XOAI21X1_1432 BUFX4_304/Y NAND2X1_815/Y OAI21X1_1431/Y gnd OAI21X1_1432/Y vdd OAI21X1
XOAI21X1_1421 BUFX4_460/Y BUFX4_388/Y INVX1_389/A gnd OAI21X1_1422/C vdd OAI21X1
XOAI21X1_1410 BUFX4_125/Y NAND2X1_814/Y OAI21X1_1409/Y gnd OAI21X1_1410/Y vdd OAI21X1
XOAI21X1_1465 BUFX4_167/Y INVX2_8/A INVX1_264/A gnd OAI21X1_1465/Y vdd OAI21X1
XOAI21X1_1443 INVX1_134/Y NOR2X1_321/Y NAND2X1_818/Y gnd DFFPOSX1_147/D vdd OAI21X1
XOAI21X1_1454 INVX1_327/Y NOR2X1_331/Y NAND2X1_829/Y gnd OAI21X1_1454/Y vdd OAI21X1
XOAI21X1_1487 BUFX4_417/Y BUFX4_392/Y NAND2X1_697/B gnd OAI21X1_1487/Y vdd OAI21X1
XOAI21X1_1476 BUFX4_420/Y NAND2X1_833/Y OAI21X1_1476/C gnd OAI21X1_1476/Y vdd OAI21X1
XOAI21X1_1498 BUFX4_402/Y NAND2X1_834/Y OAI21X1_1498/C gnd OAI21X1_1498/Y vdd OAI21X1
XDFFPOSX1_1017 MUX2X1_26/A CLKBUF1_66/Y AOI21X1_187/Y gnd vdd DFFPOSX1
XDFFPOSX1_1006 NOR2X1_225/A CLKBUF1_79/Y AOI21X1_183/Y gnd vdd DFFPOSX1
XDFFPOSX1_1028 BUFX2_4/A CLKBUF1_65/Y NAND2X1_478/Y gnd vdd DFFPOSX1
XFILL_46_2_1 gnd vdd FILL
XDFFPOSX1_307 INVX1_144/A CLKBUF1_32/Y DFFPOSX1_307/D gnd vdd DFFPOSX1
XDFFPOSX1_329 NOR2X1_380/A CLKBUF1_6/Y AOI21X1_302/Y gnd vdd DFFPOSX1
XDFFPOSX1_318 NAND2X1_568/B CLKBUF1_53/Y DFFPOSX1_318/D gnd vdd DFFPOSX1
XFILL_37_2_1 gnd vdd FILL
XBUFX4_350 BUFX4_354/A gnd BUFX4_350/Y vdd BUFX4
XBUFX4_361 a[2] gnd MUX2X1_84/S vdd BUFX4
XBUFX4_372 INVX8_9/Y gnd BUFX4_372/Y vdd BUFX4
XBUFX4_383 BUFX4_385/A gnd NOR2X1_61/A vdd BUFX4
XBUFX4_394 INVX8_6/Y gnd BUFX4_394/Y vdd BUFX4
XOAI21X1_905 INVX1_117/Y BUFX4_196/Y NAND2X1_331/Y gnd MUX2X1_85/B vdd OAI21X1
XOAI21X1_916 INVX1_128/Y BUFX4_218/Y OAI21X1_916/C gnd MUX2X1_92/A vdd OAI21X1
XOAI21X1_949 INVX1_161/Y MUX2X1_9/S NAND2X1_379/Y gnd MUX2X1_118/B vdd OAI21X1
XOAI21X1_927 INVX1_139/Y BUFX4_240/Y NAND2X1_355/Y gnd MUX2X1_101/B vdd OAI21X1
XFILL_20_1_1 gnd vdd FILL
XOAI21X1_938 INVX1_150/Y BUFX4_262/Y NAND2X1_367/Y gnd MUX2X1_109/A vdd OAI21X1
XOAI21X1_1240 INVX1_452/Y BUFX4_272/Y NAND2X1_693/Y gnd MUX2X1_335/A vdd OAI21X1
XDFFPOSX1_841 MUX2X1_8/A CLKBUF1_7/Y OAI21X1_639/Y gnd vdd DFFPOSX1
XOAI21X1_1273 INVX1_485/Y BUFX4_239/Y NAND2X1_728/Y gnd MUX2X1_361/B vdd OAI21X1
XDFFPOSX1_830 NOR2X1_141/A CLKBUF1_40/Y AOI21X1_113/Y gnd vdd DFFPOSX1
XOAI21X1_1262 INVX1_474/Y BUFX4_217/Y NAND2X1_716/Y gnd MUX2X1_352/A vdd OAI21X1
XOAI21X1_1251 INVX1_463/Y BUFX4_195/Y NAND2X1_705/Y gnd MUX2X1_344/B vdd OAI21X1
XDFFPOSX1_863 NOR2X1_153/A CLKBUF1_95/Y AOI21X1_123/Y gnd vdd DFFPOSX1
XOAI21X1_1295 INVX1_507/Y MUX2X1_8/S NAND2X1_751/Y gnd MUX2X1_377/B vdd OAI21X1
XOAI21X1_1284 INVX1_496/Y BUFX4_261/Y NAND2X1_740/Y gnd MUX2X1_368/A vdd OAI21X1
XDFFPOSX1_852 INVX1_242/A CLKBUF1_54/Y OAI21X1_656/Y gnd vdd DFFPOSX1
XDFFPOSX1_874 NOR2X1_159/A CLKBUF1_13/Y AOI21X1_127/Y gnd vdd DFFPOSX1
XDFFPOSX1_896 NOR2X1_176/A CLKBUF1_81/Y AOI21X1_142/Y gnd vdd DFFPOSX1
XDFFPOSX1_885 INVX1_308/A CLKBUF1_53/Y OAI21X1_671/Y gnd vdd DFFPOSX1
XFILL_3_2_1 gnd vdd FILL
XFILL_28_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XDFFPOSX1_115 INVX1_132/A CLKBUF1_17/Y OAI21X1_1382/Y gnd vdd DFFPOSX1
XDFFPOSX1_137 NAND2X1_247/B CLKBUF1_98/Y OAI21X1_1426/Y gnd vdd DFFPOSX1
XDFFPOSX1_104 INVX1_451/A CLKBUF1_25/Y OAI21X1_1376/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 NAND2X1_555/B CLKBUF1_55/Y OAI21X1_1404/Y gnd vdd DFFPOSX1
XDFFPOSX1_148 INVX1_198/A CLKBUF1_61/Y OAI21X1_1444/Y gnd vdd DFFPOSX1
XDFFPOSX1_159 NOR2X1_329/A CLKBUF1_98/Y AOI21X1_261/Y gnd vdd DFFPOSX1
XNAND2X1_207 BUFX4_136/Y NOR2X1_228/Y gnd OAI21X1_797/C vdd NAND2X1
XNAND2X1_218 BUFX4_207/Y OAI21X1_17/C gnd NAND2X1_218/Y vdd NAND2X1
XNAND2X1_229 BUFX4_223/Y NAND2X1_229/B gnd NAND2X1_229/Y vdd NAND2X1
XBUFX4_191 BUFX4_28/Y gnd BUFX4_191/Y vdd BUFX4
XBUFX4_180 BUFX4_27/Y gnd MUX2X1_1/S vdd BUFX4
XNOR2X1_251 BUFX4_362/Y BUFX4_80/Y gnd AOI22X1_1/C vdd NOR2X1
XNOR2X1_240 a[4] INVX1_7/Y gnd BUFX4_155/A vdd NOR2X1
XNOR2X1_273 NOR2X1_273/A NOR2X1_265/Y gnd NOR2X1_273/Y vdd NOR2X1
XNOR2X1_262 NOR2X1_262/A NOR2X1_256/B gnd NOR2X1_262/Y vdd NOR2X1
XNOR2X1_284 NAND3X1_7/Y INVX1_509/Y gnd NOR2X1_284/Y vdd NOR2X1
XNOR2X1_295 INVX4_2/Y NOR2X1_255/A gnd INVX8_11/A vdd NOR2X1
XOAI21X1_713 INVX1_502/Y NOR2X1_177/Y OAI21X1_713/C gnd OAI21X1_713/Y vdd OAI21X1
XOAI21X1_702 BUFX4_98/Y OAI21X1_704/B OAI21X1_702/C gnd OAI21X1_702/Y vdd OAI21X1
XOAI21X1_724 INVX1_312/Y NOR2X1_199/Y NAND2X1_193/Y gnd OAI21X1_724/Y vdd OAI21X1
XOAI21X1_746 NOR2X1_72/B BUFX4_441/Y NAND2X1_335/B gnd OAI21X1_747/C vdd OAI21X1
XOAI21X1_735 BUFX4_302/Y OAI21X1_729/B OAI21X1_735/C gnd OAI21X1_735/Y vdd OAI21X1
XOAI21X1_757 BUFX4_281/Y OAI21X1_757/B OAI21X1_757/C gnd OAI21X1_757/Y vdd OAI21X1
XOAI21X1_779 BUFX4_419/Y NAND2X1_201/Y OAI21X1_779/C gnd OAI21X1_779/Y vdd OAI21X1
XOAI21X1_768 BUFX4_409/Y BUFX4_442/Y INVX1_314/A gnd OAI21X1_769/C vdd OAI21X1
XMUX2X1_202 MUX2X1_202/A MUX2X1_202/B BUFX4_81/Y gnd MUX2X1_202/Y vdd MUX2X1
XMUX2X1_213 MUX2X1_213/A MUX2X1_213/B MUX2X1_48/S gnd AOI22X1_45/A vdd MUX2X1
XMUX2X1_246 MUX2X1_245/Y MUX2X1_244/Y MUX2X1_48/S gnd MUX2X1_246/Y vdd MUX2X1
XMUX2X1_235 MUX2X1_235/A MUX2X1_235/B BUFX4_50/Y gnd MUX2X1_235/Y vdd MUX2X1
XOAI21X1_1070 INVX1_282/Y BUFX4_229/Y NAND2X1_509/Y gnd MUX2X1_208/A vdd OAI21X1
XMUX2X1_224 MUX2X1_224/A MUX2X1_224/B BUFX4_81/Y gnd MUX2X1_224/Y vdd MUX2X1
XOAI21X1_1081 INVX1_293/Y BUFX4_251/Y NAND2X1_521/Y gnd MUX2X1_217/B vdd OAI21X1
XDFFPOSX1_693 INVX1_296/A CLKBUF1_47/Y OAI21X1_490/Y gnd vdd DFFPOSX1
XDFFPOSX1_660 INVX1_230/A CLKBUF1_96/Y OAI21X1_424/Y gnd vdd DFFPOSX1
XOAI21X1_1092 INVX1_304/Y BUFX4_273/Y NAND2X1_533/Y gnd MUX2X1_224/A vdd OAI21X1
XDFFPOSX1_682 NAND2X1_316/B CLKBUF1_99/Y OAI21X1_468/Y gnd vdd DFFPOSX1
XMUX2X1_279 MUX2X1_279/A MUX2X1_279/B MUX2X1_48/S gnd MUX2X1_279/Y vdd MUX2X1
XDFFPOSX1_671 OAI21X1_445/C CLKBUF1_58/Y OAI21X1_446/Y gnd vdd DFFPOSX1
XMUX2X1_257 MUX2X1_257/A MUX2X1_257/B BUFX4_51/Y gnd MUX2X1_258/A vdd MUX2X1
XMUX2X1_268 MUX2X1_268/A MUX2X1_268/B BUFX4_80/Y gnd MUX2X1_270/B vdd MUX2X1
XNAND2X1_730 BUFX4_242/Y NAND2X1_730/B gnd NAND2X1_730/Y vdd NAND2X1
XNAND2X1_752 MUX2X1_9/S NOR2X1_238/A gnd NAND2X1_752/Y vdd NAND2X1
XNAND2X1_763 BUFX4_428/Y NOR2X1_254/Y gnd NAND2X1_763/Y vdd NAND2X1
XNAND2X1_741 BUFX4_262/Y NAND2X1_741/B gnd NAND2X1_741/Y vdd NAND2X1
XNAND2X1_796 BUFX4_332/Y NOR2X1_297/Y gnd NAND2X1_796/Y vdd NAND2X1
XNAND2X1_774 BUFX4_188/Y AOI22X1_1/B gnd NOR2X1_265/B vdd NAND2X1
XNAND2X1_785 NAND2X1_8/A NOR2X1_284/Y gnd NAND2X1_785/Y vdd NAND2X1
XFILL_43_0_1 gnd vdd FILL
XBUFX4_20 BUFX4_70/Y gnd BUFX4_20/Y vdd BUFX4
XBUFX4_31 a[0] gnd BUFX4_31/Y vdd BUFX4
XBUFX4_42 BUFX4_41/A gnd BUFX4_42/Y vdd BUFX4
XBUFX4_53 BUFX4_52/A gnd BUFX4_53/Y vdd BUFX4
XBUFX4_64 BUFX4_64/A gnd BUFX4_64/Y vdd BUFX4
XBUFX4_75 a[1] gnd BUFX4_75/Y vdd BUFX4
XBUFX4_86 BUFX4_84/A gnd BUFX4_86/Y vdd BUFX4
XBUFX4_97 INVX8_7/Y gnd BUFX4_97/Y vdd BUFX4
XFILL_34_0_1 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XFILL_25_0_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XINVX8_12 INVX8_12/A gnd INVX8_12/Y vdd INVX8
XINVX1_7 a[3] gnd INVX1_7/Y vdd INVX1
XOAI21X1_510 BUFX4_284/Y NAND2X1_97/Y OAI21X1_510/C gnd OAI21X1_510/Y vdd OAI21X1
XOAI21X1_532 BUFX4_418/Y OAI21X1_544/B OAI21X1_532/C gnd OAI21X1_532/Y vdd OAI21X1
XOAI21X1_521 BUFX4_461/Y INVX1_2/A INVX1_297/A gnd OAI21X1_522/C vdd OAI21X1
XOAI21X1_565 INVX1_300/Y NOR2X1_101/Y OAI21X1_565/C gnd OAI21X1_565/Y vdd OAI21X1
XOAI21X1_554 INVX1_107/Y NOR2X1_91/Y OAI21X1_554/C gnd OAI21X1_554/Y vdd OAI21X1
XOAI21X1_543 BUFX4_153/Y BUFX4_293/Y OAI21X1_543/C gnd OAI21X1_543/Y vdd OAI21X1
XOAI21X1_587 BUFX4_148/Y BUFX4_107/Y OAI21X1_587/C gnd OAI21X1_588/C vdd OAI21X1
XOAI21X1_598 BUFX4_281/Y OAI21X1_590/B OAI21X1_598/C gnd OAI21X1_598/Y vdd OAI21X1
XOAI21X1_576 BUFX4_298/Y OAI21X1_584/B OAI21X1_576/C gnd OAI21X1_576/Y vdd OAI21X1
XDFFPOSX1_490 NOR2X1_24/A CLKBUF1_37/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XFILL_8_1_1 gnd vdd FILL
XNAND2X1_571 BUFX4_243/Y OAI21X1_27/C gnd NAND2X1_571/Y vdd NAND2X1
XNAND2X1_560 BUFX4_223/Y NAND2X1_560/B gnd NAND2X1_560/Y vdd NAND2X1
XNAND2X1_593 MUX2X1_11/S NAND2X1_593/B gnd NAND2X1_593/Y vdd NAND2X1
XNAND2X1_582 BUFX4_263/Y OAI21X1_251/C gnd NAND2X1_582/Y vdd NAND2X1
XFILL_45_8_0 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XFILL_36_8_0 gnd vdd FILL
XFILL_2_8_0 gnd vdd FILL
XFILL_27_8_0 gnd vdd FILL
XFILL_10_7_0 gnd vdd FILL
XOAI21X1_340 BUFX4_102/Y NAND2X1_78/Y OAI21X1_339/Y gnd OAI21X1_340/Y vdd OAI21X1
XOAI21X1_362 BUFX4_123/Y NAND2X1_80/Y OAI21X1_362/C gnd OAI21X1_362/Y vdd OAI21X1
XOAI21X1_373 BUFX4_370/Y BUFX4_384/Y NAND2X1_657/B gnd OAI21X1_373/Y vdd OAI21X1
XOAI21X1_351 BUFX4_307/Y BUFX4_387/Y INVX1_227/A gnd OAI21X1_351/Y vdd OAI21X1
XOAI21X1_384 NAND2X1_81/Y BUFX4_303/Y OAI21X1_383/Y gnd OAI21X1_384/Y vdd OAI21X1
XOAI21X1_395 BUFX4_415/Y BUFX4_386/Y NAND2X1_313/B gnd OAI21X1_396/C vdd OAI21X1
XINVX1_404 INVX1_404/A gnd INVX1_404/Y vdd INVX1
XINVX1_426 INVX1_426/A gnd INVX1_426/Y vdd INVX1
XINVX1_415 INVX1_415/A gnd INVX1_415/Y vdd INVX1
XINVX1_437 INVX1_437/A gnd INVX1_437/Y vdd INVX1
XINVX1_459 INVX1_459/A gnd INVX1_459/Y vdd INVX1
XINVX1_448 INVX1_448/A gnd INVX1_448/Y vdd INVX1
XNAND2X1_390 BUFX4_206/Y NOR2X1_105/A gnd OAI21X1_960/C vdd NAND2X1
XFILL_18_8_0 gnd vdd FILL
XOAI21X1_1614 NOR2X1_2/B BUFX4_345/Y NAND2X1_634/B gnd OAI21X1_1614/Y vdd OAI21X1
XOAI21X1_1603 BUFX4_125/Y NAND2X1_843/Y OAI21X1_1602/Y gnd OAI21X1_1603/Y vdd OAI21X1
XOAI21X1_1647 NAND2X1_860/Y BUFX4_286/Y OAI21X1_1647/C gnd DFFPOSX1_311/D vdd OAI21X1
XOAI21X1_1636 BUFX4_166/Y BUFX4_345/Y INVX1_80/A gnd OAI21X1_1637/C vdd OAI21X1
XOAI21X1_1625 INVX1_462/Y NOR2X1_358/Y NAND2X1_851/Y gnd DFFPOSX1_280/D vdd OAI21X1
XOAI21X1_1669 INVX1_209/Y NOR2X1_378/Y NAND2X1_866/Y gnd DFFPOSX1_324/D vdd OAI21X1
XOAI21X1_1658 BUFX4_416/Y INVX2_10/A NAND2X1_499/B gnd OAI21X1_1658/Y vdd OAI21X1
XMUX2X1_19 MUX2X1_19/A MUX2X1_19/B BUFX4_191/Y gnd MUX2X1_19/Y vdd MUX2X1
XFILL_42_6_0 gnd vdd FILL
XAOI22X1_2 AOI22X1_2/A AOI22X1_1/B AOI22X1_1/C AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XOAI21X1_192 BUFX4_301/Y NAND2X1_22/Y OAI21X1_191/Y gnd OAI21X1_192/Y vdd OAI21X1
XOAI21X1_181 NOR2X1_61/B BUFX4_133/Y INVX1_409/A gnd OAI21X1_181/Y vdd OAI21X1
XOAI21X1_170 AOI21X1_1/A NAND2X1_21/Y OAI21X1_169/Y gnd OAI21X1_170/Y vdd OAI21X1
XINVX1_223 INVX1_223/A gnd INVX1_223/Y vdd INVX1
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XINVX1_234 INVX1_234/A gnd INVX1_234/Y vdd INVX1
XINVX1_267 INVX1_267/A gnd INVX1_267/Y vdd INVX1
XINVX1_245 INVX1_245/A gnd INVX1_245/Y vdd INVX1
XINVX1_256 INVX1_256/A gnd INVX1_256/Y vdd INVX1
XINVX1_289 INVX1_289/A gnd INVX1_289/Y vdd INVX1
XINVX1_278 INVX1_278/A gnd INVX1_278/Y vdd INVX1
XNAND2X1_23 BUFX4_162/Y NOR2X1_11/Y gnd NAND2X1_23/Y vdd NAND2X1
XNAND2X1_34 INVX8_5/A NOR2X1_21/Y gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_12 BUFX4_136/Y NOR2X1_1/Y gnd OAI21X1_71/C vdd NAND2X1
XNAND2X1_45 BUFX4_139/Y NOR2X1_31/Y gnd NAND2X1_45/Y vdd NAND2X1
XNAND2X1_56 BUFX4_140/Y NOR2X1_41/Y gnd NAND2X1_56/Y vdd NAND2X1
XNAND2X1_67 INVX8_16/A INVX2_2/Y gnd NAND2X1_67/Y vdd NAND2X1
XNAND2X1_78 INVX2_3/Y INVX8_13/A gnd NAND2X1_78/Y vdd NAND2X1
XNAND2X1_89 INVX8_7/A NOR2X1_71/Y gnd NAND2X1_89/Y vdd NAND2X1
XFILL_33_6_0 gnd vdd FILL
XAOI21X1_216 BUFX4_426/Y NOR2X1_265/Y NOR2X1_267/Y gnd AOI21X1_216/Y vdd AOI21X1
XAOI21X1_205 AOI21X1_205/A AOI21X1_205/B MUX2X1_96/S gnd OAI21X1_832/A vdd AOI21X1
XAOI21X1_227 BUFX4_395/Y NOR2X1_279/B NOR2X1_280/Y gnd AOI21X1_227/Y vdd AOI21X1
XAOI21X1_238 BUFX4_376/Y NOR2X1_289/B NOR2X1_293/Y gnd DFFPOSX1_64/D vdd AOI21X1
XAOI21X1_249 BUFX4_112/Y NOR2X1_315/B NOR2X1_314/Y gnd AOI21X1_249/Y vdd AOI21X1
XAOI22X1_32 AOI22X1_32/A AOI22X1_7/B BUFX4_159/Y MUX2X1_156/Y gnd AOI22X1_32/Y vdd
+ AOI22X1
XAOI22X1_10 MUX2X1_45/Y BUFX4_349/Y BUFX4_156/Y MUX2X1_48/Y gnd AOI22X1_10/Y vdd AOI22X1
XAOI22X1_21 MUX2X1_99/Y BUFX4_321/Y BUFX4_288/Y MUX2X1_102/Y gnd AOI22X1_21/Y vdd
+ AOI22X1
XAOI22X1_65 AOI22X1_65/A BUFX4_352/Y BUFX4_159/Y MUX2X1_312/Y gnd AOI22X1_65/Y vdd
+ AOI22X1
XAOI22X1_54 AOI22X1_54/A AOI22X1_9/A NAND2X1_5/B AOI22X1_54/D gnd AOI22X1_54/Y vdd
+ AOI22X1
XAOI22X1_43 AOI22X1_43/A BUFX4_321/Y BUFX4_288/Y AOI22X1_43/D gnd AOI22X1_43/Y vdd
+ AOI22X1
XOAI21X1_1411 BUFX4_457/Y BUFX4_390/Y INVX1_69/A gnd OAI21X1_1411/Y vdd OAI21X1
XOAI21X1_1422 BUFX4_279/Y NAND2X1_814/Y OAI21X1_1422/C gnd OAI21X1_1422/Y vdd OAI21X1
XOAI21X1_1400 BUFX4_305/Y NAND2X1_812/Y OAI21X1_1400/C gnd DFFPOSX1_124/D vdd OAI21X1
XOAI21X1_1466 NAND2X1_832/Y BUFX4_397/Y OAI21X1_1465/Y gnd OAI21X1_1466/Y vdd OAI21X1
XAOI22X1_76 MUX2X1_363/Y BUFX4_324/Y BUFX4_290/Y AOI22X1_76/D gnd AOI22X1_76/Y vdd
+ AOI22X1
XOAI21X1_1444 INVX1_198/Y NOR2X1_321/Y NAND2X1_819/Y gnd OAI21X1_1444/Y vdd OAI21X1
XOAI21X1_1455 INVX1_391/Y NOR2X1_331/Y NAND2X1_830/Y gnd OAI21X1_1455/Y vdd OAI21X1
XOAI21X1_1433 BUFX4_151/Y BUFX4_388/Y NAND2X1_487/B gnd OAI21X1_1433/Y vdd OAI21X1
XOAI21X1_1488 BUFX4_373/Y NAND2X1_833/Y OAI21X1_1487/Y gnd OAI21X1_1488/Y vdd OAI21X1
XOAI21X1_1477 BUFX4_417/Y INVX2_8/A NAND2X1_352/B gnd OAI21X1_1477/Y vdd OAI21X1
XOAI21X1_1499 NOR2X1_61/B BUFX4_94/Y INVX1_329/A gnd OAI21X1_1499/Y vdd OAI21X1
XFILL_24_6_0 gnd vdd FILL
XDFFPOSX1_1018 NOR2X1_232/A CLKBUF1_70/Y AOI21X1_188/Y gnd vdd DFFPOSX1
XDFFPOSX1_1007 NOR2X1_226/A CLKBUF1_85/Y AOI21X1_184/Y gnd vdd DFFPOSX1
XDFFPOSX1_1029 BUFX2_5/A CLKBUF1_44/Y NAND2X1_547/Y gnd vdd DFFPOSX1
XFILL_7_7_0 gnd vdd FILL
XFILL_15_6_0 gnd vdd FILL
XDFFPOSX1_308 INVX1_208/A CLKBUF1_32/Y OAI21X1_1641/Y gnd vdd DFFPOSX1
XDFFPOSX1_319 NAND2X1_637/B CLKBUF1_17/Y DFFPOSX1_319/D gnd vdd DFFPOSX1
XBUFX4_340 BUFX4_338/A gnd BUFX4_340/Y vdd BUFX4
XBUFX4_351 BUFX4_354/A gnd AOI22X1_7/B vdd BUFX4
XBUFX4_362 a[2] gnd BUFX4_362/Y vdd BUFX4
XBUFX4_373 INVX8_9/Y gnd BUFX4_373/Y vdd BUFX4
XFILL_40_1 gnd vdd FILL
XBUFX4_384 BUFX4_385/A gnd BUFX4_384/Y vdd BUFX4
XBUFX4_395 INVX8_6/Y gnd BUFX4_395/Y vdd BUFX4
XOAI21X1_906 INVX1_118/Y INVX8_1/A OAI21X1_906/C gnd MUX2X1_85/A vdd OAI21X1
XOAI21X1_928 INVX1_140/Y BUFX4_242/Y NAND2X1_356/Y gnd MUX2X1_101/A vdd OAI21X1
XOAI21X1_939 INVX1_151/Y BUFX4_264/Y NAND2X1_368/Y gnd MUX2X1_110/B vdd OAI21X1
XOAI21X1_917 INVX1_129/Y BUFX4_220/Y OAI21X1_917/C gnd MUX2X1_94/B vdd OAI21X1
XOAI21X1_1230 INVX1_442/Y BUFX4_252/Y NAND2X1_681/Y gnd MUX2X1_328/A vdd OAI21X1
XDFFPOSX1_842 NAND2X1_327/B CLKBUF1_7/Y OAI21X1_641/Y gnd vdd DFFPOSX1
XOAI21X1_1274 INVX1_486/Y BUFX4_241/Y NAND2X1_729/Y gnd MUX2X1_361/A vdd OAI21X1
XDFFPOSX1_820 INVX1_240/A CLKBUF1_37/Y OAI21X1_617/Y gnd vdd DFFPOSX1
XDFFPOSX1_831 NOR2X1_142/A CLKBUF1_37/Y AOI21X1_114/Y gnd vdd DFFPOSX1
XOAI21X1_1263 INVX1_475/Y BUFX4_219/Y NAND2X1_717/Y gnd MUX2X1_353/B vdd OAI21X1
XOAI21X1_1241 INVX1_453/Y BUFX4_274/Y NAND2X1_694/Y gnd MUX2X1_337/B vdd OAI21X1
XOAI21X1_1252 INVX1_464/Y BUFX4_197/Y NAND2X1_706/Y gnd MUX2X1_344/A vdd OAI21X1
XDFFPOSX1_853 INVX1_306/A CLKBUF1_80/Y OAI21X1_657/Y gnd vdd DFFPOSX1
XDFFPOSX1_875 NOR2X1_160/A CLKBUF1_57/Y AOI21X1_128/Y gnd vdd DFFPOSX1
XDFFPOSX1_864 NOR2X1_154/A CLKBUF1_81/Y AOI21X1_124/Y gnd vdd DFFPOSX1
XOAI21X1_1296 INVX1_508/Y MUX2X1_11/S NAND2X1_752/Y gnd MUX2X1_377/A vdd OAI21X1
XOAI21X1_1285 INVX1_497/Y BUFX4_263/Y NAND2X1_741/Y gnd MUX2X1_370/B vdd OAI21X1
XDFFPOSX1_897 MUX2X1_15/B CLKBUF1_101/Y OAI21X1_676/Y gnd vdd DFFPOSX1
XDFFPOSX1_886 INVX1_372/A CLKBUF1_13/Y OAI21X1_672/Y gnd vdd DFFPOSX1
XFILL_47_5_0 gnd vdd FILL
XFILL_30_4_0 gnd vdd FILL
XDFFPOSX1_116 INVX1_196/A CLKBUF1_42/Y OAI21X1_1384/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 NAND2X1_624/B CLKBUF1_55/Y DFFPOSX1_127/D gnd vdd DFFPOSX1
XDFFPOSX1_105 NOR2X1_312/A CLKBUF1_55/Y AOI21X1_247/Y gnd vdd DFFPOSX1
XDFFPOSX1_149 INVX1_262/A CLKBUF1_63/Y OAI21X1_1445/Y gnd vdd DFFPOSX1
XDFFPOSX1_138 NAND2X1_280/B CLKBUF1_61/Y DFFPOSX1_138/D gnd vdd DFFPOSX1
XNAND2X1_208 BUFX4_427/Y NOR2X1_228/Y gnd OAI21X1_798/C vdd NAND2X1
XNAND2X1_219 NOR2X1_244/Y OAI21X1_807/Y gnd NAND3X1_2/B vdd NAND2X1
XFILL_38_5_0 gnd vdd FILL
XBUFX4_181 BUFX4_25/Y gnd MUX2X1_2/S vdd BUFX4
XBUFX4_170 BUFX4_168/A gnd INVX4_3/A vdd BUFX4
XNOR2X1_230 BUFX4_438/Y NOR2X1_32/B gnd NOR2X1_236/B vdd NOR2X1
XNOR2X1_241 a[3] INVX1_9/Y gnd BUFX4_321/A vdd NOR2X1
XNOR2X1_252 a[6] INVX1_13/Y gnd NAND2X1_5/B vdd NOR2X1
XBUFX4_192 BUFX4_25/Y gnd BUFX4_192/Y vdd BUFX4
XNOR2X1_285 NAND3X1_7/Y OR2X2_1/Y gnd NOR2X1_289/B vdd NOR2X1
XNOR2X1_274 NAND3X1_7/Y OAI22X1_3/A gnd NOR2X1_274/Y vdd NOR2X1
XNOR2X1_263 NOR2X1_263/A NOR2X1_256/B gnd NOR2X1_263/Y vdd NOR2X1
XNOR2X1_296 INVX4_2/Y NOR2X1_264/B gnd INVX8_12/A vdd NOR2X1
XOAI21X1_714 INVX1_119/Y NOR2X1_189/B OAI21X1_714/C gnd OAI21X1_714/Y vdd OAI21X1
XOAI21X1_703 BUFX4_146/Y INVX1_5/A NAND2X1_676/B gnd OAI21X1_704/C vdd OAI21X1
XFILL_21_4_0 gnd vdd FILL
XOAI21X1_725 INVX1_376/Y NOR2X1_199/Y OAI21X1_725/C gnd OAI21X1_725/Y vdd OAI21X1
XOAI21X1_736 BUFX4_455/Y BUFX4_443/Y INVX1_313/A gnd OAI21X1_737/C vdd OAI21X1
XOAI21X1_747 BUFX4_419/Y OAI21X1_757/B OAI21X1_747/C gnd OAI21X1_747/Y vdd OAI21X1
XOAI21X1_758 NOR2X1_72/B BUFX4_443/Y NAND2X1_749/B gnd OAI21X1_759/C vdd OAI21X1
XOAI21X1_769 BUFX4_400/Y OAI21X1_761/B OAI21X1_769/C gnd OAI21X1_769/Y vdd OAI21X1
XMUX2X1_203 MUX2X1_203/A MUX2X1_203/B BUFX4_82/Y gnd MUX2X1_203/Y vdd MUX2X1
XMUX2X1_214 MUX2X1_214/A MUX2X1_214/B BUFX4_2/Y gnd MUX2X1_214/Y vdd MUX2X1
XOAI21X1_1082 INVX1_294/Y BUFX4_253/Y NAND2X1_522/Y gnd MUX2X1_217/A vdd OAI21X1
XMUX2X1_236 MUX2X1_236/A MUX2X1_236/B BUFX4_3/Y gnd MUX2X1_236/Y vdd MUX2X1
XMUX2X1_225 MUX2X1_224/Y MUX2X1_225/B BUFX4_364/Y gnd AOI22X1_47/A vdd MUX2X1
XOAI21X1_1071 INVX1_283/Y BUFX4_231/Y NAND2X1_510/Y gnd MUX2X1_209/B vdd OAI21X1
XDFFPOSX1_650 NOR2X1_74/A CLKBUF1_100/Y AOI21X1_58/Y gnd vdd DFFPOSX1
XMUX2X1_247 MUX2X1_247/A MUX2X1_247/B BUFX4_81/Y gnd MUX2X1_249/B vdd MUX2X1
XOAI21X1_1060 INVX1_272/Y BUFX4_209/Y NAND2X1_499/Y gnd MUX2X1_200/A vdd OAI21X1
XOAI21X1_1093 INVX1_305/Y BUFX4_275/Y NAND2X1_534/Y gnd MUX2X1_226/B vdd OAI21X1
XDFFPOSX1_661 INVX1_294/A CLKBUF1_38/Y OAI21X1_426/Y gnd vdd DFFPOSX1
XDFFPOSX1_683 NAND2X1_385/B CLKBUF1_45/Y OAI21X1_470/Y gnd vdd DFFPOSX1
XDFFPOSX1_672 NAND2X1_729/B CLKBUF1_58/Y OAI21X1_448/Y gnd vdd DFFPOSX1
XMUX2X1_258 MUX2X1_258/A MUX2X1_256/Y BUFX4_364/Y gnd AOI22X1_53/D vdd MUX2X1
XMUX2X1_269 MUX2X1_269/A MUX2X1_269/B BUFX4_81/Y gnd MUX2X1_270/A vdd MUX2X1
XNAND2X1_720 BUFX4_222/Y NAND2X1_720/B gnd NAND2X1_720/Y vdd NAND2X1
XDFFPOSX1_694 INVX1_360/A CLKBUF1_99/Y OAI21X1_492/Y gnd vdd DFFPOSX1
XNAND2X1_731 BUFX4_244/Y NAND2X1_731/B gnd NAND2X1_731/Y vdd NAND2X1
XNAND2X1_764 MUX2X1_12/S AOI22X1_1/C gnd NOR2X1_255/A vdd NAND2X1
XNAND2X1_753 AOI22X1_77/Y AOI22X1_78/Y gnd AOI22X1_79/D vdd NAND2X1
XNAND2X1_742 BUFX4_264/Y NOR2X1_154/A gnd NAND2X1_742/Y vdd NAND2X1
XNAND2X1_797 BUFX4_142/Y NOR2X1_297/Y gnd NAND2X1_797/Y vdd NAND2X1
XNAND2X1_786 NAND2X1_9/A NOR2X1_284/Y gnd NAND2X1_786/Y vdd NAND2X1
XNAND2X1_775 BUFX4_163/Y NOR2X1_274/Y gnd NAND2X1_775/Y vdd NAND2X1
XFILL_4_5_0 gnd vdd FILL
XFILL_29_5_0 gnd vdd FILL
XFILL_12_4_0 gnd vdd FILL
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XBUFX4_10 clk gnd BUFX4_10/Y vdd BUFX4
XBUFX4_32 BUFX4_75/Y gnd BUFX4_32/Y vdd BUFX4
XBUFX4_43 BUFX4_41/A gnd BUFX4_43/Y vdd BUFX4
XBUFX4_21 BUFX4_70/Y gnd BUFX4_21/Y vdd BUFX4
XBUFX4_65 BUFX4_64/A gnd INVX1_5/A vdd BUFX4
XBUFX4_87 BUFX4_84/A gnd BUFX4_87/Y vdd BUFX4
XBUFX4_54 BUFX4_52/A gnd BUFX4_54/Y vdd BUFX4
XBUFX4_76 a[1] gnd BUFX4_52/A vdd BUFX4
XBUFX4_98 INVX8_7/Y gnd BUFX4_98/Y vdd BUFX4
XINVX8_13 INVX8_13/A gnd BUFX4_84/A vdd INVX8
XOAI21X1_511 BUFX4_414/Y BUFX4_342/Y NAND2X1_731/B gnd OAI21X1_511/Y vdd OAI21X1
XOAI21X1_500 BUFX4_419/Y NAND2X1_97/Y OAI21X1_500/C gnd OAI21X1_500/Y vdd OAI21X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XOAI21X1_522 BUFX4_396/Y NAND2X1_99/Y OAI21X1_522/C gnd OAI21X1_522/Y vdd OAI21X1
XOAI21X1_566 INVX1_364/Y NOR2X1_101/Y NAND2X1_122/Y gnd OAI21X1_566/Y vdd OAI21X1
XOAI21X1_555 INVX1_171/Y NOR2X1_91/Y NAND2X1_111/Y gnd OAI21X1_555/Y vdd OAI21X1
XOAI21X1_533 BUFX4_148/Y BUFX4_295/Y NAND2X1_387/B gnd OAI21X1_534/C vdd OAI21X1
XOAI21X1_544 BUFX4_372/Y OAI21X1_544/B OAI21X1_543/Y gnd OAI21X1_544/Y vdd OAI21X1
XOAI21X1_588 BUFX4_425/Y OAI21X1_590/B OAI21X1_588/C gnd OAI21X1_588/Y vdd OAI21X1
XOAI21X1_577 NOR2X1_1/B INVX1_3/A INVX1_301/A gnd OAI21X1_578/C vdd OAI21X1
XOAI21X1_599 BUFX4_148/Y INVX1_3/A NAND2X1_737/B gnd OAI21X1_599/Y vdd OAI21X1
XDFFPOSX1_480 NOR2X1_20/A CLKBUF1_40/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_491 NOR2X1_25/A CLKBUF1_24/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XNAND2X1_572 BUFX4_245/Y OAI21X1_59/C gnd NAND2X1_572/Y vdd NAND2X1
XNAND2X1_561 BUFX4_225/Y NOR2X1_347/A gnd NAND2X1_561/Y vdd NAND2X1
XNAND2X1_550 BUFX4_203/Y NOR2X1_281/A gnd NAND2X1_550/Y vdd NAND2X1
XNAND2X1_594 BUFX4_188/Y NAND2X1_594/B gnd NAND2X1_594/Y vdd NAND2X1
XNAND2X1_583 BUFX4_265/Y NOR2X1_48/A gnd NAND2X1_583/Y vdd NAND2X1
XFILL_45_8_1 gnd vdd FILL
XFILL_44_3_0 gnd vdd FILL
XFILL_9_1 gnd vdd FILL
XFILL_35_3_0 gnd vdd FILL
XFILL_36_8_1 gnd vdd FILL
XFILL_2_8_1 gnd vdd FILL
XFILL_27_8_1 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XFILL_10_7_1 gnd vdd FILL
XOAI21X1_341 BUFX4_85/Y BUFX4_381/Y NAND2X1_656/B gnd OAI21X1_342/C vdd OAI21X1
XOAI21X1_330 BUFX4_123/Y NAND2X1_78/Y OAI21X1_330/C gnd OAI21X1_330/Y vdd OAI21X1
XOAI21X1_374 BUFX4_283/Y NAND2X1_80/Y OAI21X1_373/Y gnd OAI21X1_374/Y vdd OAI21X1
XOAI21X1_363 BUFX4_370/Y INVX2_3/A NAND2X1_312/B gnd OAI21X1_364/C vdd OAI21X1
XOAI21X1_352 BUFX4_303/Y NAND2X1_79/Y OAI21X1_351/Y gnd OAI21X1_352/Y vdd OAI21X1
XOAI21X1_396 BUFX4_421/Y NAND2X1_82/Y OAI21X1_396/C gnd OAI21X1_396/Y vdd OAI21X1
XOAI21X1_385 BUFX4_172/Y BUFX4_384/Y INVX1_292/A gnd OAI21X1_386/C vdd OAI21X1
XINVX1_405 INVX1_405/A gnd INVX1_405/Y vdd INVX1
XINVX1_416 INVX1_416/A gnd INVX1_416/Y vdd INVX1
XINVX1_449 INVX1_449/A gnd INVX1_449/Y vdd INVX1
XINVX1_438 INVX1_438/A gnd INVX1_438/Y vdd INVX1
XINVX1_427 INVX1_427/A gnd INVX1_427/Y vdd INVX1
XFILL_9_4_0 gnd vdd FILL
XNAND2X1_380 MUX2X1_11/S OAI21X1_333/C gnd NAND2X1_380/Y vdd NAND2X1
XNAND2X1_391 AOI22X1_25/Y AOI22X1_26/Y gnd AOI22X1_29/A vdd NAND2X1
XFILL_18_8_1 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XOAI21X1_1604 NOR2X1_2/B BUFX4_345/Y NAND2X1_289/B gnd OAI21X1_1604/Y vdd OAI21X1
XOAI21X1_1615 BUFX4_279/Y NAND2X1_843/Y OAI21X1_1614/Y gnd OAI21X1_1615/Y vdd OAI21X1
XOAI21X1_1648 BUFX4_168/Y BUFX4_343/Y INVX1_464/A gnd OAI21X1_1649/C vdd OAI21X1
XOAI21X1_1626 INVX1_18/Y NOR2X1_368/Y NAND2X1_852/Y gnd OAI21X1_1626/Y vdd OAI21X1
XOAI21X1_1637 NAND2X1_860/Y BUFX4_420/Y OAI21X1_1637/C gnd OAI21X1_1637/Y vdd OAI21X1
XOAI21X1_1659 BUFX4_399/Y NAND2X1_861/Y OAI21X1_1658/Y gnd OAI21X1_1659/Y vdd OAI21X1
XFILL_41_1_0 gnd vdd FILL
XFILL_42_6_1 gnd vdd FILL
XAOI22X1_3 AOI22X1_3/A BUFX4_349/Y BUFX4_156/Y NAND3X1_2/Y gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_182 BUFX4_282/Y NAND2X1_21/Y OAI21X1_181/Y gnd OAI21X1_182/Y vdd OAI21X1
XOAI21X1_171 BUFX4_457/Y BUFX4_134/Y INVX1_89/A gnd OAI21X1_171/Y vdd OAI21X1
XOAI21X1_160 BUFX4_297/Y NAND2X1_19/Y OAI21X1_160/C gnd OAI21X1_160/Y vdd OAI21X1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XOAI21X1_193 BUFX4_147/Y INVX1_1/A NAND2X1_508/B gnd OAI21X1_193/Y vdd OAI21X1
XINVX1_213 INVX1_213/A gnd INVX1_213/Y vdd INVX1
XINVX1_235 INVX1_235/A gnd INVX1_235/Y vdd INVX1
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XINVX1_257 INVX1_257/A gnd INVX1_257/Y vdd INVX1
XINVX1_246 INVX1_246/A gnd INVX1_246/Y vdd INVX1
XINVX1_268 INVX1_268/A gnd INVX1_268/Y vdd INVX1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XNAND2X1_24 BUFX4_450/Y NOR2X1_11/Y gnd NAND2X1_24/Y vdd NAND2X1
XNAND2X1_13 BUFX4_427/Y NOR2X1_1/Y gnd NAND2X1_13/Y vdd NAND2X1
XNAND2X1_68 BUFX4_157/Y AOI22X1_9/D gnd BUFX4_385/A vdd NAND2X1
XNAND2X1_46 BUFX4_430/Y NOR2X1_31/Y gnd NAND2X1_46/Y vdd NAND2X1
XNAND2X1_35 INVX8_6/A NOR2X1_21/Y gnd NAND2X1_35/Y vdd NAND2X1
XNAND2X1_57 BUFX4_431/Y NOR2X1_41/Y gnd NAND2X1_57/Y vdd NAND2X1
XNAND2X1_79 INVX2_3/Y INVX8_14/A gnd NAND2X1_79/Y vdd NAND2X1
XFILL_32_1_0 gnd vdd FILL
XFILL_33_6_1 gnd vdd FILL
XAOI21X1_206 NAND2X1_252/Y AOI21X1_206/B INVX2_6/Y gnd OAI21X1_832/B vdd AOI21X1
XAOI21X1_239 BUFX4_129/Y NOR2X1_303/B NOR2X1_300/Y gnd AOI21X1_239/Y vdd AOI21X1
XAOI21X1_217 BUFX4_115/Y NOR2X1_265/Y NOR2X1_268/Y gnd DFFPOSX1_43/D vdd AOI21X1
XAOI21X1_228 BUFX4_96/Y NOR2X1_279/B NOR2X1_281/Y gnd DFFPOSX1_22/D vdd AOI21X1
XAOI22X1_33 AOI22X1_33/A BUFX4_320/Y INVX1_11/A MUX2X1_162/Y gnd AOI22X1_33/Y vdd
+ AOI22X1
XAOI22X1_11 MUX2X1_51/Y BUFX4_323/Y AOI22X1_6/C MUX2X1_54/Y gnd AOI22X1_11/Y vdd AOI22X1
XAOI22X1_22 AOI22X1_22/A BUFX4_350/Y AOI22X1_7/C MUX2X1_108/Y gnd AOI22X1_22/Y vdd
+ AOI22X1
XAOI22X1_66 MUX2X1_315/Y BUFX4_322/Y BUFX4_292/Y AOI22X1_66/D gnd AOI22X1_66/Y vdd
+ AOI22X1
XAOI22X1_55 AOI22X1_55/A BUFX4_352/Y BUFX4_159/Y MUX2X1_264/Y gnd AOI22X1_55/Y vdd
+ AOI22X1
XAOI22X1_44 AOI22X1_44/A AOI22X1_9/A NAND2X1_5/B AOI22X1_44/D gnd AOI22X1_44/Y vdd
+ AOI22X1
XOAI21X1_1412 BUFX4_420/Y NAND2X1_814/Y OAI21X1_1411/Y gnd OAI21X1_1412/Y vdd OAI21X1
XOAI21X1_1423 BUFX4_460/Y BUFX4_388/Y INVX1_453/A gnd OAI21X1_1423/Y vdd OAI21X1
XOAI21X1_1401 BUFX4_416/Y BUFX4_463/Y NAND2X1_486/B gnd OAI21X1_1401/Y vdd OAI21X1
XAOI22X1_77 AOI22X1_77/A INVX1_6/A INVX1_8/A AOI22X1_77/D gnd AOI22X1_77/Y vdd AOI22X1
XOAI21X1_1445 INVX1_262/Y NOR2X1_321/Y NAND2X1_820/Y gnd OAI21X1_1445/Y vdd OAI21X1
XOAI21X1_1456 INVX1_455/Y NOR2X1_331/Y NAND2X1_831/Y gnd OAI21X1_1456/Y vdd OAI21X1
XOAI21X1_1434 BUFX4_397/Y NAND2X1_815/Y OAI21X1_1433/Y gnd OAI21X1_1434/Y vdd OAI21X1
XOAI21X1_1467 BUFX4_167/Y BUFX4_393/Y INVX1_328/A gnd OAI21X1_1468/C vdd OAI21X1
XOAI21X1_1478 BUFX4_112/Y NAND2X1_833/Y OAI21X1_1477/Y gnd DFFPOSX1_187/D vdd OAI21X1
XOAI21X1_1489 BUFX4_462/Y BUFX4_89/Y MUX2X1_29/B gnd OAI21X1_1489/Y vdd OAI21X1
XFILL_24_6_1 gnd vdd FILL
XFILL_23_1_0 gnd vdd FILL
XDFFPOSX1_1008 NOR2X1_227/A CLKBUF1_85/Y AOI21X1_185/Y gnd vdd DFFPOSX1
XDFFPOSX1_1019 NOR2X1_233/A CLKBUF1_3/Y AOI21X1_189/Y gnd vdd DFFPOSX1
XFILL_7_7_1 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XFILL_15_6_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_309 INVX1_272/A CLKBUF1_39/Y OAI21X1_1643/Y gnd vdd DFFPOSX1
XBUFX4_330 d[5] gnd BUFX4_330/Y vdd BUFX4
XBUFX4_341 BUFX4_338/A gnd BUFX4_341/Y vdd BUFX4
XBUFX4_352 BUFX4_354/A gnd BUFX4_352/Y vdd BUFX4
XBUFX4_363 a[2] gnd BUFX4_363/Y vdd BUFX4
XBUFX4_385 BUFX4_385/A gnd BUFX4_385/Y vdd BUFX4
XBUFX4_396 INVX8_6/Y gnd BUFX4_396/Y vdd BUFX4
XBUFX4_374 INVX8_9/Y gnd BUFX4_374/Y vdd BUFX4
XOAI21X1_907 INVX1_119/Y BUFX4_200/Y NAND2X1_333/Y gnd MUX2X1_86/B vdd OAI21X1
XOAI21X1_918 INVX1_130/Y BUFX4_222/Y OAI21X1_918/C gnd MUX2X1_94/A vdd OAI21X1
XOAI21X1_929 INVX1_141/Y BUFX4_244/Y NAND2X1_358/Y gnd MUX2X1_103/B vdd OAI21X1
XOAI21X1_1231 INVX1_443/Y BUFX4_254/Y NAND2X1_682/Y gnd MUX2X1_329/B vdd OAI21X1
XOAI21X1_1220 INVX1_432/Y BUFX4_232/Y NAND2X1_671/Y gnd MUX2X1_320/A vdd OAI21X1
XDFFPOSX1_821 INVX1_304/A CLKBUF1_21/Y OAI21X1_618/Y gnd vdd DFFPOSX1
XOAI21X1_1253 INVX1_465/Y BUFX4_199/Y NAND2X1_707/Y gnd MUX2X1_346/B vdd OAI21X1
XDFFPOSX1_832 NOR2X1_143/A CLKBUF1_69/Y AOI21X1_115/Y gnd vdd DFFPOSX1
XOAI21X1_1264 INVX1_476/Y BUFX4_221/Y NAND2X1_718/Y gnd MUX2X1_353/A vdd OAI21X1
XDFFPOSX1_810 NOR2X1_126/A CLKBUF1_74/Y AOI21X1_100/Y gnd vdd DFFPOSX1
XOAI21X1_1242 INVX1_454/Y BUFX4_276/Y NAND2X1_695/Y gnd MUX2X1_337/A vdd OAI21X1
XOAI21X1_1275 INVX1_487/Y BUFX4_243/Y NAND2X1_730/Y gnd MUX2X1_362/B vdd OAI21X1
XOAI21X1_1297 INVX1_33/Y NOR2X1_254/Y NAND2X1_756/Y gnd DFFPOSX1_25/D vdd OAI21X1
XDFFPOSX1_865 MUX2X1_11/B CLKBUF1_27/Y AOI21X1_125/Y gnd vdd DFFPOSX1
XOAI21X1_1286 INVX1_498/Y BUFX4_265/Y NAND2X1_742/Y gnd MUX2X1_370/A vdd OAI21X1
XDFFPOSX1_854 INVX1_370/A CLKBUF1_54/Y OAI21X1_658/Y gnd vdd DFFPOSX1
XDFFPOSX1_843 OAI21X1_642/C CLKBUF1_7/Y OAI21X1_643/Y gnd vdd DFFPOSX1
XDFFPOSX1_876 NOR2X1_161/A CLKBUF1_15/Y AOI21X1_129/Y gnd vdd DFFPOSX1
XDFFPOSX1_898 INVX1_117/A CLKBUF1_21/Y OAI21X1_678/Y gnd vdd DFFPOSX1
XDFFPOSX1_887 INVX1_436/A CLKBUF1_84/Y OAI21X1_673/Y gnd vdd DFFPOSX1
XFILL_47_5_1 gnd vdd FILL
XFILL_46_0_0 gnd vdd FILL
XFILL_30_4_1 gnd vdd FILL
XDFFPOSX1_117 INVX1_260/A CLKBUF1_42/Y OAI21X1_1386/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 NAND2X1_693/B CLKBUF1_20/Y OAI21X1_1408/Y gnd vdd DFFPOSX1
XDFFPOSX1_106 NOR2X1_313/A CLKBUF1_53/Y AOI21X1_248/Y gnd vdd DFFPOSX1
XDFFPOSX1_139 NAND2X1_349/B CLKBUF1_102/Y DFFPOSX1_139/D gnd vdd DFFPOSX1
XNAND2X1_209 BUFX4_196/Y NOR2X1_244/Y gnd NOR2X1_275/B vdd NAND2X1
XFILL_37_0_0 gnd vdd FILL
XFILL_38_5_1 gnd vdd FILL
XBUFX4_171 BUFX4_168/A gnd BUFX4_171/Y vdd BUFX4
XBUFX4_182 BUFX4_29/Y gnd MUX2X1_4/S vdd BUFX4
XBUFX4_160 BUFX4_155/A gnd INVX1_8/A vdd BUFX4
XNOR2X1_231 MUX2X1_26/A NOR2X1_236/B gnd NOR2X1_231/Y vdd NOR2X1
XNOR2X1_220 MUX2X1_25/A NOR2X1_222/B gnd NOR2X1_220/Y vdd NOR2X1
XNOR2X1_242 INVX1_9/Y INVX1_7/Y gnd BUFX4_288/A vdd NOR2X1
XBUFX4_193 BUFX4_25/Y gnd BUFX4_193/Y vdd BUFX4
XNOR2X1_264 NAND3X1_7/Y NOR2X1_264/B gnd NOR2X1_264/Y vdd NOR2X1
XNOR2X1_275 NAND3X1_7/Y NOR2X1_275/B gnd NOR2X1_279/B vdd NOR2X1
XNOR2X1_253 a[5] INVX1_12/Y gnd AOI22X1_9/D vdd NOR2X1
XNOR2X1_286 NOR2X1_286/A NOR2X1_289/B gnd NOR2X1_286/Y vdd NOR2X1
XNOR2X1_297 BUFX4_463/Y NOR2X1_41/B gnd NOR2X1_297/Y vdd NOR2X1
XOAI21X1_715 INVX1_183/Y NOR2X1_189/B OAI21X1_715/C gnd OAI21X1_715/Y vdd OAI21X1
XOAI21X1_704 BUFX4_285/Y OAI21X1_704/B OAI21X1_704/C gnd OAI21X1_704/Y vdd OAI21X1
XFILL_21_4_1 gnd vdd FILL
XOAI21X1_726 INVX1_440/Y NOR2X1_199/Y OAI21X1_726/C gnd OAI21X1_726/Y vdd OAI21X1
XOAI21X1_748 NOR2X1_72/B BUFX4_442/Y NAND2X1_404/B gnd OAI21X1_749/C vdd OAI21X1
XOAI21X1_737 BUFX4_400/Y OAI21X1_729/B OAI21X1_737/C gnd OAI21X1_737/Y vdd OAI21X1
XOAI21X1_759 BUFX4_378/Y OAI21X1_757/B OAI21X1_759/C gnd OAI21X1_759/Y vdd OAI21X1
XMUX2X1_204 MUX2X1_203/Y MUX2X1_202/Y BUFX4_357/Y gnd MUX2X1_204/Y vdd MUX2X1
XMUX2X1_226 MUX2X1_226/A MUX2X1_226/B BUFX4_82/Y gnd MUX2X1_228/B vdd MUX2X1
XOAI21X1_1061 INVX1_273/Y BUFX4_211/Y NAND2X1_500/Y gnd MUX2X1_202/B vdd OAI21X1
XDFFPOSX1_640 OAI21X1_407/C CLKBUF1_6/Y OAI21X1_408/Y gnd vdd DFFPOSX1
XMUX2X1_215 MUX2X1_215/A MUX2X1_215/B BUFX4_33/Y gnd MUX2X1_215/Y vdd MUX2X1
XMUX2X1_237 MUX2X1_236/Y MUX2X1_235/Y BUFX4_357/Y gnd MUX2X1_237/Y vdd MUX2X1
XOAI21X1_1072 INVX1_284/Y BUFX4_233/Y NAND2X1_511/Y gnd MUX2X1_209/A vdd OAI21X1
XOAI21X1_1050 INVX1_262/Y BUFX4_189/Y NAND2X1_488/Y gnd MUX2X1_193/A vdd OAI21X1
XOAI21X1_1094 INVX1_306/Y BUFX4_277/Y NAND2X1_535/Y gnd MUX2X1_226/A vdd OAI21X1
XDFFPOSX1_673 INVX1_55/A CLKBUF1_38/Y OAI21X1_450/Y gnd vdd DFFPOSX1
XDFFPOSX1_684 NAND2X1_454/B CLKBUF1_45/Y OAI21X1_472/Y gnd vdd DFFPOSX1
XDFFPOSX1_662 INVX1_358/A CLKBUF1_96/Y OAI21X1_428/Y gnd vdd DFFPOSX1
XOAI21X1_1083 INVX1_295/Y BUFX4_255/Y NAND2X1_523/Y gnd MUX2X1_218/B vdd OAI21X1
XDFFPOSX1_651 NOR2X1_75/A CLKBUF1_88/Y AOI21X1_59/Y gnd vdd DFFPOSX1
XMUX2X1_259 MUX2X1_259/A MUX2X1_259/B BUFX4_4/Y gnd MUX2X1_261/B vdd MUX2X1
XMUX2X1_248 MUX2X1_248/A MUX2X1_248/B BUFX4_82/Y gnd MUX2X1_249/A vdd MUX2X1
XDFFPOSX1_695 INVX1_424/A CLKBUF1_38/Y OAI21X1_494/Y gnd vdd DFFPOSX1
XNAND2X1_710 BUFX4_204/Y OAI21X1_63/C gnd NAND2X1_710/Y vdd NAND2X1
XNAND2X1_721 BUFX4_224/Y NOR2X1_50/A gnd NAND2X1_721/Y vdd NAND2X1
XNAND2X1_754 AOI22X1_74/Y AOI22X1_79/Y gnd NAND2X1_754/Y vdd NAND2X1
XNAND2X1_743 BUFX4_266/Y NOR2X1_165/A gnd NAND2X1_743/Y vdd NAND2X1
XNAND2X1_732 BUFX4_246/Y OAI21X1_543/C gnd NAND2X1_732/Y vdd NAND2X1
XNAND2X1_765 INVX8_1/Y AOI22X1_1/B gnd NOR2X1_264/B vdd NAND2X1
XNAND2X1_776 BUFX4_453/Y NOR2X1_274/Y gnd NAND2X1_776/Y vdd NAND2X1
XNAND2X1_787 BUFX4_444/Y NOR2X1_284/Y gnd NAND2X1_787/Y vdd NAND2X1
XFILL_4_5_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_29_5_1 gnd vdd FILL
XNAND2X1_798 BUFX4_445/Y NOR2X1_297/Y gnd NAND2X1_798/Y vdd NAND2X1
XFILL_3_0_0 gnd vdd FILL
XFILL_12_4_1 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XBUFX4_11 clk gnd BUFX4_11/Y vdd BUFX4
XBUFX4_33 BUFX4_75/Y gnd BUFX4_33/Y vdd BUFX4
XBUFX4_44 BUFX4_71/Y gnd BUFX4_44/Y vdd BUFX4
XBUFX4_22 BUFX4_70/Y gnd BUFX4_22/Y vdd BUFX4
XBUFX4_66 BUFX4_64/A gnd BUFX4_66/Y vdd BUFX4
XBUFX4_77 a[1] gnd BUFX4_8/A vdd BUFX4
XBUFX4_55 BUFX4_52/A gnd BUFX4_55/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_88 BUFX4_84/A gnd BUFX4_88/Y vdd BUFX4
XBUFX4_99 INVX8_7/Y gnd BUFX4_99/Y vdd BUFX4
XINVX8_14 INVX8_14/A gnd INVX8_14/Y vdd INVX8
XOAI21X1_512 BUFX4_377/Y NAND2X1_97/Y OAI21X1_511/Y gnd OAI21X1_512/Y vdd OAI21X1
XOAI21X1_501 BUFX4_414/Y NOR2X1_72/A OAI21X1_501/C gnd OAI21X1_501/Y vdd OAI21X1
XINVX1_9 a[4] gnd INVX1_9/Y vdd INVX1
XOAI21X1_523 NOR2X1_1/B BUFX4_293/Y INVX1_361/A gnd OAI21X1_524/C vdd OAI21X1
XOAI21X1_534 BUFX4_110/Y OAI21X1_544/B OAI21X1_534/C gnd OAI21X1_534/Y vdd OAI21X1
XOAI21X1_556 INVX1_235/Y NOR2X1_91/Y OAI21X1_556/C gnd OAI21X1_556/Y vdd OAI21X1
XOAI21X1_545 INVX1_58/Y NOR2X1_81/Y OAI21X1_545/C gnd OAI21X1_545/Y vdd OAI21X1
XOAI21X1_567 INVX1_428/Y NOR2X1_101/Y NAND2X1_123/Y gnd OAI21X1_567/Y vdd OAI21X1
XOAI21X1_578 BUFX4_396/Y OAI21X1_584/B OAI21X1_578/C gnd OAI21X1_578/Y vdd OAI21X1
XOAI21X1_589 BUFX4_148/Y BUFX4_107/Y NAND2X1_392/B gnd OAI21X1_590/C vdd OAI21X1
XDFFPOSX1_470 INVX1_346/A CLKBUF1_3/Y OAI21X1_206/Y gnd vdd DFFPOSX1
XDFFPOSX1_492 NOR2X1_26/A CLKBUF1_31/Y AOI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_481 INVX1_30/A CLKBUF1_2/Y OAI21X1_209/Y gnd vdd DFFPOSX1
XNAND2X1_562 BUFX4_227/Y NOR2X1_355/A gnd NAND2X1_562/Y vdd NAND2X1
XNAND2X1_540 MUX2X1_12/S NOR2X1_195/A gnd NAND2X1_540/Y vdd NAND2X1
XNAND2X1_551 BUFX4_205/Y NOR2X1_291/A gnd NAND2X1_551/Y vdd NAND2X1
XNAND2X1_595 BUFX4_190/Y NOR2X1_88/A gnd NAND2X1_595/Y vdd NAND2X1
XNAND2X1_573 BUFX4_247/Y NOR2X1_8/A gnd NAND2X1_573/Y vdd NAND2X1
XNAND2X1_584 BUFX4_267/Y NOR2X1_58/A gnd NAND2X1_584/Y vdd NAND2X1
XFILL_44_3_1 gnd vdd FILL
XFILL_35_3_1 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XFILL_26_3_1 gnd vdd FILL
XOAI21X1_320 BUFX4_300/Y NAND2X1_77/Y OAI21X1_320/C gnd OAI21X1_320/Y vdd OAI21X1
XOAI21X1_331 BUFX4_88/Y BUFX4_385/Y NAND2X1_311/B gnd OAI21X1_331/Y vdd OAI21X1
XOAI21X1_342 BUFX4_284/Y NAND2X1_78/Y OAI21X1_342/C gnd OAI21X1_342/Y vdd OAI21X1
XOAI21X1_353 BUFX4_307/Y BUFX4_387/Y INVX1_291/A gnd OAI21X1_354/C vdd OAI21X1
XOAI21X1_364 BUFX4_421/Y NAND2X1_80/Y OAI21X1_364/C gnd OAI21X1_364/Y vdd OAI21X1
XOAI21X1_397 BUFX4_415/Y NOR2X1_61/A OAI21X1_397/C gnd OAI21X1_398/C vdd OAI21X1
XOAI21X1_375 NOR2X1_22/B BUFX4_384/Y OAI21X1_375/C gnd OAI21X1_375/Y vdd OAI21X1
XOAI21X1_386 NAND2X1_81/Y BUFX4_398/Y OAI21X1_386/C gnd OAI21X1_386/Y vdd OAI21X1
XINVX1_417 INVX1_417/A gnd INVX1_417/Y vdd INVX1
XINVX1_406 INVX1_406/A gnd INVX1_406/Y vdd INVX1
XINVX1_439 INVX1_439/A gnd INVX1_439/Y vdd INVX1
XINVX1_428 INVX1_428/A gnd INVX1_428/Y vdd INVX1
XFILL_9_4_1 gnd vdd FILL
XNAND2X1_381 BUFX4_188/Y NAND2X1_381/B gnd NAND2X1_381/Y vdd NAND2X1
XNAND2X1_370 BUFX4_267/Y OAI21X1_189/C gnd NAND2X1_370/Y vdd NAND2X1
XNAND2X1_392 BUFX4_208/Y NAND2X1_392/B gnd NAND2X1_392/Y vdd NAND2X1
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_1605 BUFX4_423/Y NAND2X1_843/Y OAI21X1_1604/Y gnd OAI21X1_1605/Y vdd OAI21X1
XOAI21X1_1638 BUFX4_168/Y BUFX4_343/Y INVX1_144/A gnd OAI21X1_1638/Y vdd OAI21X1
XOAI21X1_1627 INVX1_79/Y NOR2X1_368/Y NAND2X1_853/Y gnd OAI21X1_1627/Y vdd OAI21X1
XOAI21X1_1616 BUFX4_150/Y BUFX4_346/Y NAND2X1_703/B gnd OAI21X1_1617/C vdd OAI21X1
XOAI21X1_1649 NAND2X1_860/Y BUFX4_373/Y OAI21X1_1649/C gnd DFFPOSX1_312/D vdd OAI21X1
XFILL_41_1_1 gnd vdd FILL
XAOI22X1_4 AOI22X1_4/A AOI22X1_1/B AOI22X1_1/C AOI22X1_4/D gnd NAND3X1_3/C vdd AOI22X1
XOAI21X1_172 BUFX4_423/Y NAND2X1_21/Y OAI21X1_171/Y gnd OAI21X1_172/Y vdd OAI21X1
XOAI21X1_183 BUFX4_457/Y BUFX4_134/Y INVX1_473/A gnd OAI21X1_184/C vdd OAI21X1
XOAI21X1_150 NAND2X1_18/Y BUFX4_280/Y OAI21X1_150/C gnd OAI21X1_150/Y vdd OAI21X1
XOAI21X1_161 BUFX4_412/Y BUFX4_173/Y NAND2X1_507/B gnd OAI21X1_161/Y vdd OAI21X1
XINVX1_203 INVX1_203/A gnd INVX1_203/Y vdd INVX1
XOAI21X1_194 BUFX4_395/Y NAND2X1_22/Y OAI21X1_193/Y gnd OAI21X1_194/Y vdd OAI21X1
XINVX1_225 INVX1_225/A gnd INVX1_225/Y vdd INVX1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XINVX1_258 INVX1_258/A gnd INVX1_258/Y vdd INVX1
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XINVX1_236 INVX1_236/A gnd INVX1_236/Y vdd INVX1
XINVX1_269 INVX1_269/A gnd INVX1_269/Y vdd INVX1
XNAND2X1_25 BUFX4_332/Y NOR2X1_11/Y gnd NAND2X1_25/Y vdd NAND2X1
XNAND2X1_14 INVX2_1/Y INVX8_12/A gnd OAI21X1_82/B vdd NAND2X1
XNAND2X1_36 INVX8_7/A NOR2X1_21/Y gnd NAND2X1_36/Y vdd NAND2X1
XNAND2X1_47 BUFX4_350/Y AOI22X1_9/D gnd BUFX4_436/A vdd NAND2X1
XNAND2X1_58 BUFX4_162/Y NOR2X1_51/Y gnd NAND2X1_58/Y vdd NAND2X1
XNAND2X1_69 BUFX4_163/Y NOR2X1_61/Y gnd NAND2X1_69/Y vdd NAND2X1
XAOI21X1_207 AOI21X1_1/A NOR2X1_256/B NOR2X1_256/Y gnd DFFPOSX1_9/D vdd AOI21X1
XFILL_32_1_1 gnd vdd FILL
XAOI21X1_218 BUFX4_301/Y NOR2X1_265/Y NOR2X1_269/Y gnd DFFPOSX1_44/D vdd AOI21X1
XAOI21X1_229 BUFX4_285/Y NOR2X1_279/B NOR2X1_282/Y gnd DFFPOSX1_23/D vdd AOI21X1
XAOI22X1_23 AOI22X1_23/A BUFX4_323/Y AOI22X1_6/C MUX2X1_114/Y gnd AOI22X1_23/Y vdd
+ AOI22X1
XAOI22X1_12 MUX2X1_57/Y BUFX4_350/Y AOI22X1_7/C MUX2X1_60/Y gnd AOI22X1_12/Y vdd AOI22X1
XAOI22X1_56 MUX2X1_267/Y BUFX4_324/Y BUFX4_290/Y AOI22X1_56/D gnd AOI22X1_56/Y vdd
+ AOI22X1
XAOI22X1_45 AOI22X1_45/A AOI22X1_7/B BUFX4_159/Y MUX2X1_216/Y gnd AOI22X1_45/Y vdd
+ AOI22X1
XAOI22X1_34 AOI22X1_34/A AOI22X1_9/A NAND2X1_5/B AOI22X1_34/D gnd AOI22X1_34/Y vdd
+ AOI22X1
XOAI21X1_1413 BUFX4_460/Y BUFX4_388/Y INVX1_133/A gnd OAI21X1_1414/C vdd OAI21X1
XOAI21X1_1402 BUFX4_397/Y NAND2X1_812/Y OAI21X1_1401/Y gnd OAI21X1_1402/Y vdd OAI21X1
XOAI21X1_1457 BUFX4_167/Y INVX2_8/A INVX1_44/A gnd OAI21X1_1457/Y vdd OAI21X1
XAOI22X1_78 MUX2X1_375/Y BUFX4_322/Y BUFX4_290/Y MUX2X1_378/Y gnd AOI22X1_78/Y vdd
+ AOI22X1
XAOI22X1_67 AOI22X1_67/A AOI22X1_7/B BUFX4_159/Y AOI22X1_67/D gnd AOI22X1_67/Y vdd
+ AOI22X1
XOAI21X1_1446 INVX1_326/Y NOR2X1_321/Y NAND2X1_821/Y gnd DFFPOSX1_150/D vdd OAI21X1
XOAI21X1_1435 BUFX4_151/Y BUFX4_390/Y NAND2X1_556/B gnd OAI21X1_1435/Y vdd OAI21X1
XOAI21X1_1424 BUFX4_373/Y NAND2X1_814/Y OAI21X1_1423/Y gnd OAI21X1_1424/Y vdd OAI21X1
XOAI21X1_1479 BUFX4_417/Y BUFX4_392/Y NAND2X1_421/B gnd OAI21X1_1480/C vdd OAI21X1
XOAI21X1_1468 NAND2X1_832/Y BUFX4_99/Y OAI21X1_1468/C gnd OAI21X1_1468/Y vdd OAI21X1
XFILL_23_1_1 gnd vdd FILL
XDFFPOSX1_1009 MUX2X1_26/B CLKBUF1_10/Y AOI21X1_186/Y gnd vdd DFFPOSX1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XBUFX4_320 BUFX4_321/A gnd BUFX4_320/Y vdd BUFX4
XBUFX4_331 d[2] gnd NAND2X1_8/A vdd BUFX4
XBUFX4_342 BUFX4_338/A gnd BUFX4_342/Y vdd BUFX4
XBUFX4_353 BUFX4_354/A gnd INVX1_6/A vdd BUFX4
XBUFX4_364 a[2] gnd BUFX4_364/Y vdd BUFX4
XBUFX4_386 BUFX4_385/A gnd BUFX4_386/Y vdd BUFX4
XBUFX4_375 INVX8_9/Y gnd BUFX4_375/Y vdd BUFX4
XBUFX4_397 INVX8_6/Y gnd BUFX4_397/Y vdd BUFX4
XFILL_26_1 gnd vdd FILL
XOAI21X1_908 INVX1_120/Y BUFX4_202/Y OAI21X1_908/C gnd MUX2X1_86/A vdd OAI21X1
XOAI21X1_919 INVX1_131/Y BUFX4_224/Y NAND2X1_347/Y gnd MUX2X1_95/B vdd OAI21X1
XOAI21X1_1221 INVX1_433/Y BUFX4_234/Y NAND2X1_672/Y gnd MUX2X1_322/B vdd OAI21X1
XOAI21X1_1210 INVX1_422/Y BUFX4_212/Y NAND2X1_660/Y gnd MUX2X1_313/A vdd OAI21X1
XDFFPOSX1_833 MUX2X1_8/B CLKBUF1_7/Y OAI21X1_623/Y gnd vdd DFFPOSX1
XOAI21X1_1265 INVX1_477/Y BUFX4_223/Y NAND2X1_720/Y gnd MUX2X1_355/B vdd OAI21X1
XOAI21X1_1254 INVX1_466/Y BUFX4_201/Y NAND2X1_708/Y gnd MUX2X1_346/A vdd OAI21X1
XOAI21X1_1232 INVX1_444/Y BUFX4_256/Y NAND2X1_683/Y gnd MUX2X1_329/A vdd OAI21X1
XDFFPOSX1_822 INVX1_368/A CLKBUF1_30/Y OAI21X1_619/Y gnd vdd DFFPOSX1
XDFFPOSX1_811 NOR2X1_127/A CLKBUF1_26/Y AOI21X1_101/Y gnd vdd DFFPOSX1
XOAI21X1_1243 INVX1_455/Y BUFX4_278/Y NAND2X1_696/Y gnd MUX2X1_338/B vdd OAI21X1
XDFFPOSX1_800 NOR2X1_121/A CLKBUF1_92/Y AOI21X1_97/Y gnd vdd DFFPOSX1
XDFFPOSX1_844 NAND2X1_465/B CLKBUF1_15/Y OAI21X1_645/Y gnd vdd DFFPOSX1
XDFFPOSX1_855 INVX1_434/A CLKBUF1_19/Y OAI21X1_659/Y gnd vdd DFFPOSX1
XOAI21X1_1276 INVX1_488/Y BUFX4_245/Y NAND2X1_731/Y gnd MUX2X1_362/A vdd OAI21X1
XOAI21X1_1298 INVX1_61/Y NOR2X1_254/Y NAND2X1_757/Y gnd DFFPOSX1_26/D vdd OAI21X1
XDFFPOSX1_866 INVX1_115/A CLKBUF1_13/Y OAI21X1_661/Y gnd vdd DFFPOSX1
XOAI21X1_1287 INVX1_499/Y BUFX4_267/Y NAND2X1_743/Y gnd MUX2X1_371/B vdd OAI21X1
XDFFPOSX1_877 NOR2X1_162/A CLKBUF1_91/Y AOI21X1_130/Y gnd vdd DFFPOSX1
XDFFPOSX1_899 INVX1_181/A CLKBUF1_101/Y OAI21X1_680/Y gnd vdd DFFPOSX1
XDFFPOSX1_888 INVX1_500/A CLKBUF1_54/Y OAI21X1_674/Y gnd vdd DFFPOSX1
XFILL_46_0_1 gnd vdd FILL
XDFFPOSX1_118 INVX1_324/A CLKBUF1_55/Y OAI21X1_1388/Y gnd vdd DFFPOSX1
XDFFPOSX1_107 NOR2X1_314/A CLKBUF1_20/Y AOI21X1_249/Y gnd vdd DFFPOSX1
XCLKBUF1_1 BUFX4_14/Y gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_129 INVX1_41/A CLKBUF1_102/Y OAI21X1_1410/Y gnd vdd DFFPOSX1
XBUFX4_172 BUFX4_168/A gnd BUFX4_172/Y vdd BUFX4
XBUFX4_161 d[0] gnd INVX8_2/A vdd BUFX4
XBUFX4_150 INVX8_11/Y gnd BUFX4_150/Y vdd BUFX4
XFILL_37_0_1 gnd vdd FILL
XNOR2X1_232 NOR2X1_232/A NOR2X1_236/B gnd NOR2X1_232/Y vdd NOR2X1
XNOR2X1_221 NOR2X1_221/A NOR2X1_222/B gnd NOR2X1_221/Y vdd NOR2X1
XBUFX4_183 BUFX4_26/Y gnd MUX2X1_5/S vdd BUFX4
XBUFX4_194 BUFX4_30/Y gnd BUFX4_194/Y vdd BUFX4
XNOR2X1_210 BUFX4_440/Y BUFX4_88/Y gnd NOR2X1_216/B vdd NOR2X1
XNOR2X1_243 INVX1_12/Y INVX1_13/Y gnd AOI22X1_69/C vdd NOR2X1
XNOR2X1_265 NAND3X1_7/Y NOR2X1_265/B gnd NOR2X1_265/Y vdd NOR2X1
XNOR2X1_254 NOR2X1_294/B NAND3X1_7/Y gnd NOR2X1_254/Y vdd NOR2X1
XNOR2X1_276 NOR2X1_276/A NOR2X1_279/B gnd NOR2X1_276/Y vdd NOR2X1
XNOR2X1_298 INVX4_2/Y NOR2X1_265/B gnd INVX8_13/A vdd NOR2X1
XNOR2X1_287 NOR2X1_287/A NOR2X1_289/B gnd NOR2X1_287/Y vdd NOR2X1
XOAI21X1_705 BUFX4_146/Y BUFX4_66/Y NAND2X1_745/B gnd OAI21X1_706/C vdd OAI21X1
XOAI21X1_716 INVX1_247/Y NOR2X1_189/B OAI21X1_716/C gnd OAI21X1_716/Y vdd OAI21X1
XOAI21X1_727 INVX1_504/Y NOR2X1_199/Y OAI21X1_727/C gnd OAI21X1_727/Y vdd OAI21X1
XOAI21X1_749 BUFX4_117/Y OAI21X1_757/B OAI21X1_749/C gnd OAI21X1_749/Y vdd OAI21X1
XOAI21X1_738 BUFX4_455/Y BUFX4_441/Y INVX1_377/A gnd OAI21X1_738/Y vdd OAI21X1
XOAI21X1_1040 INVX1_252/Y BUFX4_268/Y NAND2X1_476/Y gnd MUX2X1_185/A vdd OAI21X1
XMUX2X1_205 MUX2X1_205/A MUX2X1_205/B BUFX4_41/Y gnd MUX2X1_205/Y vdd MUX2X1
XOAI21X1_1073 INVX1_285/Y BUFX4_235/Y NAND2X1_513/Y gnd MUX2X1_211/B vdd OAI21X1
XOAI21X1_1062 INVX1_274/Y BUFX4_213/Y NAND2X1_501/Y gnd MUX2X1_202/A vdd OAI21X1
XDFFPOSX1_630 INVX1_356/A CLKBUF1_6/Y OAI21X1_388/Y gnd vdd DFFPOSX1
XMUX2X1_216 MUX2X1_215/Y MUX2X1_214/Y MUX2X1_84/S gnd MUX2X1_216/Y vdd MUX2X1
XDFFPOSX1_641 INVX1_53/A CLKBUF1_69/Y OAI21X1_409/Y gnd vdd DFFPOSX1
XMUX2X1_238 MUX2X1_238/A MUX2X1_238/B BUFX4_34/Y gnd MUX2X1_240/B vdd MUX2X1
XOAI21X1_1051 INVX1_263/Y BUFX4_191/Y NAND2X1_489/Y gnd MUX2X1_194/B vdd OAI21X1
XMUX2X1_227 MUX2X1_227/A MUX2X1_227/B BUFX4_42/Y gnd MUX2X1_228/A vdd MUX2X1
XOAI21X1_1095 INVX1_307/Y MUX2X1_1/S NAND2X1_536/Y gnd MUX2X1_227/B vdd OAI21X1
XOAI21X1_1084 INVX1_296/Y BUFX4_257/Y NAND2X1_524/Y gnd MUX2X1_218/A vdd OAI21X1
XDFFPOSX1_663 INVX1_422/A CLKBUF1_70/Y OAI21X1_430/Y gnd vdd DFFPOSX1
XDFFPOSX1_674 INVX1_103/A CLKBUF1_96/Y OAI21X1_452/Y gnd vdd DFFPOSX1
XDFFPOSX1_652 NOR2X1_76/A CLKBUF1_88/Y AOI21X1_60/Y gnd vdd DFFPOSX1
XMUX2X1_249 MUX2X1_249/A MUX2X1_249/B MUX2X1_84/S gnd AOI22X1_52/A vdd MUX2X1
XDFFPOSX1_696 INVX1_488/A CLKBUF1_58/Y OAI21X1_496/Y gnd vdd DFFPOSX1
XNAND2X1_700 MUX2X1_11/S NOR2X1_357/A gnd NAND2X1_700/Y vdd NAND2X1
XDFFPOSX1_685 NAND2X1_523/B CLKBUF1_99/Y OAI21X1_474/Y gnd vdd DFFPOSX1
XNAND2X1_711 BUFX4_206/Y NOR2X1_10/A gnd NAND2X1_711/Y vdd NAND2X1
XNAND2X1_755 INVX8_1/Y AOI22X1_1/C gnd NOR2X1_294/B vdd NAND2X1
XNAND2X1_733 BUFX4_248/Y NOR2X1_90/A gnd NAND2X1_733/Y vdd NAND2X1
XNAND2X1_722 BUFX4_226/Y NOR2X1_60/A gnd NAND2X1_722/Y vdd NAND2X1
XNAND2X1_744 BUFX4_268/Y NOR2X1_176/A gnd NAND2X1_744/Y vdd NAND2X1
XNAND2X1_777 BUFX4_335/Y NOR2X1_274/Y gnd NAND2X1_777/Y vdd NAND2X1
XNAND2X1_766 BUFX4_162/Y NOR2X1_264/Y gnd NAND2X1_766/Y vdd NAND2X1
XNAND2X1_788 BUFX4_326/Y NOR2X1_284/Y gnd NAND2X1_788/Y vdd NAND2X1
XNAND2X1_799 BUFX4_327/Y NOR2X1_297/Y gnd NAND2X1_799/Y vdd NAND2X1
XFILL_3_0_1 gnd vdd FILL
XFILL_28_0_1 gnd vdd FILL
XINVX8_3 INVX8_3/A gnd INVX8_3/Y vdd INVX8
XFILL_40_7_0 gnd vdd FILL
XBUFX4_12 clk gnd BUFX4_12/Y vdd BUFX4
XBUFX4_34 BUFX4_75/Y gnd BUFX4_34/Y vdd BUFX4
XBUFX4_23 a[0] gnd BUFX4_23/Y vdd BUFX4
XFILL_48_8_0 gnd vdd FILL
XBUFX4_67 BUFX4_64/A gnd BUFX4_67/Y vdd BUFX4
XBUFX4_78 a[1] gnd BUFX4_78/Y vdd BUFX4
XBUFX4_45 BUFX4_71/Y gnd BUFX4_45/Y vdd BUFX4
XBUFX4_56 BUFX4_57/A gnd BUFX4_56/Y vdd BUFX4
XBUFX4_89 BUFX4_92/A gnd BUFX4_89/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XFILL_31_7_0 gnd vdd FILL
XFILL_39_8_0 gnd vdd FILL
XINVX8_15 INVX8_15/A gnd INVX8_15/Y vdd INVX8
XFILL_22_7_0 gnd vdd FILL
XOAI21X1_513 BUFX4_456/Y BUFX4_293/Y INVX1_57/A gnd OAI21X1_513/Y vdd OAI21X1
XOAI21X1_502 BUFX4_117/Y NAND2X1_97/Y OAI21X1_501/Y gnd OAI21X1_502/Y vdd OAI21X1
XOAI21X1_546 INVX1_106/Y NOR2X1_81/Y NAND2X1_102/Y gnd OAI21X1_546/Y vdd OAI21X1
XOAI21X1_557 INVX1_299/Y NOR2X1_91/Y OAI21X1_557/C gnd OAI21X1_557/Y vdd OAI21X1
XOAI21X1_535 BUFX4_150/Y NOR2X1_91/A NAND2X1_456/B gnd OAI21X1_535/Y vdd OAI21X1
XOAI21X1_524 BUFX4_104/Y NAND2X1_99/Y OAI21X1_524/C gnd OAI21X1_524/Y vdd OAI21X1
XOAI21X1_579 BUFX4_455/Y BUFX4_108/Y INVX1_365/A gnd OAI21X1_580/C vdd OAI21X1
XOAI21X1_568 INVX1_492/Y NOR2X1_101/Y OAI21X1_568/C gnd OAI21X1_568/Y vdd OAI21X1
XDFFPOSX1_471 INVX1_410/A CLKBUF1_23/Y OAI21X1_207/Y gnd vdd DFFPOSX1
XDFFPOSX1_460 OAI21X1_191/C CLKBUF1_5/Y OAI21X1_192/Y gnd vdd DFFPOSX1
XDFFPOSX1_482 INVX1_91/A CLKBUF1_37/Y OAI21X1_210/Y gnd vdd DFFPOSX1
XDFFPOSX1_493 NOR2X1_27/A CLKBUF1_24/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XNAND2X1_530 BUFX4_266/Y OAI21X1_593/C gnd NAND2X1_530/Y vdd NAND2X1
XNAND2X1_563 BUFX4_229/Y NAND2X1_563/B gnd NAND2X1_563/Y vdd NAND2X1
XNAND2X1_541 BUFX4_189/Y NOR2X1_206/A gnd NAND2X1_541/Y vdd NAND2X1
XNAND2X1_552 BUFX4_207/Y NAND2X1_552/B gnd NAND2X1_552/Y vdd NAND2X1
XFILL_5_8_0 gnd vdd FILL
XNAND2X1_596 BUFX4_192/Y NOR2X1_98/A gnd NAND2X1_596/Y vdd NAND2X1
XNAND2X1_574 BUFX4_249/Y OAI21X1_99/C gnd NAND2X1_574/Y vdd NAND2X1
XNAND2X1_585 BUFX4_269/Y NAND2X1_585/B gnd NAND2X1_585/Y vdd NAND2X1
XFILL_13_7_0 gnd vdd FILL
XOAI21X1_321 BUFX4_404/Y BUFX4_381/Y INVX1_290/A gnd OAI21X1_322/C vdd OAI21X1
XOAI21X1_332 BUFX4_419/Y NAND2X1_78/Y OAI21X1_331/Y gnd OAI21X1_332/Y vdd OAI21X1
XOAI21X1_310 INVX1_353/Y NOR2X1_61/Y NAND2X1_74/Y gnd OAI21X1_310/Y vdd OAI21X1
XOAI21X1_354 BUFX4_398/Y NAND2X1_79/Y OAI21X1_354/C gnd OAI21X1_354/Y vdd OAI21X1
XOAI21X1_365 BUFX4_367/Y BUFX4_387/Y NAND2X1_381/B gnd OAI21X1_366/C vdd OAI21X1
XOAI21X1_343 BUFX4_87/Y BUFX4_385/Y NAND2X1_725/B gnd OAI21X1_344/C vdd OAI21X1
XOAI21X1_398 BUFX4_113/Y NAND2X1_82/Y OAI21X1_398/C gnd OAI21X1_398/Y vdd OAI21X1
XOAI21X1_376 BUFX4_380/Y NAND2X1_80/Y OAI21X1_375/Y gnd OAI21X1_376/Y vdd OAI21X1
XOAI21X1_387 BUFX4_172/Y BUFX4_385/Y INVX1_356/A gnd OAI21X1_388/C vdd OAI21X1
XINVX1_407 INVX1_407/A gnd INVX1_407/Y vdd INVX1
XINVX1_418 INVX1_418/A gnd INVX1_418/Y vdd INVX1
XINVX1_429 INVX1_429/A gnd INVX1_429/Y vdd INVX1
XDFFPOSX1_290 INVX1_79/A CLKBUF1_68/Y OAI21X1_1627/Y gnd vdd DFFPOSX1
XNAND2X1_371 BUFX4_269/Y NOR2X1_15/A gnd NAND2X1_371/Y vdd NAND2X1
XNAND2X1_360 BUFX4_247/Y NOR2X1_372/A gnd NAND2X1_360/Y vdd NAND2X1
XNAND2X1_382 BUFX4_190/Y OAI21X1_397/C gnd OAI21X1_952/C vdd NAND2X1
XNAND2X1_393 BUFX4_210/Y NOR2X1_116/A gnd OAI21X1_962/C vdd NAND2X1
XFILL_45_6_0 gnd vdd FILL
XOAI21X1_1639 NAND2X1_860/Y BUFX4_114/Y OAI21X1_1638/Y gnd DFFPOSX1_307/D vdd OAI21X1
XOAI21X1_1606 BUFX4_151/Y BUFX4_345/Y NAND2X1_358/B gnd OAI21X1_1606/Y vdd OAI21X1
XOAI21X1_1617 BUFX4_379/Y NAND2X1_843/Y OAI21X1_1617/C gnd OAI21X1_1617/Y vdd OAI21X1
XOAI21X1_1628 INVX1_143/Y NOR2X1_368/Y NAND2X1_854/Y gnd DFFPOSX1_291/D vdd OAI21X1
XFILL_36_6_0 gnd vdd FILL
XFILL_2_6_0 gnd vdd FILL
XFILL_27_6_0 gnd vdd FILL
XFILL_10_5_0 gnd vdd FILL
XAOI22X1_5 AOI22X1_5/A AOI22X1_1/B AOI22X1_1/C AOI22X1_5/D gnd AOI22X1_5/Y vdd AOI22X1
XOAI21X1_140 NAND2X1_18/Y BUFX4_422/Y OAI21X1_139/Y gnd OAI21X1_140/Y vdd OAI21X1
XOAI21X1_173 BUFX4_457/Y INVX1_1/A INVX1_153/A gnd OAI21X1_174/C vdd OAI21X1
XOAI21X1_151 BUFX4_166/Y BUFX4_175/Y INVX1_472/A gnd OAI21X1_152/C vdd OAI21X1
XOAI21X1_162 BUFX4_394/Y NAND2X1_19/Y OAI21X1_161/Y gnd OAI21X1_162/Y vdd OAI21X1
XINVX1_226 INVX1_226/A gnd INVX1_226/Y vdd INVX1
XINVX1_204 INVX1_204/A gnd INVX1_204/Y vdd INVX1
XOAI21X1_195 BUFX4_147/Y INVX1_1/A OAI21X1_195/C gnd OAI21X1_196/C vdd OAI21X1
XOAI21X1_184 BUFX4_376/Y NAND2X1_21/Y OAI21X1_184/C gnd OAI21X1_184/Y vdd OAI21X1
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XINVX1_248 INVX1_248/A gnd INVX1_248/Y vdd INVX1
XINVX1_237 INVX1_237/A gnd INVX1_237/Y vdd INVX1
XINVX1_259 INVX1_259/A gnd INVX1_259/Y vdd INVX1
XNAND2X1_15 INVX2_1/Y INVX8_13/A gnd OAI21X1_96/B vdd NAND2X1
XNAND2X1_48 INVX8_10/A INVX2_2/Y gnd NAND2X1_48/Y vdd NAND2X1
XNAND2X1_59 BUFX4_449/Y NOR2X1_51/Y gnd NAND2X1_59/Y vdd NAND2X1
XNAND2X1_26 BUFX4_142/Y NOR2X1_11/Y gnd NAND2X1_26/Y vdd NAND2X1
XNAND2X1_37 INVX8_8/A NOR2X1_21/Y gnd NAND2X1_37/Y vdd NAND2X1
XNAND2X1_190 BUFX4_453/Y NOR2X1_199/Y gnd OAI21X1_721/C vdd NAND2X1
XFILL_18_6_0 gnd vdd FILL
XAOI21X1_219 BUFX4_402/Y NOR2X1_265/Y NOR2X1_270/Y gnd AOI21X1_219/Y vdd AOI21X1
XAOI21X1_208 BUFX4_426/Y NOR2X1_256/B NOR2X1_257/Y gnd AOI21X1_208/Y vdd AOI21X1
XAOI22X1_24 AOI22X1_24/A AOI22X1_9/A NAND2X1_5/B AOI22X1_24/D gnd AOI22X1_24/Y vdd
+ AOI22X1
XAOI22X1_13 MUX2X1_63/Y BUFX4_323/Y AOI22X1_6/C MUX2X1_66/Y gnd AOI22X1_13/Y vdd AOI22X1
XAOI22X1_35 AOI22X1_35/A BUFX4_352/Y BUFX4_157/Y MUX2X1_168/Y gnd AOI22X1_35/Y vdd
+ AOI22X1
XAOI22X1_46 AOI22X1_46/A BUFX4_322/Y BUFX4_292/Y AOI22X1_46/D gnd AOI22X1_46/Y vdd
+ AOI22X1
XAOI22X1_57 AOI22X1_57/A INVX1_6/A INVX1_8/A AOI22X1_57/D gnd AOI22X1_57/Y vdd AOI22X1
XOAI21X1_1403 BUFX4_416/Y BUFX4_466/Y NAND2X1_555/B gnd OAI21X1_1403/Y vdd OAI21X1
XOAI21X1_1414 BUFX4_112/Y NAND2X1_814/Y OAI21X1_1414/C gnd DFFPOSX1_131/D vdd OAI21X1
XAOI22X1_79 AOI22X1_79/A AOI22X1_9/D AOI22X1_69/C AOI22X1_79/D gnd AOI22X1_79/Y vdd
+ AOI22X1
XAOI22X1_68 MUX2X1_327/Y BUFX4_322/Y BUFX4_292/Y MUX2X1_330/Y gnd AOI22X1_68/Y vdd
+ AOI22X1
XOAI21X1_1436 BUFX4_99/Y NAND2X1_815/Y OAI21X1_1435/Y gnd OAI21X1_1436/Y vdd OAI21X1
XOAI21X1_1425 BUFX4_151/Y BUFX4_390/Y NAND2X1_247/B gnd OAI21X1_1425/Y vdd OAI21X1
XOAI21X1_1447 INVX1_390/Y NOR2X1_321/Y NAND2X1_822/Y gnd DFFPOSX1_151/D vdd OAI21X1
XOAI21X1_1469 BUFX4_167/Y BUFX4_392/Y INVX1_392/A gnd OAI21X1_1469/Y vdd OAI21X1
XOAI21X1_1458 NAND2X1_832/Y BUFX4_125/Y OAI21X1_1457/Y gnd DFFPOSX1_177/D vdd OAI21X1
XFILL_42_4_0 gnd vdd FILL
XAOI21X1_90 BUFX4_130/Y NOR2X1_118/B NOR2X1_114/Y gnd AOI21X1_90/Y vdd AOI21X1
XBUFX4_310 INVX8_14/Y gnd BUFX4_310/Y vdd BUFX4
XBUFX4_321 BUFX4_321/A gnd BUFX4_321/Y vdd BUFX4
XBUFX4_354 BUFX4_354/A gnd BUFX4_354/Y vdd BUFX4
XBUFX4_332 d[2] gnd BUFX4_332/Y vdd BUFX4
XBUFX4_343 BUFX4_344/A gnd BUFX4_343/Y vdd BUFX4
XBUFX4_387 BUFX4_385/A gnd BUFX4_387/Y vdd BUFX4
XBUFX4_398 INVX8_6/Y gnd BUFX4_398/Y vdd BUFX4
XBUFX4_376 INVX8_9/Y gnd BUFX4_376/Y vdd BUFX4
XBUFX4_365 a[2] gnd MUX2X1_96/S vdd BUFX4
XFILL_26_2 gnd vdd FILL
XFILL_33_4_0 gnd vdd FILL
XFILL_19_1 gnd vdd FILL
XOAI21X1_909 INVX1_121/Y BUFX4_204/Y NAND2X1_335/Y gnd MUX2X1_88/B vdd OAI21X1
XOAI21X1_1222 INVX1_434/Y BUFX4_236/Y NAND2X1_673/Y gnd MUX2X1_322/A vdd OAI21X1
XOAI21X1_1211 INVX1_423/Y BUFX4_214/Y NAND2X1_661/Y gnd MUX2X1_314/B vdd OAI21X1
XOAI21X1_1200 INVX1_412/Y BUFX4_192/Y NAND2X1_649/Y gnd MUX2X1_305/A vdd OAI21X1
XOAI21X1_1244 INVX1_456/Y MUX2X1_2/S NAND2X1_697/Y gnd MUX2X1_338/A vdd OAI21X1
XOAI21X1_1255 INVX1_467/Y BUFX4_203/Y NAND2X1_709/Y gnd MUX2X1_347/B vdd OAI21X1
XOAI21X1_1233 INVX1_445/Y BUFX4_258/Y NAND2X1_686/Y gnd MUX2X1_331/B vdd OAI21X1
XDFFPOSX1_823 INVX1_432/A CLKBUF1_44/Y OAI21X1_620/Y gnd vdd DFFPOSX1
XDFFPOSX1_801 MUX2X1_4/B CLKBUF1_88/Y AOI21X1_98/Y gnd vdd DFFPOSX1
XDFFPOSX1_812 NOR2X1_128/A CLKBUF1_61/Y AOI21X1_102/Y gnd vdd DFFPOSX1
XDFFPOSX1_845 NAND2X1_534/B CLKBUF1_15/Y OAI21X1_647/Y gnd vdd DFFPOSX1
XDFFPOSX1_834 INVX1_113/A CLKBUF1_81/Y OAI21X1_625/Y gnd vdd DFFPOSX1
XOAI21X1_1266 INVX1_478/Y BUFX4_225/Y NAND2X1_721/Y gnd MUX2X1_355/A vdd OAI21X1
XDFFPOSX1_856 INVX1_498/A CLKBUF1_13/Y OAI21X1_660/Y gnd vdd DFFPOSX1
XOAI21X1_1288 INVX1_500/Y BUFX4_269/Y NAND2X1_744/Y gnd MUX2X1_371/A vdd OAI21X1
XOAI21X1_1277 INVX1_489/Y BUFX4_247/Y NAND2X1_732/Y gnd MUX2X1_364/B vdd OAI21X1
XDFFPOSX1_867 INVX1_179/A CLKBUF1_19/Y OAI21X1_662/Y gnd vdd DFFPOSX1
XDFFPOSX1_878 NOR2X1_163/A CLKBUF1_81/Y AOI21X1_131/Y gnd vdd DFFPOSX1
XDFFPOSX1_889 MUX2X1_12/A CLKBUF1_1/Y AOI21X1_135/Y gnd vdd DFFPOSX1
XOAI21X1_1299 INVX1_125/Y NOR2X1_254/Y NAND2X1_758/Y gnd DFFPOSX1_27/D vdd OAI21X1
XFILL_24_4_0 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XFILL_15_4_0 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_1/S gnd MUX2X1_3/B vdd MUX2X1
XDFFPOSX1_119 INVX1_388/A CLKBUF1_42/Y OAI21X1_1390/Y gnd vdd DFFPOSX1
XDFFPOSX1_108 NOR2X1_315/A CLKBUF1_53/Y AOI21X1_250/Y gnd vdd DFFPOSX1
XCLKBUF1_2 BUFX4_11/Y gnd CLKBUF1_2/Y vdd CLKBUF1
XNOR2X1_200 MUX2X1_19/B NOR2X1_199/Y gnd NOR2X1_200/Y vdd NOR2X1
XBUFX4_140 d[6] gnd BUFX4_140/Y vdd BUFX4
XBUFX4_162 d[0] gnd BUFX4_162/Y vdd BUFX4
XBUFX4_173 BUFX4_178/A gnd BUFX4_173/Y vdd BUFX4
XBUFX4_151 INVX8_11/Y gnd BUFX4_151/Y vdd BUFX4
XNOR2X1_233 NOR2X1_233/A NOR2X1_236/B gnd NOR2X1_233/Y vdd NOR2X1
XBUFX4_184 BUFX4_26/Y gnd MUX2X1_8/S vdd BUFX4
XNOR2X1_222 NOR2X1_222/A NOR2X1_222/B gnd NOR2X1_222/Y vdd NOR2X1
XBUFX4_195 BUFX4_31/Y gnd BUFX4_195/Y vdd BUFX4
XNOR2X1_211 MUX2X1_23/A NOR2X1_216/B gnd NOR2X1_211/Y vdd NOR2X1
XNOR2X1_266 NOR2X1_266/A NOR2X1_265/Y gnd NOR2X1_266/Y vdd NOR2X1
XNOR2X1_255 NOR2X1_255/A NAND3X1_7/Y gnd NOR2X1_256/B vdd NOR2X1
XNOR2X1_244 BUFX4_52/Y INVX2_6/Y gnd NOR2X1_244/Y vdd NOR2X1
XNOR2X1_277 NOR2X1_277/A NOR2X1_279/B gnd NOR2X1_277/Y vdd NOR2X1
XNOR2X1_288 NOR2X1_288/A NOR2X1_289/B gnd NOR2X1_288/Y vdd NOR2X1
XNOR2X1_299 BUFX4_463/Y BUFX4_84/Y gnd NOR2X1_303/B vdd NOR2X1
XOAI21X1_706 BUFX4_375/Y OAI21X1_704/B OAI21X1_706/C gnd OAI21X1_706/Y vdd OAI21X1
XOAI21X1_717 INVX1_311/Y NOR2X1_189/B OAI21X1_717/C gnd OAI21X1_717/Y vdd OAI21X1
XOAI21X1_739 BUFX4_103/Y OAI21X1_729/B OAI21X1_738/Y gnd OAI21X1_739/Y vdd OAI21X1
XOAI21X1_728 BUFX4_455/Y INVX2_5/A MUX2X1_22/B gnd OAI21X1_728/Y vdd OAI21X1
XOAI21X1_1030 INVX1_242/Y BUFX4_248/Y NAND2X1_466/Y gnd MUX2X1_178/A vdd OAI21X1
XDFFPOSX1_631 INVX1_420/A CLKBUF1_79/Y OAI21X1_390/Y gnd vdd DFFPOSX1
XOAI21X1_1063 INVX1_275/Y BUFX4_215/Y NAND2X1_502/Y gnd MUX2X1_203/B vdd OAI21X1
XDFFPOSX1_620 NAND2X1_450/B CLKBUF1_28/Y OAI21X1_368/Y gnd vdd DFFPOSX1
XOAI21X1_1041 INVX1_253/Y BUFX4_270/Y NAND2X1_479/Y gnd MUX2X1_187/B vdd OAI21X1
XMUX2X1_217 MUX2X1_217/A MUX2X1_217/B BUFX4_53/Y gnd MUX2X1_217/Y vdd MUX2X1
XMUX2X1_206 MUX2X1_206/A MUX2X1_206/B BUFX4_57/Y gnd MUX2X1_207/A vdd MUX2X1
XOAI21X1_1052 INVX1_264/Y BUFX4_193/Y NAND2X1_490/Y gnd MUX2X1_194/A vdd OAI21X1
XMUX2X1_228 MUX2X1_228/A MUX2X1_228/B MUX2X1_96/S gnd AOI22X1_47/D vdd MUX2X1
XDFFPOSX1_664 INVX1_486/A CLKBUF1_96/Y OAI21X1_432/Y gnd vdd DFFPOSX1
XDFFPOSX1_675 INVX1_167/A CLKBUF1_45/Y OAI21X1_454/Y gnd vdd DFFPOSX1
XDFFPOSX1_642 INVX1_101/A CLKBUF1_88/Y OAI21X1_410/Y gnd vdd DFFPOSX1
XDFFPOSX1_653 NOR2X1_77/A CLKBUF1_88/Y AOI21X1_61/Y gnd vdd DFFPOSX1
XMUX2X1_239 MUX2X1_239/A MUX2X1_239/B BUFX4_54/Y gnd MUX2X1_240/A vdd MUX2X1
XOAI21X1_1085 INVX1_297/Y BUFX4_259/Y NAND2X1_525/Y gnd MUX2X1_220/B vdd OAI21X1
XOAI21X1_1074 INVX1_286/Y BUFX4_237/Y NAND2X1_514/Y gnd MUX2X1_211/A vdd OAI21X1
XOAI21X1_1096 INVX1_308/Y MUX2X1_4/S NAND2X1_537/Y gnd MUX2X1_227/A vdd OAI21X1
XNAND2X1_701 BUFX4_188/Y NAND2X1_701/B gnd NAND2X1_701/Y vdd NAND2X1
XDFFPOSX1_697 OAI21X1_497/C CLKBUF1_99/Y OAI21X1_498/Y gnd vdd DFFPOSX1
XDFFPOSX1_686 NAND2X1_592/B CLKBUF1_99/Y OAI21X1_476/Y gnd vdd DFFPOSX1
XNAND2X1_712 BUFX4_208/Y NAND2X1_712/B gnd NAND2X1_712/Y vdd NAND2X1
XNAND2X1_745 BUFX4_270/Y NAND2X1_745/B gnd NAND2X1_745/Y vdd NAND2X1
XNAND2X1_734 BUFX4_250/Y NOR2X1_100/A gnd NAND2X1_734/Y vdd NAND2X1
XNAND2X1_723 BUFX4_228/Y OAI21X1_303/C gnd NAND2X1_723/Y vdd NAND2X1
XNAND2X1_767 BUFX4_452/Y NOR2X1_264/Y gnd NAND2X1_767/Y vdd NAND2X1
XNAND2X1_756 BUFX4_164/Y NOR2X1_254/Y gnd NAND2X1_756/Y vdd NAND2X1
XNAND2X1_778 BUFX4_145/Y NOR2X1_274/Y gnd NAND2X1_778/Y vdd NAND2X1
XNAND2X1_789 BUFX4_136/Y NOR2X1_284/Y gnd NAND2X1_789/Y vdd NAND2X1
XFILL_40_7_1 gnd vdd FILL
XINVX8_4 INVX8_4/A gnd INVX8_4/Y vdd INVX8
XDFFPOSX1_90 NOR2X1_301/A CLKBUF1_68/Y DFFPOSX1_90/D gnd vdd DFFPOSX1
XBUFX4_24 a[0] gnd BUFX4_24/Y vdd BUFX4
XBUFX4_35 BUFX4_75/Y gnd BUFX4_35/Y vdd BUFX4
XBUFX4_13 clk gnd BUFX4_13/Y vdd BUFX4
XFILL_48_8_1 gnd vdd FILL
XBUFX4_68 a[1] gnd BUFX4_41/A vdd BUFX4
XBUFX4_46 BUFX4_71/Y gnd BUFX4_46/Y vdd BUFX4
XBUFX4_57 BUFX4_57/A gnd BUFX4_57/Y vdd BUFX4
XFILL_47_3_0 gnd vdd FILL
XBUFX4_79 a[1] gnd INVX4_1/A vdd BUFX4
XFILL_31_7_1 gnd vdd FILL
XFILL_30_2_0 gnd vdd FILL
XFILL_39_8_1 gnd vdd FILL
XFILL_38_3_0 gnd vdd FILL
XINVX8_16 INVX8_16/A gnd INVX8_16/Y vdd INVX8
XFILL_22_7_1 gnd vdd FILL
XOAI21X1_514 BUFX4_126/Y NAND2X1_99/Y OAI21X1_513/Y gnd OAI21X1_514/Y vdd OAI21X1
XOAI21X1_503 BUFX4_414/Y BUFX4_342/Y NAND2X1_455/B gnd OAI21X1_504/C vdd OAI21X1
XFILL_21_2_0 gnd vdd FILL
XOAI21X1_547 INVX1_170/Y NOR2X1_81/Y OAI21X1_547/C gnd OAI21X1_547/Y vdd OAI21X1
XOAI21X1_536 BUFX4_298/Y OAI21X1_544/B OAI21X1_535/Y gnd OAI21X1_536/Y vdd OAI21X1
XOAI21X1_525 NOR2X1_1/B BUFX4_293/Y INVX1_425/A gnd OAI21X1_525/Y vdd OAI21X1
XOAI21X1_569 NOR2X1_1/B BUFX4_108/Y MUX2X1_1/B gnd OAI21X1_570/C vdd OAI21X1
XOAI21X1_558 INVX1_363/Y NOR2X1_91/Y OAI21X1_558/C gnd OAI21X1_558/Y vdd OAI21X1
XDFFPOSX1_461 NAND2X1_508/B CLKBUF1_87/Y OAI21X1_194/Y gnd vdd DFFPOSX1
XDFFPOSX1_450 INVX1_89/A CLKBUF1_18/Y OAI21X1_172/Y gnd vdd DFFPOSX1
XDFFPOSX1_472 INVX1_474/A CLKBUF1_40/Y OAI21X1_208/Y gnd vdd DFFPOSX1
XDFFPOSX1_483 INVX1_155/A CLKBUF1_93/Y OAI21X1_211/Y gnd vdd DFFPOSX1
XNAND2X1_520 BUFX4_248/Y NAND2X1_520/B gnd NAND2X1_520/Y vdd NAND2X1
XDFFPOSX1_494 NOR2X1_28/A CLKBUF1_31/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XNAND2X1_542 BUFX4_191/Y NAND2X1_542/B gnd NAND2X1_542/Y vdd NAND2X1
XNAND2X1_531 BUFX4_268/Y NOR2X1_118/A gnd NAND2X1_531/Y vdd NAND2X1
XNAND2X1_553 BUFX4_209/Y NOR2X1_305/A gnd NAND2X1_553/Y vdd NAND2X1
XFILL_5_8_1 gnd vdd FILL
XNAND2X1_586 BUFX4_271/Y NOR2X1_68/A gnd NAND2X1_586/Y vdd NAND2X1
XNAND2X1_564 AOI22X1_50/Y AOI22X1_51/Y gnd AOI22X1_54/A vdd NAND2X1
XNAND2X1_597 BUFX4_194/Y NOR2X1_108/A gnd NAND2X1_597/Y vdd NAND2X1
XNAND2X1_575 BUFX4_251/Y OAI21X1_131/C gnd NAND2X1_575/Y vdd NAND2X1
XFILL_4_3_0 gnd vdd FILL
XFILL_29_3_0 gnd vdd FILL
XFILL_13_7_1 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XOAI21X1_322 BUFX4_401/Y NAND2X1_77/Y OAI21X1_322/C gnd OAI21X1_322/Y vdd OAI21X1
XOAI21X1_311 INVX1_417/Y NOR2X1_61/Y NAND2X1_75/Y gnd OAI21X1_311/Y vdd OAI21X1
XOAI21X1_300 AOI21X1_6/A NAND2X1_67/Y OAI21X1_299/Y gnd OAI21X1_300/Y vdd OAI21X1
XOAI21X1_333 BUFX4_85/Y INVX2_3/A OAI21X1_333/C gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_355 BUFX4_307/Y BUFX4_387/Y INVX1_355/A gnd OAI21X1_355/Y vdd OAI21X1
XOAI21X1_344 BUFX4_378/Y NAND2X1_78/Y OAI21X1_344/C gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_377 BUFX4_172/Y BUFX4_384/Y INVX1_52/A gnd OAI21X1_377/Y vdd OAI21X1
XOAI21X1_399 BUFX4_415/Y BUFX4_386/Y NAND2X1_451/B gnd OAI21X1_399/Y vdd OAI21X1
XOAI21X1_366 BUFX4_109/Y NAND2X1_80/Y OAI21X1_366/C gnd OAI21X1_366/Y vdd OAI21X1
XOAI21X1_388 NAND2X1_81/Y BUFX4_102/Y OAI21X1_388/C gnd OAI21X1_388/Y vdd OAI21X1
XINVX1_408 INVX1_408/A gnd INVX1_408/Y vdd INVX1
XINVX1_419 INVX1_419/A gnd INVX1_419/Y vdd INVX1
XDFFPOSX1_280 INVX1_462/A CLKBUF1_77/Y DFFPOSX1_280/D gnd vdd DFFPOSX1
XDFFPOSX1_291 INVX1_143/A CLKBUF1_53/Y DFFPOSX1_291/D gnd vdd DFFPOSX1
XNAND2X1_361 BUFX4_249/Y NAND2X1_361/B gnd NAND2X1_361/Y vdd NAND2X1
XNAND2X1_372 BUFX4_271/Y NOR2X1_25/A gnd OAI21X1_943/C vdd NAND2X1
XNAND2X1_350 BUFX4_229/Y NOR2X1_325/A gnd OAI21X1_922/C vdd NAND2X1
XNAND2X1_383 BUFX4_192/Y NOR2X1_75/A gnd NAND2X1_383/Y vdd NAND2X1
XNAND2X1_394 BUFX4_212/Y NOR2X1_127/A gnd OAI21X1_963/C vdd NAND2X1
XFILL_45_6_1 gnd vdd FILL
XFILL_44_1_0 gnd vdd FILL
XOAI21X1_1618 INVX1_19/Y NOR2X1_358/Y NAND2X1_844/Y gnd OAI21X1_1618/Y vdd OAI21X1
XOAI21X1_1607 AOI21X1_3/A NAND2X1_843/Y OAI21X1_1606/Y gnd OAI21X1_1607/Y vdd OAI21X1
XOAI21X1_1629 INVX1_207/Y NOR2X1_368/Y NAND2X1_855/Y gnd OAI21X1_1629/Y vdd OAI21X1
XFILL_7_1 gnd vdd FILL
XFILL_49_1 gnd vdd FILL
XFILL_36_6_1 gnd vdd FILL
XFILL_35_1_0 gnd vdd FILL
XNAND3X1_1 NAND3X1_1/A NAND3X1_1/B NAND3X1_1/C gnd AOI22X1_3/A vdd NAND3X1
XFILL_2_6_1 gnd vdd FILL
XFILL_27_6_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XFILL_10_5_1 gnd vdd FILL
XOAI21X1_130 BUFX4_399/Y NAND2X1_17/Y OAI21X1_130/C gnd OAI21X1_130/Y vdd OAI21X1
XOAI21X1_174 AOI21X1_3/A NAND2X1_21/Y OAI21X1_174/C gnd OAI21X1_174/Y vdd OAI21X1
XAOI22X1_6 AOI22X1_6/A INVX1_10/A AOI22X1_6/C AOI22X1_6/D gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_152 NAND2X1_18/Y BUFX4_374/Y OAI21X1_152/C gnd OAI21X1_152/Y vdd OAI21X1
XOAI21X1_163 BUFX4_411/Y BUFX4_178/Y OAI21X1_163/C gnd OAI21X1_163/Y vdd OAI21X1
XOAI21X1_141 INVX4_3/A BUFX4_173/Y INVX1_152/A gnd OAI21X1_141/Y vdd OAI21X1
XOAI21X1_185 BUFX4_147/Y INVX1_1/A NAND2X1_229/B gnd OAI21X1_186/C vdd OAI21X1
XOAI21X1_196 BUFX4_98/Y NAND2X1_22/Y OAI21X1_196/C gnd OAI21X1_196/Y vdd OAI21X1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XINVX1_227 INVX1_227/A gnd INVX1_227/Y vdd INVX1
XINVX1_249 INVX1_249/A gnd INVX1_249/Y vdd INVX1
XINVX1_238 INVX1_238/A gnd INVX1_238/Y vdd INVX1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_16 INVX2_1/Y INVX8_14/A gnd NAND2X1_16/Y vdd NAND2X1
XNAND2X1_180 INVX8_7/A NOR2X1_177/Y gnd OAI21X1_711/C vdd NAND2X1
XNAND2X1_27 BUFX4_445/Y NOR2X1_11/Y gnd NAND2X1_27/Y vdd NAND2X1
XNAND2X1_38 INVX8_9/A NOR2X1_21/Y gnd NAND2X1_38/Y vdd NAND2X1
XNAND2X1_49 INVX8_11/A INVX2_2/Y gnd NAND2X1_49/Y vdd NAND2X1
XNAND2X1_191 BUFX4_335/Y NOR2X1_199/Y gnd OAI21X1_722/C vdd NAND2X1
XFILL_18_6_1 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XAOI21X1_209 BUFX4_113/Y NOR2X1_256/B NOR2X1_258/Y gnd AOI21X1_209/Y vdd AOI21X1
XAOI22X1_14 AOI22X1_14/A AOI22X1_9/A NAND2X1_5/B AOI22X1_14/D gnd AOI22X1_14/Y vdd
+ AOI22X1
XAOI22X1_36 MUX2X1_171/Y BUFX4_324/Y BUFX4_290/Y AOI22X1_36/D gnd AOI22X1_36/Y vdd
+ AOI22X1
XAOI22X1_25 AOI22X1_25/A BUFX4_350/Y AOI22X1_7/C MUX2X1_120/Y gnd AOI22X1_25/Y vdd
+ AOI22X1
XAOI22X1_47 AOI22X1_47/A BUFX4_350/Y AOI22X1_7/C AOI22X1_47/D gnd AOI22X1_47/Y vdd
+ AOI22X1
XOAI21X1_1404 BUFX4_99/Y NAND2X1_812/Y OAI21X1_1403/Y gnd OAI21X1_1404/Y vdd OAI21X1
XAOI22X1_58 MUX2X1_279/Y BUFX4_324/Y BUFX4_290/Y AOI22X1_58/D gnd AOI22X1_58/Y vdd
+ AOI22X1
XAOI22X1_69 AOI22X1_69/A AOI22X1_9/D AOI22X1_69/C AOI22X1_69/D gnd AOI22X1_69/Y vdd
+ AOI22X1
XOAI21X1_1415 BUFX4_457/Y BUFX4_390/Y INVX1_197/A gnd OAI21X1_1416/C vdd OAI21X1
XOAI21X1_1426 BUFX4_125/Y NAND2X1_815/Y OAI21X1_1425/Y gnd OAI21X1_1426/Y vdd OAI21X1
XOAI21X1_1437 BUFX4_151/Y BUFX4_388/Y NAND2X1_625/B gnd OAI21X1_1437/Y vdd OAI21X1
XOAI21X1_1459 BUFX4_167/Y BUFX4_393/Y INVX1_72/A gnd OAI21X1_1459/Y vdd OAI21X1
XOAI21X1_1448 INVX1_454/Y NOR2X1_321/Y NAND2X1_823/Y gnd OAI21X1_1448/Y vdd OAI21X1
XFILL_42_4_1 gnd vdd FILL
XAOI21X1_80 BUFX4_372/Y NOR2X1_96/B AOI21X1_80/C gnd AOI21X1_80/Y vdd AOI21X1
XAOI21X1_91 BUFX4_425/Y NOR2X1_118/B NOR2X1_115/Y gnd AOI21X1_91/Y vdd AOI21X1
XBUFX4_300 INVX8_5/Y gnd BUFX4_300/Y vdd BUFX4
XBUFX4_322 BUFX4_321/A gnd BUFX4_322/Y vdd BUFX4
XBUFX4_311 INVX8_14/Y gnd NOR2X1_91/B vdd BUFX4
XBUFX4_333 d[2] gnd INVX8_4/A vdd BUFX4
XBUFX4_355 a[2] gnd MUX2X1_7/S vdd BUFX4
XBUFX4_344 BUFX4_344/A gnd BUFX4_344/Y vdd BUFX4
XBUFX4_377 INVX8_9/Y gnd BUFX4_377/Y vdd BUFX4
XBUFX4_366 INVX8_15/Y gnd NOR2X1_22/B vdd BUFX4
XBUFX4_388 BUFX4_392/A gnd BUFX4_388/Y vdd BUFX4
XBUFX4_399 INVX8_6/Y gnd BUFX4_399/Y vdd BUFX4
XFILL_33_4_1 gnd vdd FILL
XOAI21X1_1212 INVX1_424/Y BUFX4_216/Y NAND2X1_662/Y gnd MUX2X1_314/A vdd OAI21X1
XOAI21X1_1201 INVX1_413/Y BUFX4_194/Y NAND2X1_651/Y gnd MUX2X1_307/B vdd OAI21X1
XOAI21X1_1234 INVX1_446/Y BUFX4_260/Y NAND2X1_687/Y gnd MUX2X1_331/A vdd OAI21X1
XOAI21X1_1245 INVX1_457/Y MUX2X1_5/S NAND2X1_698/Y gnd MUX2X1_340/B vdd OAI21X1
XOAI21X1_1256 INVX1_468/Y BUFX4_205/Y NAND2X1_710/Y gnd MUX2X1_347/A vdd OAI21X1
XDFFPOSX1_824 INVX1_496/A CLKBUF1_69/Y OAI21X1_621/Y gnd vdd DFFPOSX1
XDFFPOSX1_813 NOR2X1_129/A CLKBUF1_2/Y AOI21X1_103/Y gnd vdd DFFPOSX1
XDFFPOSX1_802 INVX1_111/A CLKBUF1_100/Y OAI21X1_608/Y gnd vdd DFFPOSX1
XOAI21X1_1223 INVX1_435/Y BUFX4_238/Y NAND2X1_674/Y gnd MUX2X1_323/B vdd OAI21X1
XDFFPOSX1_857 MUX2X1_9/A CLKBUF1_15/Y AOI21X1_117/Y gnd vdd DFFPOSX1
XDFFPOSX1_835 INVX1_177/A CLKBUF1_7/Y OAI21X1_627/Y gnd vdd DFFPOSX1
XDFFPOSX1_846 NAND2X1_603/B CLKBUF1_7/Y OAI21X1_649/Y gnd vdd DFFPOSX1
XOAI21X1_1289 INVX1_501/Y BUFX4_271/Y NAND2X1_745/Y gnd MUX2X1_373/B vdd OAI21X1
XOAI21X1_1278 INVX1_490/Y BUFX4_249/Y NAND2X1_733/Y gnd MUX2X1_364/A vdd OAI21X1
XOAI21X1_1267 INVX1_479/Y BUFX4_227/Y NAND2X1_722/Y gnd MUX2X1_356/B vdd OAI21X1
XDFFPOSX1_879 NOR2X1_164/A CLKBUF1_80/Y AOI21X1_132/Y gnd vdd DFFPOSX1
XDFFPOSX1_868 INVX1_243/A CLKBUF1_81/Y OAI21X1_663/Y gnd vdd DFFPOSX1
XFILL_24_4_1 gnd vdd FILL
XFILL_7_5_1 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XFILL_15_4_1 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_2/S gnd MUX2X1_3/A vdd MUX2X1
XDFFPOSX1_109 NOR2X1_316/A CLKBUF1_39/Y AOI21X1_251/Y gnd vdd DFFPOSX1
XCLKBUF1_3 BUFX4_13/Y gnd CLKBUF1_3/Y vdd CLKBUF1
XBUFX4_130 INVX8_2/Y gnd BUFX4_130/Y vdd BUFX4
XBUFX4_141 d[3] gnd NAND2X1_9/A vdd BUFX4
XBUFX4_163 d[0] gnd BUFX4_163/Y vdd BUFX4
XBUFX4_152 INVX8_11/Y gnd NOR2X1_2/B vdd BUFX4
XNOR2X1_234 NOR2X1_234/A NOR2X1_236/B gnd NOR2X1_234/Y vdd NOR2X1
XNOR2X1_201 BUFX4_64/Y BUFX4_410/Y gnd NOR2X1_206/B vdd NOR2X1
XNOR2X1_223 NOR2X1_223/A NOR2X1_222/B gnd NOR2X1_223/Y vdd NOR2X1
XNOR2X1_212 NOR2X1_212/A NOR2X1_216/B gnd NOR2X1_212/Y vdd NOR2X1
XBUFX4_174 BUFX4_178/A gnd INVX2_1/A vdd BUFX4
XBUFX4_185 BUFX4_25/Y gnd MUX2X1_9/S vdd BUFX4
XBUFX4_196 BUFX4_25/Y gnd BUFX4_196/Y vdd BUFX4
XNOR2X1_267 NOR2X1_267/A NOR2X1_265/Y gnd NOR2X1_267/Y vdd NOR2X1
XNOR2X1_245 BUFX4_197/Y OR2X2_1/A gnd INVX1_509/A vdd NOR2X1
XNOR2X1_256 DFFPOSX1_9/Q NOR2X1_256/B gnd NOR2X1_256/Y vdd NOR2X1
XFILL_31_1 gnd vdd FILL
XNOR2X1_278 NOR2X1_278/A NOR2X1_279/B gnd NOR2X1_278/Y vdd NOR2X1
XNOR2X1_289 NOR2X1_289/A NOR2X1_289/B gnd NOR2X1_289/Y vdd NOR2X1
XOAI21X1_707 INVX1_118/Y NOR2X1_177/Y OAI21X1_707/C gnd OAI21X1_707/Y vdd OAI21X1
XOAI21X1_718 INVX1_375/Y NOR2X1_189/B NAND2X1_187/Y gnd OAI21X1_718/Y vdd OAI21X1
XOAI21X1_729 BUFX4_130/Y OAI21X1_729/B OAI21X1_728/Y gnd OAI21X1_729/Y vdd OAI21X1
XOAI21X1_1031 INVX1_243/Y BUFX4_250/Y NAND2X1_467/Y gnd MUX2X1_179/B vdd OAI21X1
XOAI21X1_1020 INVX1_232/Y BUFX4_228/Y NAND2X1_455/Y gnd MUX2X1_170/A vdd OAI21X1
XMUX2X1_218 MUX2X1_218/A MUX2X1_218/B BUFX4_6/Y gnd MUX2X1_218/Y vdd MUX2X1
XDFFPOSX1_621 NAND2X1_519/B CLKBUF1_22/Y OAI21X1_370/Y gnd vdd DFFPOSX1
XOAI21X1_1042 INVX1_254/Y BUFX4_272/Y NAND2X1_480/Y gnd MUX2X1_187/A vdd OAI21X1
XDFFPOSX1_632 INVX1_484/A CLKBUF1_60/Y OAI21X1_392/Y gnd vdd DFFPOSX1
XDFFPOSX1_610 INVX1_99/A CLKBUF1_28/Y OAI21X1_348/Y gnd vdd DFFPOSX1
XOAI21X1_1064 INVX1_276/Y BUFX4_217/Y NAND2X1_503/Y gnd MUX2X1_203/A vdd OAI21X1
XOAI21X1_1053 INVX1_265/Y BUFX4_195/Y NAND2X1_491/Y gnd MUX2X1_196/B vdd OAI21X1
XMUX2X1_229 MUX2X1_229/A MUX2X1_229/B BUFX4_58/Y gnd MUX2X1_229/Y vdd MUX2X1
XMUX2X1_207 MUX2X1_207/A MUX2X1_205/Y MUX2X1_42/S gnd AOI22X1_43/A vdd MUX2X1
XDFFPOSX1_665 NAND2X1_264/B CLKBUF1_96/Y OAI21X1_434/Y gnd vdd DFFPOSX1
XOAI21X1_1097 INVX1_309/Y MUX2X1_8/S NAND2X1_538/Y gnd MUX2X1_229/B vdd OAI21X1
XDFFPOSX1_654 NOR2X1_78/A CLKBUF1_33/Y AOI21X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_643 INVX1_165/A CLKBUF1_33/Y OAI21X1_411/Y gnd vdd DFFPOSX1
XOAI21X1_1086 INVX1_298/Y BUFX4_261/Y NAND2X1_526/Y gnd MUX2X1_220/A vdd OAI21X1
XOAI21X1_1075 INVX1_287/Y BUFX4_239/Y NAND2X1_515/Y gnd MUX2X1_212/B vdd OAI21X1
XDFFPOSX1_698 OAI21X1_499/C CLKBUF1_58/Y OAI21X1_500/Y gnd vdd DFFPOSX1
XDFFPOSX1_676 INVX1_231/A CLKBUF1_96/Y OAI21X1_456/Y gnd vdd DFFPOSX1
XDFFPOSX1_687 NAND2X1_661/B CLKBUF1_45/Y OAI21X1_478/Y gnd vdd DFFPOSX1
XNAND2X1_702 AOI22X1_70/Y AOI22X1_71/Y gnd AOI22X1_74/A vdd NAND2X1
XNAND2X1_746 BUFX4_272/Y NOR2X1_187/A gnd NAND2X1_746/Y vdd NAND2X1
XNAND2X1_724 BUFX4_230/Y NOR2X1_70/A gnd NAND2X1_724/Y vdd NAND2X1
XNAND2X1_713 BUFX4_210/Y NAND2X1_713/B gnd NAND2X1_713/Y vdd NAND2X1
XNAND2X1_735 BUFX4_252/Y NOR2X1_110/A gnd NAND2X1_735/Y vdd NAND2X1
XNAND2X1_768 BUFX4_334/Y NOR2X1_264/Y gnd NAND2X1_768/Y vdd NAND2X1
XNAND2X1_757 BUFX4_450/Y NOR2X1_254/Y gnd NAND2X1_757/Y vdd NAND2X1
XNAND2X1_779 BUFX4_448/Y NOR2X1_274/Y gnd NAND2X1_779/Y vdd NAND2X1
XINVX8_5 INVX8_5/A gnd INVX8_5/Y vdd INVX8
XDFFPOSX1_80 NAND2X1_690/B CLKBUF1_42/Y DFFPOSX1_80/D gnd vdd DFFPOSX1
XDFFPOSX1_91 NOR2X1_302/A CLKBUF1_78/Y AOI21X1_241/Y gnd vdd DFFPOSX1
XBUFX4_14 clk gnd BUFX4_14/Y vdd BUFX4
XBUFX4_25 a[0] gnd BUFX4_25/Y vdd BUFX4
XBUFX4_36 BUFX4_78/Y gnd BUFX4_36/Y vdd BUFX4
XBUFX4_47 BUFX4_71/Y gnd BUFX4_47/Y vdd BUFX4
XBUFX4_69 a[1] gnd BUFX4_57/A vdd BUFX4
XBUFX4_58 BUFX4_57/A gnd BUFX4_58/Y vdd BUFX4
XFILL_47_3_1 gnd vdd FILL
XFILL_30_2_1 gnd vdd FILL
XFILL_38_3_1 gnd vdd FILL
XOAI21X1_504 BUFX4_302/Y NAND2X1_97/Y OAI21X1_504/C gnd OAI21X1_504/Y vdd OAI21X1
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_548 INVX1_234/Y NOR2X1_81/Y NAND2X1_104/Y gnd OAI21X1_548/Y vdd OAI21X1
XOAI21X1_537 NOR2X1_2/B BUFX4_295/Y NAND2X1_525/B gnd OAI21X1_538/C vdd OAI21X1
XOAI21X1_526 BUFX4_287/Y NAND2X1_99/Y OAI21X1_525/Y gnd OAI21X1_526/Y vdd OAI21X1
XOAI21X1_515 BUFX4_461/Y INVX1_2/A INVX1_105/A gnd OAI21X1_516/C vdd OAI21X1
XOAI21X1_559 INVX1_427/Y NOR2X1_91/Y OAI21X1_559/C gnd OAI21X1_559/Y vdd OAI21X1
XDFFPOSX1_440 INVX1_472/A CLKBUF1_77/Y OAI21X1_152/Y gnd vdd DFFPOSX1
XDFFPOSX1_462 OAI21X1_195/C CLKBUF1_87/Y OAI21X1_196/Y gnd vdd DFFPOSX1
XDFFPOSX1_451 INVX1_153/A CLKBUF1_50/Y OAI21X1_174/Y gnd vdd DFFPOSX1
XDFFPOSX1_473 NOR2X1_13/A CLKBUF1_44/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_495 NOR2X1_29/A CLKBUF1_2/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_484 INVX1_219/A CLKBUF1_31/Y OAI21X1_212/Y gnd vdd DFFPOSX1
XNAND2X1_510 BUFX4_230/Y NOR2X1_27/A gnd NAND2X1_510/Y vdd NAND2X1
XNAND2X1_521 BUFX4_250/Y NOR2X1_77/A gnd NAND2X1_521/Y vdd NAND2X1
XNAND2X1_543 BUFX4_193/Y NOR2X1_215/A gnd NAND2X1_543/Y vdd NAND2X1
XNAND2X1_532 BUFX4_270/Y NOR2X1_129/A gnd NAND2X1_532/Y vdd NAND2X1
XNAND2X1_554 BUFX4_211/Y NOR2X1_317/A gnd NAND2X1_554/Y vdd NAND2X1
XNAND2X1_587 BUFX4_273/Y OAI21X1_339/C gnd NAND2X1_587/Y vdd NAND2X1
XNAND2X1_565 BUFX4_231/Y NAND2X1_565/B gnd NAND2X1_565/Y vdd NAND2X1
XNAND2X1_576 BUFX4_253/Y OAI21X1_163/C gnd NAND2X1_576/Y vdd NAND2X1
XFILL_4_3_1 gnd vdd FILL
XNAND2X1_598 AOI22X1_55/Y AOI22X1_56/Y gnd AOI22X1_59/A vdd NAND2X1
XFILL_29_3_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XOAI21X1_323 BUFX4_404/Y BUFX4_381/Y INVX1_354/A gnd OAI21X1_323/Y vdd OAI21X1
XOAI21X1_312 INVX1_481/Y NOR2X1_61/Y NAND2X1_76/Y gnd OAI21X1_312/Y vdd OAI21X1
XOAI21X1_301 BUFX4_411/Y BUFX4_433/Y NAND2X1_654/B gnd OAI21X1_301/Y vdd OAI21X1
XOAI21X1_345 NOR2X1_21/B BUFX4_386/Y INVX1_51/A gnd OAI21X1_345/Y vdd OAI21X1
XOAI21X1_334 BUFX4_117/Y NAND2X1_78/Y OAI21X1_333/Y gnd OAI21X1_334/Y vdd OAI21X1
XOAI21X1_356 BUFX4_102/Y NAND2X1_79/Y OAI21X1_355/Y gnd OAI21X1_356/Y vdd OAI21X1
XOAI21X1_378 NAND2X1_81/Y BUFX4_123/Y OAI21X1_377/Y gnd OAI21X1_378/Y vdd OAI21X1
XOAI21X1_389 BUFX4_172/Y BUFX4_384/Y INVX1_420/A gnd OAI21X1_389/Y vdd OAI21X1
XOAI21X1_367 BUFX4_367/Y BUFX4_387/Y NAND2X1_450/B gnd OAI21X1_367/Y vdd OAI21X1
XINVX1_409 INVX1_409/A gnd INVX1_409/Y vdd INVX1
XDFFPOSX1_281 NOR2X1_360/A CLKBUF1_93/Y AOI21X1_286/Y gnd vdd DFFPOSX1
XDFFPOSX1_270 NAND2X1_565/B CLKBUF1_89/Y OAI21X1_1613/Y gnd vdd DFFPOSX1
XDFFPOSX1_292 INVX1_207/A CLKBUF1_102/Y OAI21X1_1629/Y gnd vdd DFFPOSX1
XNAND2X1_362 BUFX4_251/Y NOR2X1_382/A gnd NAND2X1_362/Y vdd NAND2X1
XNAND2X1_340 AOI22X1_14/Y AOI22X1_19/Y gnd NAND2X1_340/Y vdd NAND2X1
XNAND2X1_351 BUFX4_231/Y NOR2X1_335/A gnd OAI21X1_923/C vdd NAND2X1
XNAND2X1_384 BUFX4_194/Y NAND2X1_384/B gnd NAND2X1_384/Y vdd NAND2X1
XNAND2X1_395 BUFX4_214/Y NOR2X1_138/A gnd NAND2X1_395/Y vdd NAND2X1
XNAND2X1_373 BUFX4_273/Y NOR2X1_35/A gnd OAI21X1_944/C vdd NAND2X1
XFILL_44_1_1 gnd vdd FILL
XOAI21X1_1619 INVX1_78/Y NOR2X1_358/Y NAND2X1_845/Y gnd OAI21X1_1619/Y vdd OAI21X1
XOAI21X1_1608 NOR2X1_2/B BUFX4_346/Y NAND2X1_427/B gnd OAI21X1_1609/C vdd OAI21X1
XOAI21X1_890 INVX1_102/Y BUFX4_265/Y OAI21X1_890/C gnd MUX2X1_73/A vdd OAI21X1
XFILL_49_2 gnd vdd FILL
XFILL_35_1_1 gnd vdd FILL
XNAND3X1_2 NAND3X1_2/A NAND3X1_2/B AOI22X1_2/Y gnd NAND3X1_2/Y vdd NAND3X1
XFILL_1_1_1 gnd vdd FILL
XFILL_26_1_1 gnd vdd FILL
XOAI21X1_120 BUFX4_379/Y NAND2X1_16/Y OAI21X1_120/C gnd OAI21X1_120/Y vdd OAI21X1
XOAI21X1_131 NOR2X1_52/B BUFX4_178/Y OAI21X1_131/C gnd OAI21X1_131/Y vdd OAI21X1
XAOI22X1_7 AOI22X1_7/A AOI22X1_7/B AOI22X1_7/C MUX2X1_36/Y gnd AOI22X1_7/Y vdd AOI22X1
XOAI21X1_153 NOR2X1_32/B NOR2X1_2/A OAI21X1_153/C gnd OAI21X1_154/C vdd OAI21X1
XOAI21X1_164 AOI21X1_6/A NAND2X1_19/Y OAI21X1_163/Y gnd OAI21X1_164/Y vdd OAI21X1
XOAI21X1_142 NAND2X1_18/Y BUFX4_114/Y OAI21X1_141/Y gnd OAI21X1_142/Y vdd OAI21X1
XOAI21X1_186 BUFX4_131/Y NAND2X1_22/Y OAI21X1_186/C gnd OAI21X1_186/Y vdd OAI21X1
XOAI21X1_175 NOR2X1_61/B BUFX4_133/Y INVX1_217/A gnd OAI21X1_175/Y vdd OAI21X1
XOAI21X1_197 NOR2X1_2/B BUFX4_133/Y NAND2X1_646/B gnd OAI21X1_198/C vdd OAI21X1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XINVX1_206 INVX1_206/A gnd INVX1_206/Y vdd INVX1
XINVX1_228 INVX1_228/A gnd INVX1_228/Y vdd INVX1
XINVX1_239 INVX1_239/A gnd INVX1_239/Y vdd INVX1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_28 BUFX4_327/Y NOR2X1_11/Y gnd NAND2X1_28/Y vdd NAND2X1
XNAND2X1_39 BUFX4_164/Y NOR2X1_31/Y gnd NAND2X1_39/Y vdd NAND2X1
XNAND2X1_17 INVX2_1/Y INVX8_15/A gnd NAND2X1_17/Y vdd NAND2X1
XNAND2X1_170 BUFX4_327/Y NOR2X1_166/Y gnd NAND2X1_170/Y vdd NAND2X1
XNAND2X1_181 INVX8_8/A NOR2X1_177/Y gnd NAND2X1_181/Y vdd NAND2X1
XNAND2X1_192 BUFX4_145/Y NOR2X1_199/Y gnd OAI21X1_723/C vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_15 MUX2X1_69/Y BUFX4_352/Y BUFX4_157/Y MUX2X1_72/Y gnd AOI22X1_15/Y vdd AOI22X1
XAOI22X1_48 MUX2X1_231/Y INVX1_10/A INVX1_11/A MUX2X1_234/Y gnd AOI22X1_48/Y vdd AOI22X1
XAOI22X1_26 MUX2X1_123/Y BUFX4_320/Y INVX1_11/A AOI22X1_26/D gnd AOI22X1_26/Y vdd
+ AOI22X1
XAOI22X1_37 MUX2X1_177/Y INVX1_6/A INVX1_8/A AOI22X1_37/D gnd AOI22X1_37/Y vdd AOI22X1
XOAI21X1_1405 BUFX4_416/Y BUFX4_466/Y NAND2X1_624/B gnd OAI21X1_1405/Y vdd OAI21X1
XAOI22X1_59 AOI22X1_59/A AOI22X1_9/D AOI22X1_69/C AOI22X1_59/D gnd AOI22X1_59/Y vdd
+ AOI22X1
XOAI21X1_1416 BUFX4_304/Y NAND2X1_814/Y OAI21X1_1416/C gnd DFFPOSX1_132/D vdd OAI21X1
XOAI21X1_1427 BUFX4_151/Y BUFX4_389/Y NAND2X1_280/B gnd OAI21X1_1427/Y vdd OAI21X1
XOAI21X1_1438 BUFX4_286/Y NAND2X1_815/Y OAI21X1_1437/Y gnd OAI21X1_1438/Y vdd OAI21X1
XOAI21X1_1449 INVX1_43/Y NOR2X1_331/Y NAND2X1_824/Y gnd OAI21X1_1449/Y vdd OAI21X1
XFILL_20_8_0 gnd vdd FILL
XFILL_11_8_0 gnd vdd FILL
XAOI21X1_70 BUFX4_103/Y NOR2X1_90/B NOR2X1_88/Y gnd AOI21X1_70/Y vdd AOI21X1
XAOI21X1_92 BUFX4_110/Y NOR2X1_118/B NOR2X1_116/Y gnd AOI21X1_92/Y vdd AOI21X1
XAOI21X1_81 BUFX4_126/Y NOR2X1_103/B AOI21X1_81/C gnd AOI21X1_81/Y vdd AOI21X1
XBUFX4_312 INVX8_14/Y gnd BUFX4_312/Y vdd BUFX4
XBUFX4_301 INVX8_5/Y gnd BUFX4_301/Y vdd BUFX4
XBUFX4_323 BUFX4_321/A gnd BUFX4_323/Y vdd BUFX4
XBUFX4_334 d[2] gnd BUFX4_334/Y vdd BUFX4
XBUFX4_345 BUFX4_344/A gnd BUFX4_345/Y vdd BUFX4
XBUFX4_367 INVX8_15/Y gnd BUFX4_367/Y vdd BUFX4
XBUFX4_378 INVX8_9/Y gnd BUFX4_378/Y vdd BUFX4
XBUFX4_356 a[2] gnd MUX2X1_69/S vdd BUFX4
XBUFX4_389 BUFX4_392/A gnd BUFX4_389/Y vdd BUFX4
XOAI21X1_1213 INVX1_425/Y BUFX4_218/Y NAND2X1_663/Y gnd MUX2X1_316/B vdd OAI21X1
XOAI21X1_1202 INVX1_414/Y BUFX4_196/Y NAND2X1_652/Y gnd MUX2X1_307/A vdd OAI21X1
XOAI21X1_1246 INVX1_458/Y MUX2X1_9/S NAND2X1_699/Y gnd MUX2X1_340/A vdd OAI21X1
XOAI21X1_1235 INVX1_447/Y BUFX4_262/Y NAND2X1_688/Y gnd MUX2X1_332/B vdd OAI21X1
XDFFPOSX1_814 NOR2X1_130/A CLKBUF1_40/Y AOI21X1_104/Y gnd vdd DFFPOSX1
XDFFPOSX1_803 INVX1_175/A CLKBUF1_100/Y OAI21X1_609/Y gnd vdd DFFPOSX1
XOAI21X1_1224 INVX1_436/Y BUFX4_240/Y NAND2X1_675/Y gnd MUX2X1_323/A vdd OAI21X1
XDFFPOSX1_836 INVX1_241/A CLKBUF1_15/Y OAI21X1_629/Y gnd vdd DFFPOSX1
XDFFPOSX1_847 NAND2X1_672/B CLKBUF1_15/Y OAI21X1_651/Y gnd vdd DFFPOSX1
XDFFPOSX1_825 MUX2X1_5/A CLKBUF1_96/Y AOI21X1_108/Y gnd vdd DFFPOSX1
XOAI21X1_1257 INVX1_469/Y BUFX4_207/Y NAND2X1_711/Y gnd MUX2X1_349/B vdd OAI21X1
XOAI21X1_1279 INVX1_491/Y BUFX4_251/Y NAND2X1_734/Y gnd MUX2X1_365/B vdd OAI21X1
XOAI21X1_1268 INVX1_480/Y BUFX4_229/Y NAND2X1_723/Y gnd MUX2X1_356/A vdd OAI21X1
XDFFPOSX1_869 INVX1_307/A CLKBUF1_91/Y OAI21X1_664/Y gnd vdd DFFPOSX1
XDFFPOSX1_858 NOR2X1_148/A CLKBUF1_54/Y AOI21X1_118/Y gnd vdd DFFPOSX1
XFILL_6_0_1 gnd vdd FILL
XFILL_43_7_0 gnd vdd FILL
XMUX2X1_3 MUX2X1_3/A MUX2X1_3/B MUX2X1_3/S gnd MUX2X1_7/B vdd MUX2X1
XCLKBUF1_4 BUFX4_13/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XBUFX4_120 BUFX4_121/A gnd BUFX4_120/Y vdd BUFX4
XBUFX4_131 INVX8_2/Y gnd BUFX4_131/Y vdd BUFX4
XBUFX4_142 d[3] gnd BUFX4_142/Y vdd BUFX4
XBUFX4_164 d[0] gnd BUFX4_164/Y vdd BUFX4
XBUFX4_153 INVX8_11/Y gnd BUFX4_153/Y vdd BUFX4
XBUFX4_197 BUFX4_24/Y gnd BUFX4_197/Y vdd BUFX4
XNOR2X1_202 MUX2X1_19/A NOR2X1_206/B gnd NOR2X1_202/Y vdd NOR2X1
XNOR2X1_224 NOR2X1_224/A NOR2X1_222/B gnd NOR2X1_224/Y vdd NOR2X1
XNOR2X1_213 NOR2X1_213/A NOR2X1_216/B gnd NOR2X1_213/Y vdd NOR2X1
XBUFX4_175 BUFX4_178/A gnd BUFX4_175/Y vdd BUFX4
XBUFX4_186 BUFX4_27/Y gnd MUX2X1_11/S vdd BUFX4
XNOR2X1_235 NOR2X1_235/A NOR2X1_236/B gnd NOR2X1_235/Y vdd NOR2X1
XNOR2X1_257 NOR2X1_257/A NOR2X1_256/B gnd NOR2X1_257/Y vdd NOR2X1
XNOR2X1_246 NOR2X1_246/A OAI22X1_3/Y gnd NOR2X1_246/Y vdd NOR2X1
XFILL_31_2 gnd vdd FILL
XFILL_34_7_0 gnd vdd FILL
XNOR2X1_268 NOR2X1_268/A NOR2X1_265/Y gnd NOR2X1_268/Y vdd NOR2X1
XNOR2X1_279 NOR2X1_279/A NOR2X1_279/B gnd NOR2X1_279/Y vdd NOR2X1
XFILL_24_1 gnd vdd FILL
XOAI21X1_708 INVX1_182/Y NOR2X1_177/Y OAI21X1_708/C gnd OAI21X1_708/Y vdd OAI21X1
XOAI21X1_719 INVX1_439/Y NOR2X1_189/B OAI21X1_719/C gnd OAI21X1_719/Y vdd OAI21X1
XOAI21X1_1021 INVX1_233/Y BUFX4_230/Y NAND2X1_456/Y gnd MUX2X1_172/B vdd OAI21X1
XOAI21X1_1010 INVX1_222/Y BUFX4_208/Y NAND2X1_445/Y gnd MUX2X1_163/A vdd OAI21X1
XOAI21X1_1032 INVX1_244/Y BUFX4_252/Y NAND2X1_468/Y gnd MUX2X1_179/A vdd OAI21X1
XDFFPOSX1_600 INVX1_482/A CLKBUF1_79/Y OAI21X1_328/Y gnd vdd DFFPOSX1
XOAI21X1_1054 INVX1_266/Y BUFX4_197/Y NAND2X1_492/Y gnd MUX2X1_196/A vdd OAI21X1
XDFFPOSX1_622 NAND2X1_588/B CLKBUF1_60/Y OAI21X1_372/Y gnd vdd DFFPOSX1
XDFFPOSX1_611 INVX1_163/A CLKBUF1_34/Y OAI21X1_350/Y gnd vdd DFFPOSX1
XMUX2X1_208 MUX2X1_208/A MUX2X1_208/B BUFX4_20/Y gnd MUX2X1_208/Y vdd MUX2X1
XOAI21X1_1043 INVX1_255/Y BUFX4_274/Y NAND2X1_481/Y gnd MUX2X1_188/B vdd OAI21X1
XMUX2X1_219 MUX2X1_218/Y MUX2X1_217/Y BUFX4_362/Y gnd AOI22X1_46/A vdd MUX2X1
XOAI21X1_1098 INVX1_310/Y MUX2X1_11/S NAND2X1_539/Y gnd MUX2X1_229/A vdd OAI21X1
XDFFPOSX1_666 NAND2X1_315/B CLKBUF1_58/Y OAI21X1_436/Y gnd vdd DFFPOSX1
XDFFPOSX1_633 OAI21X1_393/C CLKBUF1_97/Y OAI21X1_394/Y gnd vdd DFFPOSX1
XDFFPOSX1_644 INVX1_229/A CLKBUF1_69/Y OAI21X1_412/Y gnd vdd DFFPOSX1
XDFFPOSX1_655 NOR2X1_79/A CLKBUF1_100/Y AOI21X1_63/Y gnd vdd DFFPOSX1
XOAI21X1_1087 INVX1_299/Y BUFX4_263/Y NAND2X1_527/Y gnd MUX2X1_221/B vdd OAI21X1
XOAI21X1_1065 INVX1_277/Y BUFX4_219/Y NAND2X1_504/Y gnd MUX2X1_205/B vdd OAI21X1
XOAI21X1_1076 INVX1_288/Y BUFX4_241/Y NAND2X1_516/Y gnd MUX2X1_212/A vdd OAI21X1
XDFFPOSX1_688 NAND2X1_730/B CLKBUF1_70/Y OAI21X1_480/Y gnd vdd DFFPOSX1
XDFFPOSX1_677 INVX1_295/A CLKBUF1_99/Y OAI21X1_458/Y gnd vdd DFFPOSX1
XDFFPOSX1_699 OAI21X1_501/C CLKBUF1_97/Y OAI21X1_502/Y gnd vdd DFFPOSX1
XNAND2X1_703 BUFX4_190/Y NAND2X1_703/B gnd NAND2X1_703/Y vdd NAND2X1
XNAND2X1_725 BUFX4_232/Y NAND2X1_725/B gnd NAND2X1_725/Y vdd NAND2X1
XNAND2X1_736 AOI22X1_75/Y AOI22X1_76/Y gnd AOI22X1_79/A vdd NAND2X1
XNAND2X1_714 BUFX4_212/Y NAND2X1_714/B gnd NAND2X1_714/Y vdd NAND2X1
XNAND2X1_747 BUFX4_274/Y NOR2X1_198/A gnd NAND2X1_747/Y vdd NAND2X1
XNAND2X1_758 BUFX4_332/Y NOR2X1_254/Y gnd NAND2X1_758/Y vdd NAND2X1
XNAND2X1_769 BUFX4_144/Y NOR2X1_264/Y gnd NAND2X1_769/Y vdd NAND2X1
XFILL_0_7_0 gnd vdd FILL
XFILL_25_7_0 gnd vdd FILL
XINVX8_6 INVX8_6/A gnd INVX8_6/Y vdd INVX8
XDFFPOSX1_81 INVX1_38/A CLKBUF1_17/Y DFFPOSX1_81/D gnd vdd DFFPOSX1
XDFFPOSX1_70 INVX1_321/A CLKBUF1_17/Y DFFPOSX1_70/D gnd vdd DFFPOSX1
XDFFPOSX1_92 NOR2X1_303/A CLKBUF1_78/Y AOI21X1_242/Y gnd vdd DFFPOSX1
XFILL_8_8_0 gnd vdd FILL
XBUFX4_15 clk gnd BUFX4_15/Y vdd BUFX4
XBUFX4_26 a[0] gnd BUFX4_26/Y vdd BUFX4
XBUFX4_37 BUFX4_78/Y gnd BUFX4_37/Y vdd BUFX4
XBUFX4_48 BUFX4_50/A gnd BUFX4_48/Y vdd BUFX4
XBUFX4_59 BUFX4_57/A gnd BUFX4_59/Y vdd BUFX4
XFILL_16_7_0 gnd vdd FILL
XOAI21X1_505 BUFX4_414/Y INVX2_4/A NAND2X1_524/B gnd OAI21X1_506/C vdd OAI21X1
XOAI21X1_527 BUFX4_456/Y BUFX4_293/Y INVX1_489/A gnd OAI21X1_528/C vdd OAI21X1
XOAI21X1_538 BUFX4_396/Y OAI21X1_544/B OAI21X1_538/C gnd OAI21X1_538/Y vdd OAI21X1
XOAI21X1_516 BUFX4_418/Y NAND2X1_99/Y OAI21X1_516/C gnd OAI21X1_516/Y vdd OAI21X1
XOAI21X1_549 INVX1_298/Y NOR2X1_81/Y OAI21X1_549/C gnd OAI21X1_549/Y vdd OAI21X1
XDFFPOSX1_430 OAI21X1_131/C CLKBUF1_41/Y OAI21X1_132/Y gnd vdd DFFPOSX1
XDFFPOSX1_452 INVX1_217/A CLKBUF1_5/Y OAI21X1_176/Y gnd vdd DFFPOSX1
XDFFPOSX1_463 NAND2X1_646/B CLKBUF1_56/Y OAI21X1_198/Y gnd vdd DFFPOSX1
XDFFPOSX1_474 NOR2X1_14/A CLKBUF1_44/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_441 OAI21X1_153/C CLKBUF1_30/Y OAI21X1_154/Y gnd vdd DFFPOSX1
XNAND2X1_500 BUFX4_210/Y NOR2X1_384/A gnd NAND2X1_500/Y vdd NAND2X1
XDFFPOSX1_496 NOR2X1_30/A CLKBUF1_2/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XNAND2X1_511 BUFX4_232/Y NOR2X1_37/A gnd NAND2X1_511/Y vdd NAND2X1
XDFFPOSX1_485 INVX1_283/A CLKBUF1_93/Y OAI21X1_213/Y gnd vdd DFFPOSX1
XNAND2X1_533 BUFX4_272/Y NOR2X1_140/A gnd NAND2X1_533/Y vdd NAND2X1
XNAND2X1_522 BUFX4_252/Y NAND2X1_522/B gnd NAND2X1_522/Y vdd NAND2X1
XNAND2X1_544 BUFX4_195/Y NOR2X1_224/A gnd NAND2X1_544/Y vdd NAND2X1
XNAND2X1_588 BUFX4_275/Y NAND2X1_588/B gnd NAND2X1_588/Y vdd NAND2X1
XNAND2X1_577 BUFX4_255/Y OAI21X1_195/C gnd NAND2X1_577/Y vdd NAND2X1
XNAND2X1_555 BUFX4_213/Y NAND2X1_555/B gnd NAND2X1_555/Y vdd NAND2X1
XNAND2X1_566 BUFX4_233/Y NOR2X1_365/A gnd NAND2X1_566/Y vdd NAND2X1
XNAND2X1_599 BUFX4_196/Y OAI21X1_595/C gnd NAND2X1_599/Y vdd NAND2X1
XFILL_40_5_0 gnd vdd FILL
XAOI21X1_190 BUFX4_300/Y NOR2X1_236/B NOR2X1_234/Y gnd AOI21X1_190/Y vdd AOI21X1
XFILL_48_6_0 gnd vdd FILL
XFILL_31_5_0 gnd vdd FILL
XFILL_39_6_0 gnd vdd FILL
XFILL_22_5_0 gnd vdd FILL
XOAI21X1_313 BUFX4_404/Y BUFX4_387/Y INVX1_50/A gnd OAI21X1_314/C vdd OAI21X1
XOAI21X1_302 BUFX4_287/Y NAND2X1_67/Y OAI21X1_301/Y gnd OAI21X1_302/Y vdd OAI21X1
XOAI21X1_324 BUFX4_102/Y NAND2X1_77/Y OAI21X1_323/Y gnd OAI21X1_324/Y vdd OAI21X1
XOAI21X1_335 BUFX4_85/Y BUFX4_381/Y OAI21X1_335/C gnd OAI21X1_336/C vdd OAI21X1
XOAI21X1_346 BUFX4_123/Y NAND2X1_79/Y OAI21X1_345/Y gnd OAI21X1_346/Y vdd OAI21X1
XOAI21X1_379 BUFX4_172/Y BUFX4_384/Y INVX1_100/A gnd OAI21X1_380/C vdd OAI21X1
XOAI21X1_368 BUFX4_303/Y NAND2X1_80/Y OAI21X1_367/Y gnd OAI21X1_368/Y vdd OAI21X1
XOAI21X1_357 BUFX4_308/Y BUFX4_385/Y INVX1_419/A gnd OAI21X1_357/Y vdd OAI21X1
XDFFPOSX1_282 NOR2X1_361/A CLKBUF1_93/Y AOI21X1_287/Y gnd vdd DFFPOSX1
XDFFPOSX1_271 NAND2X1_634/B CLKBUF1_12/Y OAI21X1_1615/Y gnd vdd DFFPOSX1
XDFFPOSX1_260 INVX1_205/A CLKBUF1_48/Y DFFPOSX1_260/D gnd vdd DFFPOSX1
XDFFPOSX1_293 INVX1_271/A CLKBUF1_25/Y OAI21X1_1630/Y gnd vdd DFFPOSX1
XNAND2X1_352 BUFX4_233/Y NAND2X1_352/B gnd NAND2X1_352/Y vdd NAND2X1
XNAND2X1_363 BUFX4_253/Y NAND2X1_363/B gnd NAND2X1_363/Y vdd NAND2X1
XNAND2X1_341 BUFX4_211/Y NOR2X1_258/A gnd NAND2X1_341/Y vdd NAND2X1
XNAND2X1_330 BUFX4_193/Y NOR2X1_170/A gnd OAI21X1_904/C vdd NAND2X1
XNAND2X1_385 BUFX4_196/Y NAND2X1_385/B gnd NAND2X1_385/Y vdd NAND2X1
XFILL_5_6_0 gnd vdd FILL
XNAND2X1_374 AOI22X1_22/Y AOI22X1_23/Y gnd AOI22X1_24/D vdd NAND2X1
XNAND2X1_396 BUFX4_216/Y OAI21X1_642/C gnd OAI21X1_965/C vdd NAND2X1
XFILL_13_5_0 gnd vdd FILL
XOAI21X1_1609 BUFX4_297/Y NAND2X1_843/Y OAI21X1_1609/C gnd DFFPOSX1_268/D vdd OAI21X1
XOAI21X1_880 INVX1_92/Y BUFX4_245/Y OAI21X1_880/C gnd MUX2X1_65/A vdd OAI21X1
XOAI21X1_891 INVX1_103/Y BUFX4_267/Y NAND2X1_316/Y gnd MUX2X1_74/B vdd OAI21X1
XFILL_49_3 gnd vdd FILL
XNAND3X1_3 NAND3X1_3/A NAND3X1_3/B NAND3X1_3/C gnd AOI22X1_6/A vdd NAND3X1
XOAI21X1_121 BUFX4_371/Y BUFX4_179/Y OAI21X1_121/C gnd OAI21X1_122/C vdd OAI21X1
XOAI21X1_110 BUFX4_116/Y NAND2X1_16/Y OAI21X1_110/C gnd OAI21X1_110/Y vdd OAI21X1
XAOI22X1_8 MUX2X1_39/Y BUFX4_320/Y INVX1_11/A AOI22X1_8/D gnd AOI22X1_8/Y vdd AOI22X1
XOAI21X1_154 BUFX4_127/Y NAND2X1_19/Y OAI21X1_154/C gnd OAI21X1_154/Y vdd OAI21X1
XOAI21X1_165 NOR2X1_32/B BUFX4_175/Y NAND2X1_645/B gnd OAI21X1_165/Y vdd OAI21X1
XOAI21X1_132 AOI21X1_6/A NAND2X1_17/Y OAI21X1_131/Y gnd OAI21X1_132/Y vdd OAI21X1
XOAI21X1_143 INVX4_3/A BUFX4_173/Y INVX1_216/A gnd OAI21X1_144/C vdd OAI21X1
XOAI21X1_176 BUFX4_301/Y NAND2X1_21/Y OAI21X1_175/Y gnd OAI21X1_176/Y vdd OAI21X1
XOAI21X1_198 BUFX4_282/Y NAND2X1_22/Y OAI21X1_198/C gnd OAI21X1_198/Y vdd OAI21X1
XOAI21X1_187 NOR2X1_2/B BUFX4_134/Y OAI21X1_187/C gnd OAI21X1_187/Y vdd OAI21X1
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XINVX1_218 INVX1_218/A gnd INVX1_218/Y vdd INVX1
XINVX1_229 INVX1_229/A gnd INVX1_229/Y vdd INVX1
XNAND2X1_160 NAND2X1_8/A NOR2X1_155/Y gnd OAI21X1_662/C vdd NAND2X1
XNAND2X1_29 BUFX4_137/Y NOR2X1_11/Y gnd NAND2X1_29/Y vdd NAND2X1
XNAND2X1_18 INVX2_1/Y INVX4_3/Y gnd NAND2X1_18/Y vdd NAND2X1
XNAND2X1_171 BUFX4_137/Y NOR2X1_166/Y gnd NAND2X1_171/Y vdd NAND2X1
XNAND2X1_182 INVX8_9/A NOR2X1_177/Y gnd OAI21X1_713/C vdd NAND2X1
XNAND2X1_193 BUFX4_448/Y NOR2X1_199/Y gnd NAND2X1_193/Y vdd NAND2X1
XFILL_45_4_0 gnd vdd FILL
XAOI22X1_38 MUX2X1_183/Y BUFX4_322/Y BUFX4_292/Y AOI22X1_38/D gnd AOI22X1_38/Y vdd
+ AOI22X1
XAOI22X1_16 MUX2X1_75/Y BUFX4_322/Y BUFX4_292/Y MUX2X1_78/Y gnd AOI22X1_16/Y vdd AOI22X1
XAOI22X1_27 AOI22X1_27/A AOI22X1_7/B AOI22X1_7/C AOI22X1_27/D gnd AOI22X1_27/Y vdd
+ AOI22X1
XAOI22X1_49 AOI22X1_49/A AOI22X1_9/D AOI22X1_69/C AOI22X1_49/D gnd AOI22X1_49/Y vdd
+ AOI22X1
XOAI21X1_1428 BUFX4_420/Y NAND2X1_815/Y OAI21X1_1427/Y gnd DFFPOSX1_138/D vdd OAI21X1
XOAI21X1_1406 BUFX4_279/Y NAND2X1_812/Y OAI21X1_1405/Y gnd DFFPOSX1_127/D vdd OAI21X1
XOAI21X1_1417 BUFX4_457/Y BUFX4_389/Y INVX1_261/A gnd OAI21X1_1417/Y vdd OAI21X1
XOAI21X1_1439 BUFX4_154/Y INVX2_8/A NAND2X1_694/B gnd OAI21X1_1439/Y vdd OAI21X1
XFILL_36_4_0 gnd vdd FILL
XFILL_20_8_1 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XFILL_27_4_0 gnd vdd FILL
XFILL_11_8_1 gnd vdd FILL
XFILL_10_3_0 gnd vdd FILL
XAOI21X1_60 BUFX4_298/Y NOR2X1_77/B NOR2X1_76/Y gnd AOI21X1_60/Y vdd AOI21X1
XAOI21X1_71 BUFX4_281/Y NOR2X1_90/B NOR2X1_89/Y gnd AOI21X1_71/Y vdd AOI21X1
XAOI21X1_93 BUFX4_298/Y NOR2X1_118/B AOI21X1_93/C gnd AOI21X1_93/Y vdd AOI21X1
XAOI21X1_82 BUFX4_422/Y NOR2X1_103/B NOR2X1_104/Y gnd AOI21X1_82/Y vdd AOI21X1
XBUFX4_302 INVX8_5/Y gnd BUFX4_302/Y vdd BUFX4
XBUFX4_313 BUFX4_316/A gnd OAI21X1_1/B vdd BUFX4
XBUFX4_324 BUFX4_321/A gnd BUFX4_324/Y vdd BUFX4
XBUFX4_335 d[2] gnd BUFX4_335/Y vdd BUFX4
XBUFX4_346 BUFX4_344/A gnd BUFX4_346/Y vdd BUFX4
XBUFX4_368 INVX8_15/Y gnd BUFX4_368/Y vdd BUFX4
XFILL_18_4_0 gnd vdd FILL
XBUFX4_357 a[2] gnd BUFX4_357/Y vdd BUFX4
XBUFX4_379 INVX8_9/Y gnd BUFX4_379/Y vdd BUFX4
XOAI21X1_1203 INVX1_415/Y INVX8_1/A NAND2X1_653/Y gnd MUX2X1_308/B vdd OAI21X1
XOAI21X1_1225 INVX1_437/Y BUFX4_242/Y NAND2X1_676/Y gnd MUX2X1_325/B vdd OAI21X1
XOAI21X1_1247 INVX1_459/Y MUX2X1_12/S NAND2X1_700/Y gnd MUX2X1_341/B vdd OAI21X1
XOAI21X1_1236 INVX1_448/Y BUFX4_264/Y NAND2X1_689/Y gnd MUX2X1_332/A vdd OAI21X1
XDFFPOSX1_815 NOR2X1_131/A CLKBUF1_93/Y AOI21X1_105/Y gnd vdd DFFPOSX1
XDFFPOSX1_804 INVX1_239/A CLKBUF1_61/Y OAI21X1_610/Y gnd vdd DFFPOSX1
XOAI21X1_1214 INVX1_426/Y BUFX4_220/Y NAND2X1_664/Y gnd MUX2X1_316/A vdd OAI21X1
XDFFPOSX1_837 INVX1_305/A CLKBUF1_15/Y OAI21X1_631/Y gnd vdd DFFPOSX1
XDFFPOSX1_848 NAND2X1_741/B CLKBUF1_81/Y OAI21X1_653/Y gnd vdd DFFPOSX1
XDFFPOSX1_826 NOR2X1_137/A CLKBUF1_99/Y AOI21X1_109/Y gnd vdd DFFPOSX1
XOAI21X1_1269 INVX1_481/Y BUFX4_231/Y NAND2X1_724/Y gnd MUX2X1_358/B vdd OAI21X1
XOAI21X1_1258 INVX1_470/Y BUFX4_209/Y NAND2X1_712/Y gnd MUX2X1_349/A vdd OAI21X1
XDFFPOSX1_859 NOR2X1_149/A CLKBUF1_95/Y AOI21X1_119/Y gnd vdd DFFPOSX1
XFILL_43_7_1 gnd vdd FILL
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_4/S gnd MUX2X1_6/B vdd MUX2X1
XFILL_42_2_0 gnd vdd FILL
XCLKBUF1_5 BUFX4_17/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XBUFX4_121 BUFX4_121/A gnd BUFX4_121/Y vdd BUFX4
XBUFX4_110 INVX8_4/Y gnd BUFX4_110/Y vdd BUFX4
XBUFX4_132 BUFX4_135/A gnd INVX1_1/A vdd BUFX4
XBUFX4_143 d[3] gnd INVX8_5/A vdd BUFX4
XBUFX4_154 INVX8_11/Y gnd BUFX4_154/Y vdd BUFX4
XBUFX4_165 BUFX4_168/A gnd BUFX4_165/Y vdd BUFX4
XNOR2X1_203 NOR2X1_203/A NOR2X1_206/B gnd NOR2X1_203/Y vdd NOR2X1
XNOR2X1_225 NOR2X1_225/A NOR2X1_222/B gnd NOR2X1_225/Y vdd NOR2X1
XNOR2X1_214 NOR2X1_214/A NOR2X1_216/B gnd NOR2X1_214/Y vdd NOR2X1
XBUFX4_176 BUFX4_178/A gnd NOR2X1_1/A vdd BUFX4
XBUFX4_187 BUFX4_25/Y gnd MUX2X1_12/S vdd BUFX4
XNOR2X1_247 BUFX4_36/Y MUX2X1_29/Y gnd NOR2X1_247/Y vdd NOR2X1
XNOR2X1_258 NOR2X1_258/A NOR2X1_256/B gnd NOR2X1_258/Y vdd NOR2X1
XNOR2X1_236 NOR2X1_236/A NOR2X1_236/B gnd NOR2X1_236/Y vdd NOR2X1
XBUFX4_198 BUFX4_26/Y gnd INVX8_1/A vdd BUFX4
XFILL_34_7_1 gnd vdd FILL
XNOR2X1_269 NOR2X1_269/A NOR2X1_265/Y gnd NOR2X1_269/Y vdd NOR2X1
XFILL_33_2_0 gnd vdd FILL
XFILL_17_1 gnd vdd FILL
XOAI21X1_709 INVX1_246/Y NOR2X1_177/Y OAI21X1_709/C gnd OAI21X1_709/Y vdd OAI21X1
XOAI21X1_1000 INVX1_212/Y BUFX4_188/Y NAND2X1_434/Y gnd MUX2X1_155/A vdd OAI21X1
XOAI21X1_1022 INVX1_234/Y BUFX4_232/Y NAND2X1_457/Y gnd MUX2X1_172/A vdd OAI21X1
XOAI21X1_1011 INVX1_223/Y BUFX4_210/Y NAND2X1_446/Y gnd MUX2X1_164/B vdd OAI21X1
XDFFPOSX1_623 NAND2X1_657/B CLKBUF1_79/Y OAI21X1_374/Y gnd vdd DFFPOSX1
XOAI21X1_1055 INVX1_267/Y BUFX4_199/Y NAND2X1_493/Y gnd MUX2X1_197/B vdd OAI21X1
XDFFPOSX1_601 NAND2X1_260/B CLKBUF1_60/Y OAI21X1_330/Y gnd vdd DFFPOSX1
XOAI21X1_1033 INVX1_245/Y BUFX4_254/Y NAND2X1_469/Y gnd MUX2X1_181/B vdd OAI21X1
XDFFPOSX1_612 INVX1_227/A CLKBUF1_8/Y OAI21X1_352/Y gnd vdd DFFPOSX1
XOAI21X1_1044 INVX1_256/Y BUFX4_276/Y NAND2X1_482/Y gnd MUX2X1_188/A vdd OAI21X1
XMUX2X1_209 MUX2X1_209/A MUX2X1_209/B BUFX4_45/Y gnd MUX2X1_210/A vdd MUX2X1
XDFFPOSX1_634 NAND2X1_313/B CLKBUF1_60/Y OAI21X1_396/Y gnd vdd DFFPOSX1
XOAI21X1_1077 INVX1_289/Y BUFX4_243/Y NAND2X1_517/Y gnd MUX2X1_214/B vdd OAI21X1
XDFFPOSX1_656 NOR2X1_80/A CLKBUF1_59/Y AOI21X1_64/Y gnd vdd DFFPOSX1
XDFFPOSX1_645 INVX1_293/A CLKBUF1_88/Y OAI21X1_413/Y gnd vdd DFFPOSX1
XOAI21X1_1088 INVX1_300/Y BUFX4_265/Y NAND2X1_528/Y gnd MUX2X1_221/A vdd OAI21X1
XOAI21X1_1066 INVX1_278/Y BUFX4_221/Y NAND2X1_505/Y gnd MUX2X1_205/A vdd OAI21X1
XOAI21X1_1099 INVX1_311/Y BUFX4_188/Y NAND2X1_540/Y gnd MUX2X1_230/B vdd OAI21X1
XDFFPOSX1_678 INVX1_359/A CLKBUF1_96/Y OAI21X1_460/Y gnd vdd DFFPOSX1
XDFFPOSX1_689 INVX1_56/A CLKBUF1_45/Y OAI21X1_482/Y gnd vdd DFFPOSX1
XDFFPOSX1_667 NAND2X1_384/B CLKBUF1_58/Y OAI21X1_438/Y gnd vdd DFFPOSX1
XNAND2X1_726 BUFX4_234/Y OAI21X1_375/C gnd NAND2X1_726/Y vdd NAND2X1
XNAND2X1_715 BUFX4_214/Y NAND2X1_715/B gnd NAND2X1_715/Y vdd NAND2X1
XNAND2X1_737 BUFX4_254/Y NAND2X1_737/B gnd NAND2X1_737/Y vdd NAND2X1
XNAND2X1_704 BUFX4_192/Y NOR2X1_367/A gnd NAND2X1_704/Y vdd NAND2X1
XINVX1_390 INVX1_390/A gnd INVX1_390/Y vdd INVX1
XNAND2X1_748 BUFX4_276/Y NOR2X1_209/A gnd NAND2X1_748/Y vdd NAND2X1
XNAND2X1_759 BUFX4_142/Y NOR2X1_254/Y gnd NAND2X1_759/Y vdd NAND2X1
XFILL_0_7_1 gnd vdd FILL
XFILL_25_7_1 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XINVX8_7 INVX8_7/A gnd INVX8_7/Y vdd INVX8
XDFFPOSX1_60 NOR2X1_289/A CLKBUF1_2/Y AOI21X1_234/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 INVX1_385/A CLKBUF1_102/Y DFFPOSX1_71/D gnd vdd DFFPOSX1
XDFFPOSX1_93 NOR2X1_304/A CLKBUF1_42/Y DFFPOSX1_93/D gnd vdd DFFPOSX1
XDFFPOSX1_82 INVX1_66/A CLKBUF1_20/Y DFFPOSX1_82/D gnd vdd DFFPOSX1
XFILL_8_8_1 gnd vdd FILL
XBUFX4_16 clk gnd BUFX4_16/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XBUFX4_38 BUFX4_78/Y gnd BUFX4_38/Y vdd BUFX4
XBUFX4_49 BUFX4_50/A gnd BUFX4_49/Y vdd BUFX4
XBUFX4_27 a[0] gnd BUFX4_27/Y vdd BUFX4
XFILL_16_7_1 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XOAI21X1_528 BUFX4_372/Y NAND2X1_99/Y OAI21X1_528/C gnd OAI21X1_528/Y vdd OAI21X1
XOAI21X1_506 BUFX4_400/Y NAND2X1_97/Y OAI21X1_506/C gnd OAI21X1_506/Y vdd OAI21X1
XOAI21X1_539 BUFX4_150/Y NOR2X1_91/A NAND2X1_594/B gnd OAI21X1_539/Y vdd OAI21X1
XOAI21X1_517 NOR2X1_1/B NOR2X1_91/A INVX1_169/A gnd OAI21X1_517/Y vdd OAI21X1
XDFFPOSX1_431 OAI21X1_133/C CLKBUF1_49/Y OAI21X1_134/Y gnd vdd DFFPOSX1
XDFFPOSX1_420 INVX1_215/A CLKBUF1_82/Y OAI21X1_112/Y gnd vdd DFFPOSX1
XDFFPOSX1_464 NAND2X1_715/B CLKBUF1_87/Y OAI21X1_200/Y gnd vdd DFFPOSX1
XDFFPOSX1_453 INVX1_281/A CLKBUF1_18/Y OAI21X1_178/Y gnd vdd DFFPOSX1
XDFFPOSX1_442 NAND2X1_300/B CLKBUF1_41/Y OAI21X1_156/Y gnd vdd DFFPOSX1
XNAND2X1_501 BUFX4_212/Y NAND2X1_501/B gnd NAND2X1_501/Y vdd NAND2X1
XDFFPOSX1_475 NOR2X1_15/A CLKBUF1_56/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_497 INVX1_29/A CLKBUF1_30/Y OAI21X1_217/Y gnd vdd DFFPOSX1
XNAND2X1_512 AOI22X1_42/Y AOI22X1_43/Y gnd AOI22X1_44/D vdd NAND2X1
XDFFPOSX1_486 INVX1_347/A CLKBUF1_31/Y OAI21X1_214/Y gnd vdd DFFPOSX1
XNAND2X1_534 BUFX4_274/Y NAND2X1_534/B gnd NAND2X1_534/Y vdd NAND2X1
XNAND2X1_523 BUFX4_254/Y NAND2X1_523/B gnd NAND2X1_523/Y vdd NAND2X1
XNAND2X1_545 BUFX4_197/Y NOR2X1_235/A gnd NAND2X1_545/Y vdd NAND2X1
XNAND2X1_578 BUFX4_257/Y NOR2X1_18/A gnd NAND2X1_578/Y vdd NAND2X1
XNAND2X1_556 BUFX4_215/Y NAND2X1_556/B gnd NAND2X1_556/Y vdd NAND2X1
XNAND2X1_567 BUFX4_235/Y NOR2X1_375/A gnd NAND2X1_567/Y vdd NAND2X1
XNAND2X1_589 BUFX4_277/Y NAND2X1_589/B gnd NAND2X1_589/Y vdd NAND2X1
XFILL_40_5_1 gnd vdd FILL
XAOI21X1_191 BUFX4_398/Y NOR2X1_236/B NOR2X1_235/Y gnd AOI21X1_191/Y vdd AOI21X1
XAOI21X1_180 BUFX4_113/Y NOR2X1_222/B NOR2X1_222/Y gnd AOI21X1_180/Y vdd AOI21X1
XFILL_48_6_1 gnd vdd FILL
XFILL_47_1_0 gnd vdd FILL
XFILL_31_5_1 gnd vdd FILL
XFILL_30_0_0 gnd vdd FILL
XFILL_39_6_1 gnd vdd FILL
XFILL_38_1_0 gnd vdd FILL
XFILL_22_5_1 gnd vdd FILL
XOAI21X1_314 BUFX4_123/Y NAND2X1_77/Y OAI21X1_314/C gnd OAI21X1_314/Y vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_303 BUFX4_411/Y BUFX4_433/Y OAI21X1_303/C gnd OAI21X1_304/C vdd OAI21X1
XOAI21X1_325 BUFX4_404/Y BUFX4_381/Y INVX1_418/A gnd OAI21X1_326/C vdd OAI21X1
XOAI21X1_336 BUFX4_300/Y NAND2X1_78/Y OAI21X1_336/C gnd OAI21X1_336/Y vdd OAI21X1
XOAI21X1_347 BUFX4_307/Y INVX2_3/A INVX1_99/A gnd OAI21X1_347/Y vdd OAI21X1
XOAI21X1_369 NOR2X1_22/B BUFX4_386/Y NAND2X1_519/B gnd OAI21X1_369/Y vdd OAI21X1
XOAI21X1_358 BUFX4_284/Y NAND2X1_79/Y OAI21X1_357/Y gnd OAI21X1_358/Y vdd OAI21X1
XBUFX4_1 BUFX4_3/A gnd BUFX4_1/Y vdd BUFX4
XDFFPOSX1_250 NAND2X1_287/B CLKBUF1_35/Y DFFPOSX1_250/D gnd vdd DFFPOSX1
XDFFPOSX1_261 INVX1_269/A CLKBUF1_75/Y OAI21X1_1595/Y gnd vdd DFFPOSX1
XDFFPOSX1_272 NAND2X1_703/B CLKBUF1_27/Y OAI21X1_1617/Y gnd vdd DFFPOSX1
XDFFPOSX1_283 NOR2X1_362/A CLKBUF1_75/Y AOI21X1_288/Y gnd vdd DFFPOSX1
XNAND2X1_320 BUFX4_274/Y NOR2X1_94/A gnd NAND2X1_320/Y vdd NAND2X1
XDFFPOSX1_294 INVX1_335/A CLKBUF1_53/Y DFFPOSX1_294/D gnd vdd DFFPOSX1
XNAND2X1_342 BUFX4_213/Y NOR2X1_268/A gnd NAND2X1_342/Y vdd NAND2X1
XNAND2X1_353 BUFX4_235/Y NAND2X1_353/B gnd NAND2X1_353/Y vdd NAND2X1
XNAND2X1_331 BUFX4_195/Y OAI21X1_693/C gnd NAND2X1_331/Y vdd NAND2X1
XNAND2X1_375 BUFX4_275/Y OAI21X1_245/C gnd OAI21X1_945/C vdd NAND2X1
XFILL_5_6_1 gnd vdd FILL
XNAND2X1_364 BUFX4_255/Y OAI21X1_21/C gnd NAND2X1_364/Y vdd NAND2X1
XNAND2X1_386 INVX8_1/A OAI21X1_501/C gnd NAND2X1_386/Y vdd NAND2X1
XFILL_4_1_0 gnd vdd FILL
XFILL_29_1_0 gnd vdd FILL
XNAND2X1_397 BUFX4_218/Y NOR2X1_149/A gnd NAND2X1_397/Y vdd NAND2X1
XFILL_13_5_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XOAI21X1_881 INVX1_93/Y BUFX4_247/Y OAI21X1_881/C gnd MUX2X1_67/B vdd OAI21X1
XOAI21X1_870 INVX1_82/Y BUFX4_225/Y NAND2X1_294/Y gnd MUX2X1_58/A vdd OAI21X1
XOAI21X1_892 INVX1_104/Y BUFX4_269/Y NAND2X1_317/Y gnd MUX2X1_74/A vdd OAI21X1
XMUX2X1_370 MUX2X1_370/A MUX2X1_370/B BUFX4_48/Y gnd MUX2X1_372/B vdd MUX2X1
XNAND3X1_4 NAND3X1_4/A NAND3X1_4/B AOI22X1_5/Y gnd AOI22X1_6/D vdd NAND3X1
XOAI21X1_100 AOI21X1_6/A OAI21X1_96/B OAI21X1_99/Y gnd OAI21X1_100/Y vdd OAI21X1
XOAI21X1_122 BUFX4_127/Y NAND2X1_17/Y OAI21X1_122/C gnd OAI21X1_122/Y vdd OAI21X1
XOAI21X1_111 NOR2X1_91/B BUFX4_178/Y INVX1_215/A gnd OAI21X1_111/Y vdd OAI21X1
XAOI22X1_9 AOI22X1_9/A AOI22X1_9/B AOI22X1_9/C AOI22X1_9/D gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_155 NOR2X1_32/B BUFX4_175/Y NAND2X1_300/B gnd OAI21X1_156/C vdd OAI21X1
XOAI21X1_133 BUFX4_371/Y BUFX4_179/Y OAI21X1_133/C gnd OAI21X1_134/C vdd OAI21X1
XOAI21X1_144 NAND2X1_18/Y BUFX4_297/Y OAI21X1_144/C gnd OAI21X1_144/Y vdd OAI21X1
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XOAI21X1_188 BUFX4_423/Y NAND2X1_22/Y OAI21X1_187/Y gnd OAI21X1_188/Y vdd OAI21X1
XOAI21X1_177 BUFX4_457/Y BUFX4_134/Y INVX1_281/A gnd OAI21X1_178/C vdd OAI21X1
XOAI21X1_166 BUFX4_280/Y NAND2X1_19/Y OAI21X1_165/Y gnd OAI21X1_166/Y vdd OAI21X1
XOAI21X1_199 BUFX4_147/Y INVX1_1/A NAND2X1_715/B gnd OAI21X1_200/C vdd OAI21X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XNAND2X1_161 NAND2X1_9/A NOR2X1_155/Y gnd OAI21X1_663/C vdd NAND2X1
XNAND2X1_150 INVX8_10/A INVX1_4/Y gnd OAI21X1_635/B vdd NAND2X1
XNAND2X1_19 INVX8_16/A INVX2_1/Y gnd NAND2X1_19/Y vdd NAND2X1
XNAND2X1_183 BUFX4_452/Y NOR2X1_189/B gnd OAI21X1_714/C vdd NAND2X1
XNAND2X1_194 BUFX4_330/Y NOR2X1_199/Y gnd OAI21X1_725/C vdd NAND2X1
XNAND2X1_172 BUFX4_428/Y NOR2X1_166/Y gnd NAND2X1_172/Y vdd NAND2X1
XFILL_45_4_1 gnd vdd FILL
XAOI22X1_28 MUX2X1_135/Y INVX1_10/A INVX1_11/A MUX2X1_138/Y gnd AOI22X1_28/Y vdd AOI22X1
XAOI22X1_39 AOI22X1_39/A AOI22X1_9/D AOI22X1_69/C AOI22X1_39/D gnd AOI22X1_39/Y vdd
+ AOI22X1
XAOI22X1_17 MUX2X1_81/Y INVX1_6/A INVX1_8/A MUX2X1_84/Y gnd AOI22X1_17/Y vdd AOI22X1
XOAI21X1_1418 BUFX4_397/Y NAND2X1_814/Y OAI21X1_1417/Y gnd DFFPOSX1_133/D vdd OAI21X1
XOAI21X1_1407 BUFX4_416/Y BUFX4_466/Y NAND2X1_693/B gnd OAI21X1_1408/C vdd OAI21X1
XOAI21X1_1429 BUFX4_151/Y BUFX4_388/Y NAND2X1_349/B gnd OAI21X1_1429/Y vdd OAI21X1
XFILL_5_1 gnd vdd FILL
XFILL_47_1 gnd vdd FILL
XFILL_36_4_1 gnd vdd FILL
XFILL_2_4_1 gnd vdd FILL
XFILL_27_4_1 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XAOI21X1_50 BUFX4_424/Y NOR2X1_67/B NOR2X1_64/Y gnd AOI21X1_50/Y vdd AOI21X1
XAOI21X1_61 BUFX4_396/Y NOR2X1_77/B NOR2X1_77/Y gnd AOI21X1_61/Y vdd AOI21X1
XAOI21X1_83 AOI21X1_3/A NOR2X1_103/B NOR2X1_105/Y gnd AOI21X1_83/Y vdd AOI21X1
XAOI21X1_72 BUFX4_379/Y NOR2X1_90/B NOR2X1_90/Y gnd AOI21X1_72/Y vdd AOI21X1
XAOI21X1_94 BUFX4_396/Y NOR2X1_118/B AOI21X1_94/C gnd AOI21X1_94/Y vdd AOI21X1
XOAI21X1_1 NOR2X1_21/B OAI21X1_1/B INVX1_22/A gnd OAI21X1_2/C vdd OAI21X1
XFILL_9_0_0 gnd vdd FILL
XBUFX4_303 INVX8_5/Y gnd BUFX4_303/Y vdd BUFX4
XBUFX4_336 BUFX4_338/A gnd BUFX4_336/Y vdd BUFX4
XBUFX4_314 BUFX4_316/A gnd BUFX4_314/Y vdd BUFX4
XBUFX4_325 BUFX4_321/A gnd INVX1_10/A vdd BUFX4
XFILL_18_4_1 gnd vdd FILL
XBUFX4_358 a[2] gnd MUX2X1_42/S vdd BUFX4
XBUFX4_369 INVX8_15/Y gnd NOR2X1_52/B vdd BUFX4
XBUFX4_347 BUFX4_344/A gnd INVX2_10/A vdd BUFX4
XOAI21X1_1204 INVX1_416/Y BUFX4_200/Y NAND2X1_654/Y gnd MUX2X1_308/A vdd OAI21X1
XOAI21X1_1226 INVX1_438/Y BUFX4_244/Y NAND2X1_677/Y gnd MUX2X1_325/A vdd OAI21X1
XDFFPOSX1_805 INVX1_303/A CLKBUF1_2/Y OAI21X1_611/Y gnd vdd DFFPOSX1
XOAI21X1_1215 INVX1_427/Y BUFX4_222/Y NAND2X1_665/Y gnd MUX2X1_317/B vdd OAI21X1
XOAI21X1_1237 INVX1_449/Y BUFX4_266/Y NAND2X1_690/Y gnd MUX2X1_334/B vdd OAI21X1
XDFFPOSX1_838 INVX1_369/A CLKBUF1_81/Y OAI21X1_633/Y gnd vdd DFFPOSX1
XOAI21X1_1248 INVX1_460/Y BUFX4_189/Y NAND2X1_701/Y gnd MUX2X1_341/A vdd OAI21X1
XDFFPOSX1_827 NOR2X1_138/A CLKBUF1_85/Y AOI21X1_110/Y gnd vdd DFFPOSX1
XDFFPOSX1_816 NOR2X1_132/A CLKBUF1_33/Y AOI21X1_106/Y gnd vdd DFFPOSX1
XOAI21X1_1259 INVX1_471/Y BUFX4_211/Y NAND2X1_713/Y gnd MUX2X1_350/B vdd OAI21X1
XDFFPOSX1_849 MUX2X1_9/B CLKBUF1_7/Y AOI21X1_116/Y gnd vdd DFFPOSX1
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B MUX2X1_5/S gnd MUX2X1_5/Y vdd MUX2X1
XFILL_42_2_1 gnd vdd FILL
XCLKBUF1_6 BUFX4_10/Y gnd CLKBUF1_6/Y vdd CLKBUF1
XBUFX4_111 INVX8_4/Y gnd AOI21X1_3/A vdd BUFX4
XBUFX4_100 INVX8_7/Y gnd AOI21X1_6/A vdd BUFX4
XBUFX4_133 BUFX4_135/A gnd BUFX4_133/Y vdd BUFX4
XBUFX4_122 INVX8_2/Y gnd AOI21X1_1/A vdd BUFX4
XBUFX4_144 d[3] gnd BUFX4_144/Y vdd BUFX4
XBUFX4_155 BUFX4_155/A gnd BUFX4_155/Y vdd BUFX4
XNOR2X1_204 NOR2X1_204/A NOR2X1_206/B gnd NOR2X1_204/Y vdd NOR2X1
XBUFX4_188 BUFX4_26/Y gnd BUFX4_188/Y vdd BUFX4
XNOR2X1_215 NOR2X1_215/A NOR2X1_216/B gnd NOR2X1_215/Y vdd NOR2X1
XBUFX4_177 BUFX4_178/A gnd NOR2X1_2/A vdd BUFX4
XBUFX4_166 BUFX4_168/A gnd BUFX4_166/Y vdd BUFX4
XNOR2X1_248 INVX4_1/Y MUX2X1_30/Y gnd NOR2X1_248/Y vdd NOR2X1
XNOR2X1_226 NOR2X1_226/A NOR2X1_222/B gnd NOR2X1_226/Y vdd NOR2X1
XNOR2X1_237 NOR2X1_237/A NOR2X1_236/B gnd NOR2X1_237/Y vdd NOR2X1
XBUFX4_199 BUFX4_30/Y gnd BUFX4_199/Y vdd BUFX4
XNOR2X1_259 NOR2X1_259/A NOR2X1_256/B gnd NOR2X1_259/Y vdd NOR2X1
XFILL_33_2_1 gnd vdd FILL
XOAI21X1_1001 INVX1_213/Y BUFX4_190/Y NAND2X1_435/Y gnd MUX2X1_157/B vdd OAI21X1
XOAI21X1_1012 INVX1_224/Y BUFX4_212/Y NAND2X1_447/Y gnd MUX2X1_164/A vdd OAI21X1
XOAI21X1_1045 INVX1_257/Y BUFX4_278/Y NAND2X1_483/Y gnd MUX2X1_190/B vdd OAI21X1
XOAI21X1_1034 INVX1_246/Y BUFX4_256/Y NAND2X1_470/Y gnd MUX2X1_181/A vdd OAI21X1
XDFFPOSX1_613 INVX1_291/A CLKBUF1_60/Y OAI21X1_354/Y gnd vdd DFFPOSX1
XDFFPOSX1_602 NAND2X1_311/B CLKBUF1_97/Y OAI21X1_332/Y gnd vdd DFFPOSX1
XOAI21X1_1023 INVX1_235/Y BUFX4_234/Y NAND2X1_458/Y gnd MUX2X1_173/B vdd OAI21X1
XDFFPOSX1_635 OAI21X1_397/C CLKBUF1_10/Y OAI21X1_398/Y gnd vdd DFFPOSX1
XOAI21X1_1078 INVX1_290/Y BUFX4_245/Y NAND2X1_518/Y gnd MUX2X1_214/A vdd OAI21X1
XDFFPOSX1_624 OAI21X1_375/C CLKBUF1_60/Y OAI21X1_376/Y gnd vdd DFFPOSX1
XOAI21X1_1056 INVX1_268/Y BUFX4_201/Y NAND2X1_494/Y gnd MUX2X1_197/A vdd OAI21X1
XDFFPOSX1_657 INVX1_54/A CLKBUF1_58/Y OAI21X1_418/Y gnd vdd DFFPOSX1
XDFFPOSX1_646 INVX1_357/A CLKBUF1_33/Y OAI21X1_414/Y gnd vdd DFFPOSX1
XOAI21X1_1089 INVX1_301/Y BUFX4_267/Y NAND2X1_530/Y gnd MUX2X1_223/B vdd OAI21X1
XOAI21X1_1067 INVX1_279/Y BUFX4_223/Y NAND2X1_506/Y gnd MUX2X1_206/B vdd OAI21X1
XDFFPOSX1_668 OAI21X1_439/C CLKBUF1_58/Y OAI21X1_440/Y gnd vdd DFFPOSX1
XDFFPOSX1_679 INVX1_423/A CLKBUF1_38/Y OAI21X1_462/Y gnd vdd DFFPOSX1
XINVX1_380 INVX1_380/A gnd INVX1_380/Y vdd INVX1
XNAND2X1_727 BUFX4_236/Y OAI21X1_407/C gnd NAND2X1_727/Y vdd NAND2X1
XNAND2X1_716 BUFX4_216/Y NOR2X1_20/A gnd NAND2X1_716/Y vdd NAND2X1
XINVX1_391 INVX1_391/A gnd INVX1_391/Y vdd INVX1
XNAND2X1_705 BUFX4_194/Y NOR2X1_377/A gnd NAND2X1_705/Y vdd NAND2X1
XNAND2X1_749 BUFX4_278/Y NAND2X1_749/B gnd NAND2X1_749/Y vdd NAND2X1
XNAND2X1_738 BUFX4_256/Y NOR2X1_121/A gnd NAND2X1_738/Y vdd NAND2X1
XFILL_24_2_1 gnd vdd FILL
XINVX8_8 INVX8_8/A gnd INVX8_8/Y vdd INVX8
XDFFPOSX1_72 INVX1_449/A CLKBUF1_43/Y DFFPOSX1_72/D gnd vdd DFFPOSX1
XDFFPOSX1_50 INVX1_64/A CLKBUF1_56/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XDFFPOSX1_61 NOR2X1_290/A CLKBUF1_37/Y DFFPOSX1_61/D gnd vdd DFFPOSX1
XDFFPOSX1_83 INVX1_130/A CLKBUF1_78/Y DFFPOSX1_83/D gnd vdd DFFPOSX1
XOAI21X1_1590 BUFX4_454/Y INVX2_10/A INVX1_141/A gnd OAI21X1_1591/C vdd OAI21X1
XDFFPOSX1_94 NOR2X1_305/A CLKBUF1_25/Y DFFPOSX1_94/D gnd vdd DFFPOSX1
XBUFX4_17 clk gnd BUFX4_17/Y vdd BUFX4
XFILL_7_3_1 gnd vdd FILL
XBUFX4_39 BUFX4_78/Y gnd BUFX4_39/Y vdd BUFX4
XBUFX4_28 a[0] gnd BUFX4_28/Y vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XOAI21X1_507 BUFX4_414/Y BUFX4_340/Y NAND2X1_593/B gnd OAI21X1_507/Y vdd OAI21X1
XOAI21X1_518 BUFX4_116/Y NAND2X1_99/Y OAI21X1_517/Y gnd OAI21X1_518/Y vdd OAI21X1
XOAI21X1_529 BUFX4_153/Y BUFX4_293/Y NAND2X1_267/B gnd OAI21X1_529/Y vdd OAI21X1
XDFFPOSX1_410 OAI21X1_91/C CLKBUF1_72/Y OAI21X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_421 INVX1_279/A CLKBUF1_48/Y OAI21X1_114/Y gnd vdd DFFPOSX1
XDFFPOSX1_454 INVX1_345/A CLKBUF1_50/Y OAI21X1_180/Y gnd vdd DFFPOSX1
XDFFPOSX1_465 INVX1_31/A CLKBUF1_71/Y OAI21X1_201/Y gnd vdd DFFPOSX1
XDFFPOSX1_432 NAND2X1_713/B CLKBUF1_77/Y OAI21X1_136/Y gnd vdd DFFPOSX1
XDFFPOSX1_443 OAI21X1_157/C CLKBUF1_11/Y OAI21X1_158/Y gnd vdd DFFPOSX1
XDFFPOSX1_498 INVX1_92/A CLKBUF1_24/Y OAI21X1_218/Y gnd vdd DFFPOSX1
XNAND2X1_502 BUFX4_214/Y OAI21X1_25/C gnd NAND2X1_502/Y vdd NAND2X1
XDFFPOSX1_476 NOR2X1_16/A CLKBUF1_56/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_487 INVX1_411/A CLKBUF1_2/Y OAI21X1_215/Y gnd vdd DFFPOSX1
XNAND2X1_535 BUFX4_276/Y NOR2X1_151/A gnd NAND2X1_535/Y vdd NAND2X1
XNAND2X1_513 BUFX4_234/Y NAND2X1_513/B gnd NAND2X1_513/Y vdd NAND2X1
XNAND2X1_524 BUFX4_256/Y NAND2X1_524/B gnd NAND2X1_524/Y vdd NAND2X1
XNAND2X1_546 AOI22X1_47/Y AOI22X1_48/Y gnd AOI22X1_49/D vdd NAND2X1
XNAND2X1_579 BUFX4_259/Y NOR2X1_28/A gnd NAND2X1_579/Y vdd NAND2X1
XNAND2X1_557 BUFX4_217/Y NOR2X1_328/A gnd NAND2X1_557/Y vdd NAND2X1
XNAND2X1_568 BUFX4_237/Y NAND2X1_568/B gnd NAND2X1_568/Y vdd NAND2X1
XAOI21X1_181 BUFX4_302/Y NOR2X1_222/B NOR2X1_223/Y gnd AOI21X1_181/Y vdd AOI21X1
XAOI21X1_192 BUFX4_102/Y NOR2X1_236/B NOR2X1_236/Y gnd AOI21X1_192/Y vdd AOI21X1
XAOI21X1_170 BUFX4_130/Y NOR2X1_216/B NOR2X1_211/Y gnd AOI21X1_170/Y vdd AOI21X1
XFILL_47_1_1 gnd vdd FILL
XFILL_30_0_1 gnd vdd FILL
XFILL_38_1_1 gnd vdd FILL
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_304 BUFX4_379/Y NAND2X1_67/Y OAI21X1_304/C gnd OAI21X1_304/Y vdd OAI21X1
XOAI21X1_315 BUFX4_403/Y BUFX4_381/Y INVX1_98/A gnd OAI21X1_316/C vdd OAI21X1
XOAI21X1_326 BUFX4_284/Y NAND2X1_77/Y OAI21X1_326/C gnd OAI21X1_326/Y vdd OAI21X1
XOAI21X1_337 BUFX4_85/Y INVX2_3/A NAND2X1_518/B gnd OAI21X1_338/C vdd OAI21X1
XOAI21X1_348 BUFX4_421/Y NAND2X1_79/Y OAI21X1_347/Y gnd OAI21X1_348/Y vdd OAI21X1
XOAI21X1_359 BUFX4_310/Y INVX2_3/A INVX1_483/A gnd OAI21X1_360/C vdd OAI21X1
XDFFPOSX1_240 NOR2X1_357/A CLKBUF1_64/Y AOI21X1_285/Y gnd vdd DFFPOSX1
XBUFX4_2 BUFX4_3/A gnd BUFX4_2/Y vdd BUFX4
XDFFPOSX1_251 NAND2X1_356/B CLKBUF1_76/Y OAI21X1_1575/Y gnd vdd DFFPOSX1
XDFFPOSX1_273 INVX1_19/A CLKBUF1_31/Y OAI21X1_1618/Y gnd vdd DFFPOSX1
XDFFPOSX1_262 INVX1_333/A CLKBUF1_75/Y OAI21X1_1597/Y gnd vdd DFFPOSX1
XNAND2X1_310 BUFX4_254/Y NOR2X1_64/A gnd NAND2X1_310/Y vdd NAND2X1
XDFFPOSX1_284 NOR2X1_363/A CLKBUF1_94/Y AOI21X1_289/Y gnd vdd DFFPOSX1
XDFFPOSX1_295 INVX1_399/A CLKBUF1_68/Y DFFPOSX1_295/D gnd vdd DFFPOSX1
XNAND2X1_332 BUFX4_197/Y NOR2X1_181/A gnd OAI21X1_906/C vdd NAND2X1
XNAND2X1_354 BUFX4_237/Y NOR2X1_344/A gnd NAND2X1_354/Y vdd NAND2X1
XNAND2X1_343 BUFX4_215/Y NOR2X1_278/A gnd NAND2X1_343/Y vdd NAND2X1
XNAND2X1_321 BUFX4_276/Y NOR2X1_104/A gnd OAI21X1_896/C vdd NAND2X1
XNAND2X1_365 BUFX4_257/Y OAI21X1_53/C gnd NAND2X1_365/Y vdd NAND2X1
XNAND2X1_387 BUFX4_200/Y NAND2X1_387/B gnd OAI21X1_957/C vdd NAND2X1
XNAND2X1_376 BUFX4_277/Y NOR2X1_45/A gnd OAI21X1_946/C vdd NAND2X1
XNAND2X1_398 BUFX4_220/Y NOR2X1_160/A gnd OAI21X1_967/C vdd NAND2X1
XFILL_4_1_1 gnd vdd FILL
XFILL_29_1_1 gnd vdd FILL
XFILL_41_8_0 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XINVX4_2 we gnd INVX4_2/Y vdd INVX4
XOAI21X1_860 INVX1_72/Y BUFX4_205/Y OAI21X1_860/C gnd MUX2X1_50/A vdd OAI21X1
XOAI21X1_882 INVX1_94/Y BUFX4_249/Y OAI21X1_882/C gnd MUX2X1_67/A vdd OAI21X1
XOAI21X1_871 INVX1_83/Y BUFX4_227/Y NAND2X1_295/Y gnd MUX2X1_59/B vdd OAI21X1
XOAI21X1_893 INVX1_105/Y BUFX4_271/Y OAI21X1_893/C gnd MUX2X1_76/B vdd OAI21X1
XMUX2X1_360 MUX2X1_359/Y MUX2X1_358/Y MUX2X1_96/S gnd MUX2X1_360/Y vdd MUX2X1
XMUX2X1_371 MUX2X1_371/A MUX2X1_371/B BUFX4_1/Y gnd MUX2X1_372/A vdd MUX2X1
XFILL_32_8_0 gnd vdd FILL
XNAND3X1_5 NAND3X1_5/A NAND3X1_5/B NAND3X1_5/C gnd AOI22X1_9/B vdd NAND3X1
XFILL_23_8_0 gnd vdd FILL
XOAI21X1_101 BUFX4_84/Y BUFX4_179/Y NAND2X1_643/B gnd OAI21X1_102/C vdd OAI21X1
XOAI21X1_112 BUFX4_297/Y NAND2X1_16/Y OAI21X1_111/Y gnd OAI21X1_112/Y vdd OAI21X1
XOAI21X1_156 BUFX4_425/Y NAND2X1_19/Y OAI21X1_156/C gnd OAI21X1_156/Y vdd OAI21X1
XOAI21X1_134 BUFX4_280/Y NAND2X1_17/Y OAI21X1_134/C gnd OAI21X1_134/Y vdd OAI21X1
XOAI21X1_123 BUFX4_371/Y BUFX4_175/Y NAND2X1_299/B gnd OAI21X1_123/Y vdd OAI21X1
XOAI21X1_145 INVX4_3/A BUFX4_173/Y INVX1_280/A gnd OAI21X1_145/Y vdd OAI21X1
XOAI21X1_189 BUFX4_147/Y BUFX4_133/Y OAI21X1_189/C gnd OAI21X1_190/C vdd OAI21X1
XOAI21X1_178 BUFX4_395/Y NAND2X1_21/Y OAI21X1_178/C gnd OAI21X1_178/Y vdd OAI21X1
XOAI21X1_167 NOR2X1_32/B INVX2_1/A NAND2X1_714/B gnd OAI21X1_168/C vdd OAI21X1
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XNAND2X1_140 INVX8_8/A NOR2X1_122/Y gnd OAI21X1_613/C vdd NAND2X1
XNAND2X1_151 INVX8_11/A INVX1_4/Y gnd OAI21X1_651/B vdd NAND2X1
XNAND2X1_162 BUFX4_444/Y NOR2X1_155/Y gnd NAND2X1_162/Y vdd NAND2X1
XNAND2X1_184 BUFX4_334/Y NOR2X1_189/B gnd OAI21X1_715/C vdd NAND2X1
XNAND2X1_195 BUFX4_140/Y NOR2X1_199/Y gnd OAI21X1_726/C vdd NAND2X1
XNAND2X1_173 INVX1_10/A AOI22X1_69/C gnd BUFX4_64/A vdd NAND2X1
XFILL_14_8_0 gnd vdd FILL
XAOI22X1_18 MUX2X1_87/Y BUFX4_324/Y BUFX4_290/Y MUX2X1_90/Y gnd AOI22X1_18/Y vdd AOI22X1
XAOI22X1_29 AOI22X1_29/A AOI22X1_9/D AOI22X1_69/C AOI22X1_29/D gnd AOI22X1_29/Y vdd
+ AOI22X1
XOAI21X1_1419 BUFX4_457/Y BUFX4_389/Y INVX1_325/A gnd OAI21X1_1420/C vdd OAI21X1
XOAI21X1_1408 BUFX4_376/Y NAND2X1_812/Y OAI21X1_1408/C gnd OAI21X1_1408/Y vdd OAI21X1
XOAI21X1_690 BUFX4_375/Y NAND2X1_174/Y OAI21X1_690/C gnd OAI21X1_690/Y vdd OAI21X1
XMUX2X1_190 MUX2X1_190/A MUX2X1_190/B BUFX4_48/Y gnd MUX2X1_192/B vdd MUX2X1
XFILL_47_2 gnd vdd FILL
XAOI21X1_51 BUFX4_113/Y NOR2X1_67/B NOR2X1_65/Y gnd AOI21X1_51/Y vdd AOI21X1
XAOI21X1_62 BUFX4_103/Y NOR2X1_77/B NOR2X1_78/Y gnd AOI21X1_62/Y vdd AOI21X1
XAOI21X1_40 BUFX4_379/Y NOR2X1_43/B NOR2X1_50/Y gnd AOI21X1_40/Y vdd AOI21X1
XAOI21X1_95 BUFX4_104/Y NOR2X1_118/B AOI21X1_95/C gnd AOI21X1_95/Y vdd AOI21X1
XAOI21X1_84 BUFX4_298/Y NOR2X1_103/B AOI21X1_84/C gnd AOI21X1_84/Y vdd AOI21X1
XAOI21X1_73 BUFX4_129/Y NOR2X1_96/B NOR2X1_93/Y gnd AOI21X1_73/Y vdd AOI21X1
XOAI21X1_2 BUFX4_128/Y NAND2X1_1/Y OAI21X1_2/C gnd OAI21X1_2/Y vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XBUFX4_304 INVX8_5/Y gnd BUFX4_304/Y vdd BUFX4
XBUFX4_337 BUFX4_338/A gnd BUFX4_337/Y vdd BUFX4
XBUFX4_315 BUFX4_316/A gnd OAI21X1_5/B vdd BUFX4
XBUFX4_326 d[5] gnd BUFX4_326/Y vdd BUFX4
XFILL_46_7_0 gnd vdd FILL
XBUFX4_359 a[2] gnd INVX2_6/A vdd BUFX4
XBUFX4_348 BUFX4_344/A gnd BUFX4_348/Y vdd BUFX4
XOAI21X1_1227 INVX1_439/Y BUFX4_246/Y NAND2X1_678/Y gnd MUX2X1_326/B vdd OAI21X1
XOAI21X1_1205 INVX1_417/Y BUFX4_202/Y NAND2X1_655/Y gnd MUX2X1_310/B vdd OAI21X1
XDFFPOSX1_806 INVX1_367/A CLKBUF1_30/Y OAI21X1_612/Y gnd vdd DFFPOSX1
XOAI21X1_1216 INVX1_428/Y BUFX4_224/Y NAND2X1_666/Y gnd MUX2X1_317/A vdd OAI21X1
XOAI21X1_1238 INVX1_450/Y BUFX4_268/Y NAND2X1_691/Y gnd MUX2X1_334/A vdd OAI21X1
XDFFPOSX1_839 INVX1_433/A CLKBUF1_15/Y OAI21X1_635/Y gnd vdd DFFPOSX1
XDFFPOSX1_817 MUX2X1_5/B CLKBUF1_96/Y AOI21X1_107/Y gnd vdd DFFPOSX1
XDFFPOSX1_828 NOR2X1_139/A CLKBUF1_24/Y AOI21X1_111/Y gnd vdd DFFPOSX1
XOAI21X1_1249 INVX1_461/Y BUFX4_191/Y NAND2X1_703/Y gnd MUX2X1_343/B vdd OAI21X1
XFILL_37_7_0 gnd vdd FILL
XFILL_20_6_0 gnd vdd FILL
XFILL_3_7_0 gnd vdd FILL
XFILL_28_7_0 gnd vdd FILL
XMUX2X1_6 MUX2X1_5/Y MUX2X1_6/B BUFX4_56/Y gnd MUX2X1_6/Y vdd MUX2X1
XFILL_11_6_0 gnd vdd FILL
XCLKBUF1_7 BUFX4_18/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XBUFX4_101 INVX8_7/Y gnd BUFX4_101/Y vdd BUFX4
XBUFX4_112 INVX8_4/Y gnd BUFX4_112/Y vdd BUFX4
XBUFX4_123 INVX8_2/Y gnd BUFX4_123/Y vdd BUFX4
XBUFX4_134 BUFX4_135/A gnd BUFX4_134/Y vdd BUFX4
XFILL_19_7_0 gnd vdd FILL
XBUFX4_145 d[3] gnd BUFX4_145/Y vdd BUFX4
XBUFX4_167 BUFX4_168/A gnd BUFX4_167/Y vdd BUFX4
XNOR2X1_205 NOR2X1_205/A NOR2X1_206/B gnd NOR2X1_205/Y vdd NOR2X1
XBUFX4_156 BUFX4_155/A gnd BUFX4_156/Y vdd BUFX4
XNOR2X1_216 NOR2X1_216/A NOR2X1_216/B gnd NOR2X1_216/Y vdd NOR2X1
XBUFX4_178 BUFX4_178/A gnd BUFX4_178/Y vdd BUFX4
XNOR2X1_227 NOR2X1_227/A NOR2X1_222/B gnd NOR2X1_227/Y vdd NOR2X1
XNOR2X1_238 NOR2X1_238/A NOR2X1_236/B gnd NOR2X1_238/Y vdd NOR2X1
XBUFX4_189 BUFX4_26/Y gnd BUFX4_189/Y vdd BUFX4
XNOR2X1_249 a[6] a[5] gnd AOI22X1_9/A vdd NOR2X1
XOAI21X1_1013 INVX1_225/Y BUFX4_214/Y NAND2X1_448/Y gnd MUX2X1_166/B vdd OAI21X1
XOAI21X1_1002 INVX1_214/Y BUFX4_192/Y NAND2X1_436/Y gnd MUX2X1_157/A vdd OAI21X1
XOAI21X1_1046 INVX1_258/Y MUX2X1_2/S NAND2X1_484/Y gnd MUX2X1_190/A vdd OAI21X1
XDFFPOSX1_603 OAI21X1_333/C CLKBUF1_47/Y OAI21X1_334/Y gnd vdd DFFPOSX1
XDFFPOSX1_614 INVX1_355/A CLKBUF1_28/Y OAI21X1_356/Y gnd vdd DFFPOSX1
XOAI21X1_1035 INVX1_247/Y BUFX4_258/Y NAND2X1_471/Y gnd MUX2X1_182/B vdd OAI21X1
XOAI21X1_1024 INVX1_236/Y BUFX4_236/Y NAND2X1_459/Y gnd MUX2X1_173/A vdd OAI21X1
XDFFPOSX1_625 INVX1_52/A CLKBUF1_60/Y OAI21X1_378/Y gnd vdd DFFPOSX1
XDFFPOSX1_636 NAND2X1_451/B CLKBUF1_22/Y OAI21X1_400/Y gnd vdd DFFPOSX1
XOAI21X1_1079 INVX1_291/Y BUFX4_247/Y NAND2X1_519/Y gnd MUX2X1_215/B vdd OAI21X1
XDFFPOSX1_647 INVX1_421/A CLKBUF1_33/Y OAI21X1_415/Y gnd vdd DFFPOSX1
XOAI21X1_1057 INVX1_269/Y BUFX4_203/Y NAND2X1_496/Y gnd MUX2X1_199/B vdd OAI21X1
XOAI21X1_1068 INVX1_280/Y BUFX4_225/Y NAND2X1_507/Y gnd MUX2X1_206/A vdd OAI21X1
XDFFPOSX1_669 NAND2X1_522/B CLKBUF1_70/Y OAI21X1_442/Y gnd vdd DFFPOSX1
XDFFPOSX1_658 INVX1_102/A CLKBUF1_85/Y OAI21X1_420/Y gnd vdd DFFPOSX1
XINVX1_370 INVX1_370/A gnd INVX1_370/Y vdd INVX1
XINVX1_392 INVX1_392/A gnd INVX1_392/Y vdd INVX1
XINVX1_381 INVX1_381/A gnd INVX1_381/Y vdd INVX1
XNAND2X1_728 BUFX4_238/Y NOR2X1_80/A gnd NAND2X1_728/Y vdd NAND2X1
XNAND2X1_717 BUFX4_218/Y NOR2X1_30/A gnd NAND2X1_717/Y vdd NAND2X1
XNAND2X1_706 BUFX4_196/Y NAND2X1_706/B gnd NAND2X1_706/Y vdd NAND2X1
XNAND2X1_739 BUFX4_258/Y NOR2X1_132/A gnd NAND2X1_739/Y vdd NAND2X1
XINVX8_9 INVX8_9/A gnd INVX8_9/Y vdd INVX8
XDFFPOSX1_62 NOR2X1_291/A CLKBUF1_3/Y DFFPOSX1_62/D gnd vdd DFFPOSX1
XDFFPOSX1_40 INVX1_447/A CLKBUF1_56/Y DFFPOSX1_40/D gnd vdd DFFPOSX1
XDFFPOSX1_51 INVX1_128/A CLKBUF1_2/Y DFFPOSX1_51/D gnd vdd DFFPOSX1
XDFFPOSX1_84 INVX1_194/A CLKBUF1_78/Y DFFPOSX1_84/D gnd vdd DFFPOSX1
XDFFPOSX1_73 DFFPOSX1_73/Q CLKBUF1_42/Y DFFPOSX1_73/D gnd vdd DFFPOSX1
XOAI21X1_1580 BUFX4_410/Y BUFX4_95/Y NAND2X1_563/B gnd OAI21X1_1581/C vdd OAI21X1
XOAI21X1_1591 BUFX4_114/Y NAND2X1_842/Y OAI21X1_1591/C gnd OAI21X1_1591/Y vdd OAI21X1
XDFFPOSX1_95 NOR2X1_306/A CLKBUF1_20/Y DFFPOSX1_95/D gnd vdd DFFPOSX1
XBUFX4_18 clk gnd BUFX4_18/Y vdd BUFX4
XBUFX4_29 a[0] gnd BUFX4_29/Y vdd BUFX4
XFILL_43_5_0 gnd vdd FILL
XFILL_34_5_0 gnd vdd FILL
XFILL_22_1 gnd vdd FILL
XOAI21X1_508 BUFX4_101/Y NAND2X1_97/Y OAI21X1_507/Y gnd OAI21X1_508/Y vdd OAI21X1
XOAI21X1_519 BUFX4_461/Y INVX1_2/A INVX1_233/A gnd OAI21X1_520/C vdd OAI21X1
XDFFPOSX1_400 NOR2X1_10/A CLKBUF1_72/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_411 OAI21X1_93/C CLKBUF1_72/Y OAI21X1_94/Y gnd vdd DFFPOSX1
XDFFPOSX1_422 INVX1_343/A CLKBUF1_77/Y OAI21X1_116/Y gnd vdd DFFPOSX1
XDFFPOSX1_455 INVX1_409/A CLKBUF1_50/Y OAI21X1_182/Y gnd vdd DFFPOSX1
XDFFPOSX1_433 INVX1_25/A CLKBUF1_48/Y OAI21X1_138/Y gnd vdd DFFPOSX1
XDFFPOSX1_444 OAI21X1_159/C CLKBUF1_82/Y OAI21X1_160/Y gnd vdd DFFPOSX1
XNAND2X1_503 BUFX4_216/Y OAI21X1_57/C gnd NAND2X1_503/Y vdd NAND2X1
XDFFPOSX1_477 NOR2X1_17/A CLKBUF1_23/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_466 INVX1_90/A CLKBUF1_71/Y OAI21X1_202/Y gnd vdd DFFPOSX1
XDFFPOSX1_488 INVX1_475/A CLKBUF1_89/Y OAI21X1_216/Y gnd vdd DFFPOSX1
XDFFPOSX1_499 INVX1_156/A CLKBUF1_24/Y OAI21X1_219/Y gnd vdd DFFPOSX1
XNAND2X1_536 BUFX4_278/Y NOR2X1_162/A gnd NAND2X1_536/Y vdd NAND2X1
XNAND2X1_514 BUFX4_236/Y NOR2X1_47/A gnd NAND2X1_514/Y vdd NAND2X1
XNAND2X1_525 BUFX4_258/Y NAND2X1_525/B gnd NAND2X1_525/Y vdd NAND2X1
XNAND2X1_569 BUFX4_239/Y NOR2X1_385/A gnd NAND2X1_569/Y vdd NAND2X1
XNAND2X1_547 AOI22X1_44/Y AOI22X1_49/Y gnd NAND2X1_547/Y vdd NAND2X1
XNAND2X1_558 BUFX4_219/Y NOR2X1_338/A gnd NAND2X1_558/Y vdd NAND2X1
XFILL_0_5_0 gnd vdd FILL
XFILL_25_5_0 gnd vdd FILL
XAOI21X1_160 BUFX4_375/Y NOR2X1_197/B NOR2X1_198/Y gnd AOI21X1_160/Y vdd AOI21X1
XAOI21X1_193 BUFX4_283/Y NOR2X1_236/B NOR2X1_237/Y gnd AOI21X1_193/Y vdd AOI21X1
XAOI21X1_182 BUFX4_400/Y NOR2X1_222/B NOR2X1_224/Y gnd AOI21X1_182/Y vdd AOI21X1
XAOI21X1_171 BUFX4_425/Y NOR2X1_216/B NOR2X1_212/Y gnd AOI21X1_171/Y vdd AOI21X1
XFILL_8_6_0 gnd vdd FILL
XFILL_16_5_0 gnd vdd FILL
XOAI21X1_305 INVX1_49/Y NOR2X1_61/Y NAND2X1_69/Y gnd OAI21X1_305/Y vdd OAI21X1
XOAI21X1_327 BUFX4_403/Y BUFX4_381/Y INVX1_482/A gnd OAI21X1_327/Y vdd OAI21X1
XOAI21X1_316 BUFX4_421/Y NAND2X1_77/Y OAI21X1_316/C gnd OAI21X1_316/Y vdd OAI21X1
XOAI21X1_338 BUFX4_401/Y NAND2X1_78/Y OAI21X1_338/C gnd OAI21X1_338/Y vdd OAI21X1
XOAI21X1_349 BUFX4_307/Y BUFX4_387/Y INVX1_163/A gnd OAI21X1_350/C vdd OAI21X1
XDFFPOSX1_230 INVX1_331/A CLKBUF1_52/Y DFFPOSX1_230/D gnd vdd DFFPOSX1
XBUFX4_3 BUFX4_3/A gnd BUFX4_3/Y vdd BUFX4
XDFFPOSX1_241 NAND2X1_211/A CLKBUF1_66/Y DFFPOSX1_241/D gnd vdd DFFPOSX1
XDFFPOSX1_252 NAND2X1_425/B CLKBUF1_52/Y DFFPOSX1_252/D gnd vdd DFFPOSX1
XDFFPOSX1_263 INVX1_397/A CLKBUF1_12/Y OAI21X1_1599/Y gnd vdd DFFPOSX1
XNAND2X1_311 BUFX4_256/Y NAND2X1_311/B gnd NAND2X1_311/Y vdd NAND2X1
XDFFPOSX1_274 INVX1_78/A CLKBUF1_89/Y OAI21X1_1619/Y gnd vdd DFFPOSX1
XDFFPOSX1_285 NOR2X1_364/A CLKBUF1_12/Y AOI21X1_290/Y gnd vdd DFFPOSX1
XNAND2X1_300 BUFX4_236/Y NAND2X1_300/B gnd NAND2X1_300/Y vdd NAND2X1
XDFFPOSX1_296 INVX1_463/A CLKBUF1_39/Y OAI21X1_1633/Y gnd vdd DFFPOSX1
XNAND2X1_333 BUFX4_199/Y NOR2X1_192/A gnd NAND2X1_333/Y vdd NAND2X1
XNAND2X1_344 BUFX4_217/Y NOR2X1_288/A gnd OAI21X1_916/C vdd NAND2X1
XNAND2X1_322 AOI22X1_15/Y AOI22X1_16/Y gnd AOI22X1_19/A vdd NAND2X1
XNAND2X1_377 MUX2X1_1/S NOR2X1_55/A gnd OAI21X1_947/C vdd NAND2X1
XNAND2X1_355 BUFX4_239/Y NOR2X1_352/A gnd NAND2X1_355/Y vdd NAND2X1
XNAND2X1_366 BUFX4_259/Y NOR2X1_5/A gnd OAI21X1_937/C vdd NAND2X1
XNAND2X1_399 BUFX4_222/Y NOR2X1_171/A gnd OAI21X1_968/C vdd NAND2X1
XNAND2X1_388 BUFX4_202/Y NOR2X1_85/A gnd NAND2X1_388/Y vdd NAND2X1
XFILL_41_8_1 gnd vdd FILL
XFILL_40_3_0 gnd vdd FILL
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XOAI21X1_850 INVX1_62/Y MUX2X1_9/S OAI21X1_850/C gnd MUX2X1_43/A vdd OAI21X1
XOAI21X1_883 INVX1_95/Y BUFX4_251/Y OAI21X1_883/C gnd MUX2X1_68/B vdd OAI21X1
XOAI21X1_861 INVX1_73/Y BUFX4_207/Y OAI21X1_861/C gnd MUX2X1_52/B vdd OAI21X1
XOAI21X1_872 INVX1_84/Y BUFX4_229/Y NAND2X1_296/Y gnd MUX2X1_59/A vdd OAI21X1
XOAI21X1_894 INVX1_106/Y BUFX4_273/Y NAND2X1_319/Y gnd MUX2X1_76/A vdd OAI21X1
XMUX2X1_350 MUX2X1_350/A MUX2X1_350/B BUFX4_35/Y gnd MUX2X1_351/A vdd MUX2X1
XMUX2X1_361 MUX2X1_361/A MUX2X1_361/B BUFX4_82/Y gnd MUX2X1_361/Y vdd MUX2X1
XMUX2X1_372 MUX2X1_372/A MUX2X1_372/B MUX2X1_42/S gnd AOI22X1_77/D vdd MUX2X1
XFILL_48_4_0 gnd vdd FILL
XFILL_32_8_1 gnd vdd FILL
XFILL_31_3_0 gnd vdd FILL
XNAND3X1_6 NAND3X1_6/A NAND3X1_6/B AOI22X1_9/Y gnd NAND3X1_6/Y vdd NAND3X1
XFILL_39_4_0 gnd vdd FILL
XFILL_23_8_1 gnd vdd FILL
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_102 BUFX4_280/Y OAI21X1_96/B OAI21X1_102/C gnd OAI21X1_102/Y vdd OAI21X1
XOAI21X1_113 NOR2X1_51/B BUFX4_179/Y INVX1_279/A gnd OAI21X1_114/C vdd OAI21X1
XOAI21X1_135 NOR2X1_52/B NOR2X1_1/A NAND2X1_713/B gnd OAI21X1_135/Y vdd OAI21X1
XOAI21X1_124 BUFX4_422/Y NAND2X1_17/Y OAI21X1_123/Y gnd OAI21X1_124/Y vdd OAI21X1
XOAI21X1_146 NAND2X1_18/Y BUFX4_394/Y OAI21X1_145/Y gnd OAI21X1_146/Y vdd OAI21X1
XOAI21X1_179 BUFX4_457/Y BUFX4_134/Y INVX1_345/A gnd OAI21X1_180/C vdd OAI21X1
XOAI21X1_168 BUFX4_374/Y NAND2X1_19/Y OAI21X1_168/C gnd OAI21X1_168/Y vdd OAI21X1
XOAI21X1_157 BUFX4_412/Y BUFX4_173/Y OAI21X1_157/C gnd OAI21X1_158/C vdd OAI21X1
XNAND2X1_141 INVX8_9/A NOR2X1_122/Y gnd OAI21X1_614/C vdd NAND2X1
XNAND2X1_130 BUFX4_142/Y NOR2X1_111/Y gnd OAI21X1_603/C vdd NAND2X1
XNAND2X1_152 BUFX4_453/Y NOR2X1_145/B gnd OAI21X1_654/C vdd NAND2X1
XNAND2X1_174 INVX8_10/A INVX1_5/Y gnd NAND2X1_174/Y vdd NAND2X1
XFILL_5_4_0 gnd vdd FILL
XNAND2X1_185 BUFX4_144/Y NOR2X1_189/B gnd OAI21X1_716/C vdd NAND2X1
XNAND2X1_196 BUFX4_431/Y NOR2X1_199/Y gnd OAI21X1_727/C vdd NAND2X1
XNAND2X1_163 BUFX4_326/Y NOR2X1_155/Y gnd OAI21X1_665/C vdd NAND2X1
XFILL_14_8_1 gnd vdd FILL
XFILL_13_3_0 gnd vdd FILL
XAOI22X1_19 AOI22X1_19/A AOI22X1_9/D AOI22X1_69/C AOI22X1_19/D gnd AOI22X1_19/Y vdd
+ AOI22X1
XOAI21X1_1409 BUFX4_460/Y BUFX4_388/Y INVX1_41/A gnd OAI21X1_1409/Y vdd OAI21X1
XOAI21X1_691 BUFX4_146/Y BUFX4_66/Y MUX2X1_15/A gnd OAI21X1_692/C vdd OAI21X1
XOAI21X1_680 BUFX4_115/Y NAND2X1_174/Y OAI21X1_679/Y gnd OAI21X1_680/Y vdd OAI21X1
XMUX2X1_180 MUX2X1_180/A MUX2X1_180/B MUX2X1_48/S gnd AOI22X1_37/D vdd MUX2X1
XMUX2X1_191 MUX2X1_191/A MUX2X1_191/B BUFX4_1/Y gnd MUX2X1_191/Y vdd MUX2X1
XAOI21X1_41 BUFX4_129/Y NOR2X1_55/B NOR2X1_53/Y gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_52 BUFX4_300/Y NOR2X1_67/B NOR2X1_66/Y gnd AOI21X1_52/Y vdd AOI21X1
XAOI21X1_30 BUFX4_97/Y NOR2X1_38/B NOR2X1_38/Y gnd AOI21X1_30/Y vdd AOI21X1
XAOI21X1_63 BUFX4_281/Y NOR2X1_77/B NOR2X1_79/Y gnd AOI21X1_63/Y vdd AOI21X1
XAOI21X1_85 BUFX4_396/Y NOR2X1_103/B AOI21X1_85/C gnd AOI21X1_85/Y vdd AOI21X1
XAOI21X1_74 BUFX4_418/Y NOR2X1_96/B NOR2X1_94/Y gnd AOI21X1_74/Y vdd AOI21X1
XOAI21X1_3 BUFX4_312/Y OAI21X1_1/B INVX1_83/A gnd OAI21X1_4/C vdd OAI21X1
XAOI21X1_96 BUFX4_281/Y NOR2X1_118/B AOI21X1_96/C gnd AOI21X1_96/Y vdd AOI21X1
XBUFX4_316 BUFX4_316/A gnd INVX2_11/A vdd BUFX4
XBUFX4_327 d[5] gnd BUFX4_327/Y vdd BUFX4
XBUFX4_305 INVX8_5/Y gnd BUFX4_305/Y vdd BUFX4
XFILL_46_7_1 gnd vdd FILL
XBUFX4_338 BUFX4_338/A gnd NOR2X1_72/A vdd BUFX4
XBUFX4_349 BUFX4_354/A gnd BUFX4_349/Y vdd BUFX4
XFILL_45_2_0 gnd vdd FILL
XOAI21X1_1206 INVX1_418/Y BUFX4_204/Y NAND2X1_656/Y gnd MUX2X1_310/A vdd OAI21X1
XOAI21X1_1228 INVX1_440/Y BUFX4_248/Y NAND2X1_679/Y gnd MUX2X1_326/A vdd OAI21X1
XOAI21X1_1217 INVX1_429/Y BUFX4_226/Y NAND2X1_668/Y gnd MUX2X1_319/B vdd OAI21X1
XDFFPOSX1_829 NOR2X1_140/A CLKBUF1_21/Y AOI21X1_112/Y gnd vdd DFFPOSX1
XDFFPOSX1_818 INVX1_112/A CLKBUF1_70/Y OAI21X1_615/Y gnd vdd DFFPOSX1
XDFFPOSX1_807 INVX1_431/A CLKBUF1_93/Y OAI21X1_613/Y gnd vdd DFFPOSX1
XOAI21X1_1239 INVX1_451/Y BUFX4_270/Y NAND2X1_692/Y gnd MUX2X1_335/B vdd OAI21X1
XFILL_37_7_1 gnd vdd FILL
XFILL_36_2_0 gnd vdd FILL
XFILL_20_6_1 gnd vdd FILL
XFILL_3_7_1 gnd vdd FILL
XFILL_28_7_1 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XMUX2X1_7 MUX2X1_6/Y MUX2X1_7/B MUX2X1_7/S gnd MUX2X1_7/Y vdd MUX2X1
XFILL_11_6_1 gnd vdd FILL
XFILL_10_1_0 gnd vdd FILL
XCLKBUF1_8 BUFX4_17/Y gnd CLKBUF1_8/Y vdd CLKBUF1
XBUFX4_102 INVX8_7/Y gnd BUFX4_102/Y vdd BUFX4
XBUFX4_113 INVX8_4/Y gnd BUFX4_113/Y vdd BUFX4
XBUFX4_146 INVX8_11/Y gnd BUFX4_146/Y vdd BUFX4
XBUFX4_124 INVX8_2/Y gnd BUFX4_124/Y vdd BUFX4
XFILL_19_7_1 gnd vdd FILL
XBUFX4_135 BUFX4_135/A gnd BUFX4_135/Y vdd BUFX4
XBUFX4_168 BUFX4_168/A gnd BUFX4_168/Y vdd BUFX4
XNOR2X1_206 NOR2X1_206/A NOR2X1_206/B gnd NOR2X1_206/Y vdd NOR2X1
XFILL_18_2_0 gnd vdd FILL
XBUFX4_157 BUFX4_155/A gnd BUFX4_157/Y vdd BUFX4
XBUFX4_179 BUFX4_178/A gnd BUFX4_179/Y vdd BUFX4
XNOR2X1_228 BUFX4_438/Y BUFX4_172/Y gnd NOR2X1_228/Y vdd NOR2X1
XNOR2X1_239 a[4] a[3] gnd BUFX4_354/A vdd NOR2X1
XNOR2X1_217 NOR2X1_217/A NOR2X1_216/B gnd NOR2X1_217/Y vdd NOR2X1
XOAI21X1_1003 INVX1_215/Y BUFX4_194/Y NAND2X1_437/Y gnd MUX2X1_158/B vdd OAI21X1
XOAI21X1_1014 INVX1_226/Y BUFX4_216/Y NAND2X1_449/Y gnd MUX2X1_166/A vdd OAI21X1
XDFFPOSX1_604 OAI21X1_335/C CLKBUF1_47/Y OAI21X1_336/Y gnd vdd DFFPOSX1
XOAI21X1_1036 INVX1_248/Y BUFX4_260/Y NAND2X1_472/Y gnd MUX2X1_182/A vdd OAI21X1
XOAI21X1_1025 INVX1_237/Y BUFX4_238/Y NAND2X1_461/Y gnd MUX2X1_175/B vdd OAI21X1
XDFFPOSX1_626 INVX1_100/A CLKBUF1_60/Y OAI21X1_380/Y gnd vdd DFFPOSX1
XDFFPOSX1_615 INVX1_419/A CLKBUF1_97/Y OAI21X1_358/Y gnd vdd DFFPOSX1
XDFFPOSX1_637 NAND2X1_520/B CLKBUF1_6/Y OAI21X1_402/Y gnd vdd DFFPOSX1
XOAI21X1_1069 INVX1_281/Y BUFX4_227/Y NAND2X1_508/Y gnd MUX2X1_208/B vdd OAI21X1
XDFFPOSX1_648 INVX1_485/A CLKBUF1_83/Y OAI21X1_416/Y gnd vdd DFFPOSX1
XOAI21X1_1058 INVX1_270/Y BUFX4_205/Y NAND2X1_497/Y gnd MUX2X1_199/A vdd OAI21X1
XOAI21X1_1047 INVX1_259/Y MUX2X1_5/S NAND2X1_485/Y gnd MUX2X1_191/B vdd OAI21X1
XINVX1_360 INVX1_360/A gnd INVX1_360/Y vdd INVX1
XDFFPOSX1_659 INVX1_166/A CLKBUF1_85/Y OAI21X1_422/Y gnd vdd DFFPOSX1
XINVX1_371 INVX1_371/A gnd INVX1_371/Y vdd INVX1
XINVX1_393 INVX1_393/A gnd INVX1_393/Y vdd INVX1
XINVX1_382 INVX1_382/A gnd INVX1_382/Y vdd INVX1
XNAND2X1_707 INVX8_1/A NOR2X1_387/A gnd NAND2X1_707/Y vdd NAND2X1
XNAND2X1_718 BUFX4_220/Y NOR2X1_40/A gnd NAND2X1_718/Y vdd NAND2X1
XNAND2X1_729 BUFX4_240/Y NAND2X1_729/B gnd NAND2X1_729/Y vdd NAND2X1
XDFFPOSX1_41 NOR2X1_266/A CLKBUF1_86/Y DFFPOSX1_41/D gnd vdd DFFPOSX1
XDFFPOSX1_63 NOR2X1_292/A CLKBUF1_3/Y DFFPOSX1_63/D gnd vdd DFFPOSX1
XDFFPOSX1_30 INVX1_317/A CLKBUF1_87/Y DFFPOSX1_30/D gnd vdd DFFPOSX1
XDFFPOSX1_52 INVX1_192/A CLKBUF1_31/Y DFFPOSX1_52/D gnd vdd DFFPOSX1
XDFFPOSX1_96 NOR2X1_307/A CLKBUF1_32/Y DFFPOSX1_96/D gnd vdd DFFPOSX1
XDFFPOSX1_85 INVX1_258/A CLKBUF1_43/Y DFFPOSX1_85/D gnd vdd DFFPOSX1
XOAI21X1_1570 BUFX4_410/Y BUFX4_93/Y INVX1_16/A gnd OAI21X1_1570/Y vdd OAI21X1
XOAI21X1_1581 BUFX4_96/Y NAND2X1_840/Y OAI21X1_1581/C gnd DFFPOSX1_254/D vdd OAI21X1
XOAI21X1_1592 BUFX4_454/Y BUFX4_346/Y INVX1_205/A gnd OAI21X1_1592/Y vdd OAI21X1
XDFFPOSX1_74 NAND2X1_276/B CLKBUF1_68/Y DFFPOSX1_74/D gnd vdd DFFPOSX1
XBUFX4_19 BUFX4_70/Y gnd BUFX4_19/Y vdd BUFX4
XFILL_43_5_1 gnd vdd FILL
XFILL_42_0_0 gnd vdd FILL
XFILL_34_5_1 gnd vdd FILL
XFILL_33_0_0 gnd vdd FILL
XOAI21X1_509 BUFX4_414/Y BUFX4_341/Y NAND2X1_662/B gnd OAI21X1_510/C vdd OAI21X1
XFILL_15_1 gnd vdd FILL
XDFFPOSX1_401 INVX1_27/A CLKBUF1_4/Y OAI21X1_74/Y gnd vdd DFFPOSX1
XDFFPOSX1_412 OAI21X1_95/C CLKBUF1_77/Y OAI21X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_456 INVX1_473/A CLKBUF1_50/Y OAI21X1_184/Y gnd vdd DFFPOSX1
XDFFPOSX1_423 INVX1_407/A CLKBUF1_48/Y OAI21X1_118/Y gnd vdd DFFPOSX1
XDFFPOSX1_434 INVX1_88/A CLKBUF1_49/Y OAI21X1_140/Y gnd vdd DFFPOSX1
XDFFPOSX1_445 NAND2X1_507/B CLKBUF1_11/Y OAI21X1_162/Y gnd vdd DFFPOSX1
XDFFPOSX1_478 NOR2X1_18/A CLKBUF1_40/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_489 NOR2X1_23/A CLKBUF1_50/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_467 INVX1_154/A CLKBUF1_2/Y OAI21X1_203/Y gnd vdd DFFPOSX1
XINVX1_190 INVX1_190/A gnd INVX1_190/Y vdd INVX1
XNAND2X1_526 BUFX4_260/Y NOR2X1_87/A gnd NAND2X1_526/Y vdd NAND2X1
XNAND2X1_504 BUFX4_218/Y NOR2X1_7/A gnd NAND2X1_504/Y vdd NAND2X1
XNAND2X1_515 BUFX4_238/Y NOR2X1_57/A gnd NAND2X1_515/Y vdd NAND2X1
XNAND2X1_559 BUFX4_221/Y NAND2X1_559/B gnd NAND2X1_559/Y vdd NAND2X1
XNAND2X1_537 MUX2X1_2/S NOR2X1_173/A gnd NAND2X1_537/Y vdd NAND2X1
XNAND2X1_548 BUFX4_199/Y NOR2X1_261/A gnd NAND2X1_548/Y vdd NAND2X1
XFILL_0_5_1 gnd vdd FILL
XFILL_25_5_1 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XAOI21X1_150 BUFX4_285/Y NOR2X1_186/B NOR2X1_186/Y gnd AOI21X1_150/Y vdd AOI21X1
XAOI21X1_161 BUFX4_131/Y NOR2X1_199/Y NOR2X1_200/Y gnd AOI21X1_161/Y vdd AOI21X1
XAOI21X1_183 BUFX4_102/Y NOR2X1_222/B NOR2X1_225/Y gnd AOI21X1_183/Y vdd AOI21X1
XAOI21X1_194 BUFX4_378/Y NOR2X1_236/B NOR2X1_238/Y gnd AOI21X1_194/Y vdd AOI21X1
XAOI21X1_172 BUFX4_110/Y NOR2X1_216/B NOR2X1_213/Y gnd AOI21X1_172/Y vdd AOI21X1
XFILL_8_6_1 gnd vdd FILL
XDFFPOSX1_990 NOR2X1_216/A CLKBUF1_33/Y AOI21X1_175/Y gnd vdd DFFPOSX1
XFILL_7_1_0 gnd vdd FILL
XFILL_16_5_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XOAI21X1_328 BUFX4_377/Y NAND2X1_77/Y OAI21X1_327/Y gnd OAI21X1_328/Y vdd OAI21X1
XOAI21X1_317 BUFX4_406/Y INVX2_3/A INVX1_162/A gnd OAI21X1_317/Y vdd OAI21X1
XOAI21X1_306 INVX1_97/Y NOR2X1_61/Y NAND2X1_70/Y gnd OAI21X1_306/Y vdd OAI21X1
XOAI21X1_339 BUFX4_87/Y BUFX4_384/Y OAI21X1_339/C gnd OAI21X1_339/Y vdd OAI21X1
XDFFPOSX1_220 NOR2X1_345/A CLKBUF1_5/Y AOI21X1_274/Y gnd vdd DFFPOSX1
XDFFPOSX1_231 INVX1_395/A CLKBUF1_35/Y OAI21X1_1550/Y gnd vdd DFFPOSX1
XBUFX4_4 BUFX4_3/A gnd BUFX4_4/Y vdd BUFX4
XDFFPOSX1_242 INVX1_76/A CLKBUF1_66/Y DFFPOSX1_242/D gnd vdd DFFPOSX1
XDFFPOSX1_253 NAND2X1_494/B CLKBUF1_52/Y OAI21X1_1579/Y gnd vdd DFFPOSX1
XDFFPOSX1_264 INVX1_461/A CLKBUF1_48/Y DFFPOSX1_264/D gnd vdd DFFPOSX1
XNAND2X1_301 BUFX4_238/Y OAI21X1_187/C gnd NAND2X1_301/Y vdd NAND2X1
XDFFPOSX1_297 NOR2X1_370/A CLKBUF1_24/Y AOI21X1_294/Y gnd vdd DFFPOSX1
XDFFPOSX1_286 NOR2X1_365/A CLKBUF1_48/Y AOI21X1_291/Y gnd vdd DFFPOSX1
XDFFPOSX1_275 INVX1_142/A CLKBUF1_39/Y DFFPOSX1_275/D gnd vdd DFFPOSX1
XNAND2X1_345 BUFX4_219/Y DFFPOSX1_75/Q gnd OAI21X1_917/C vdd NAND2X1
XNAND2X1_334 BUFX4_201/Y NOR2X1_203/A gnd OAI21X1_908/C vdd NAND2X1
XNAND2X1_312 BUFX4_258/Y NAND2X1_312/B gnd NAND2X1_312/Y vdd NAND2X1
XNAND2X1_323 BUFX4_278/Y OAI21X1_587/C gnd OAI21X1_897/C vdd NAND2X1
XNAND2X1_356 BUFX4_241/Y NAND2X1_356/B gnd NAND2X1_356/Y vdd NAND2X1
XNAND2X1_367 BUFX4_261/Y OAI21X1_93/C gnd NAND2X1_367/Y vdd NAND2X1
XNAND2X1_378 MUX2X1_4/S NAND2X1_378/B gnd OAI21X1_948/C vdd NAND2X1
XNAND2X1_389 BUFX4_204/Y NOR2X1_95/A gnd OAI21X1_959/C vdd NAND2X1
XFILL_40_3_1 gnd vdd FILL
XOAI21X1_840 INVX1_52/Y BUFX4_264/Y OAI21X1_840/C gnd MUX2X1_35/A vdd OAI21X1
XOAI21X1_851 INVX1_63/Y MUX2X1_12/S OAI21X1_851/C gnd MUX2X1_44/B vdd OAI21X1
XOAI21X1_884 INVX1_96/Y BUFX4_253/Y OAI21X1_884/C gnd MUX2X1_68/A vdd OAI21X1
XOAI21X1_862 INVX1_74/Y BUFX4_209/Y OAI21X1_862/C gnd MUX2X1_52/A vdd OAI21X1
XOAI21X1_873 INVX1_85/Y BUFX4_231/Y NAND2X1_297/Y gnd MUX2X1_61/B vdd OAI21X1
XOAI21X1_895 INVX1_107/Y BUFX4_275/Y NAND2X1_320/Y gnd MUX2X1_77/B vdd OAI21X1
XMUX2X1_340 MUX2X1_340/A MUX2X1_340/B BUFX4_43/Y gnd MUX2X1_340/Y vdd MUX2X1
XMUX2X1_373 MUX2X1_373/A MUX2X1_373/B BUFX4_32/Y gnd MUX2X1_373/Y vdd MUX2X1
XMUX2X1_362 MUX2X1_362/A MUX2X1_362/B MUX2X1_3/S gnd MUX2X1_362/Y vdd MUX2X1
XMUX2X1_351 MUX2X1_351/A MUX2X1_349/Y BUFX4_362/Y gnd AOI22X1_73/A vdd MUX2X1
XFILL_48_4_1 gnd vdd FILL
XFILL_31_3_1 gnd vdd FILL
XNAND3X1_7 we BUFX4_349/Y AOI22X1_9/A gnd NAND3X1_7/Y vdd NAND3X1
XFILL_39_4_1 gnd vdd FILL
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_103 BUFX4_86/Y INVX2_1/A NAND2X1_712/B gnd OAI21X1_103/Y vdd OAI21X1
XOAI21X1_136 BUFX4_374/Y NAND2X1_17/Y OAI21X1_135/Y gnd OAI21X1_136/Y vdd OAI21X1
XOAI21X1_147 INVX4_3/A BUFX4_175/Y INVX1_344/A gnd OAI21X1_148/C vdd OAI21X1
XOAI21X1_114 BUFX4_399/Y NAND2X1_16/Y OAI21X1_114/C gnd OAI21X1_114/Y vdd OAI21X1
XOAI21X1_125 NOR2X1_52/B BUFX4_178/Y NAND2X1_368/B gnd OAI21X1_125/Y vdd OAI21X1
XOAI21X1_169 BUFX4_457/Y BUFX4_134/Y INVX1_32/A gnd OAI21X1_169/Y vdd OAI21X1
XOAI21X1_158 BUFX4_116/Y NAND2X1_19/Y OAI21X1_158/C gnd OAI21X1_158/Y vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd q[0] vdd BUFX2
XNAND2X1_142 BUFX4_452/Y NOR2X1_133/Y gnd OAI21X1_615/C vdd NAND2X1
XNAND2X1_120 NAND2X1_9/A NOR2X1_101/Y gnd NAND2X1_120/Y vdd NAND2X1
XNAND2X1_153 BUFX4_335/Y NOR2X1_145/B gnd OAI21X1_655/C vdd NAND2X1
XNAND2X1_131 BUFX4_445/Y NOR2X1_111/Y gnd OAI21X1_604/C vdd NAND2X1
XNAND2X1_186 BUFX4_447/Y NOR2X1_189/B gnd OAI21X1_717/C vdd NAND2X1
XNAND2X1_175 INVX8_11/A INVX1_5/Y gnd OAI21X1_704/B vdd NAND2X1
XFILL_5_4_1 gnd vdd FILL
XNAND2X1_164 BUFX4_136/Y NOR2X1_155/Y gnd NAND2X1_164/Y vdd NAND2X1
XNAND2X1_197 BUFX4_290/Y AOI22X1_69/C gnd BUFX4_439/A vdd NAND2X1
XFILL_13_3_1 gnd vdd FILL
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 AOI21X1_1/A NOR2X1_2/Y NOR2X1_3/Y gnd AOI21X1_1/Y vdd AOI21X1
XOAI21X1_670 INVX1_244/Y NOR2X1_166/Y NAND2X1_168/Y gnd OAI21X1_670/Y vdd OAI21X1
XOAI21X1_681 BUFX4_462/Y BUFX4_67/Y INVX1_245/A gnd OAI21X1_682/C vdd OAI21X1
XOAI21X1_692 BUFX4_131/Y OAI21X1_704/B OAI21X1_692/C gnd OAI21X1_692/Y vdd OAI21X1
XMUX2X1_170 MUX2X1_170/A MUX2X1_170/B BUFX4_35/Y gnd MUX2X1_170/Y vdd MUX2X1
XMUX2X1_181 MUX2X1_181/A MUX2X1_181/B BUFX4_82/Y gnd MUX2X1_181/Y vdd MUX2X1
XMUX2X1_192 MUX2X1_191/Y MUX2X1_192/B BUFX4_364/Y gnd AOI22X1_40/D vdd MUX2X1
XAOI21X1_42 BUFX4_418/Y NOR2X1_55/B NOR2X1_54/Y gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_53 BUFX4_398/Y NOR2X1_67/B NOR2X1_67/Y gnd AOI21X1_53/Y vdd AOI21X1
XAOI21X1_20 BUFX4_304/Y NOR2X1_27/B NOR2X1_26/Y gnd AOI21X1_20/Y vdd AOI21X1
XAOI21X1_31 BUFX4_279/Y NOR2X1_38/B NOR2X1_39/Y gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_64 BUFX4_374/Y NOR2X1_77/B NOR2X1_80/Y gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_86 BUFX4_103/Y NOR2X1_103/B NOR2X1_108/Y gnd AOI21X1_86/Y vdd AOI21X1
XAOI21X1_75 AOI21X1_3/A NOR2X1_96/B NOR2X1_95/Y gnd AOI21X1_75/Y vdd AOI21X1
XOAI21X1_4 BUFX4_424/Y NAND2X1_1/Y OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_97 BUFX4_372/Y NOR2X1_118/B NOR2X1_121/Y gnd AOI21X1_97/Y vdd AOI21X1
XBUFX4_317 BUFX4_316/A gnd BUFX4_317/Y vdd BUFX4
XBUFX4_306 INVX8_14/Y gnd NOR2X1_21/B vdd BUFX4
XBUFX4_328 d[5] gnd INVX8_7/A vdd BUFX4
XBUFX4_339 BUFX4_338/A gnd INVX2_4/A vdd BUFX4
XFILL_45_2_1 gnd vdd FILL
XOAI21X1_1207 INVX1_419/Y BUFX4_206/Y NAND2X1_657/Y gnd MUX2X1_311/B vdd OAI21X1
XOAI21X1_1229 INVX1_441/Y BUFX4_250/Y NAND2X1_680/Y gnd MUX2X1_328/B vdd OAI21X1
XOAI21X1_1218 INVX1_430/Y BUFX4_228/Y NAND2X1_669/Y gnd MUX2X1_319/A vdd OAI21X1
XDFFPOSX1_819 INVX1_176/A CLKBUF1_83/Y OAI21X1_616/Y gnd vdd DFFPOSX1
XDFFPOSX1_808 INVX1_495/A CLKBUF1_69/Y OAI21X1_614/Y gnd vdd DFFPOSX1
XFILL_45_1 gnd vdd FILL
XFILL_36_2_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XFILL_27_2_1 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A MUX2X1_8/B MUX2X1_8/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 BUFX4_16/Y gnd CLKBUF1_9/Y vdd CLKBUF1
XBUFX4_103 INVX8_7/Y gnd BUFX4_103/Y vdd BUFX4
XBUFX4_136 d[6] gnd BUFX4_136/Y vdd BUFX4
XBUFX4_114 INVX8_4/Y gnd BUFX4_114/Y vdd BUFX4
XBUFX4_125 INVX8_2/Y gnd BUFX4_125/Y vdd BUFX4
XNOR2X1_207 NOR2X1_207/A NOR2X1_206/B gnd NOR2X1_207/Y vdd NOR2X1
XBUFX4_169 BUFX4_168/A gnd BUFX4_169/Y vdd BUFX4
XBUFX4_147 INVX8_11/Y gnd BUFX4_147/Y vdd BUFX4
XFILL_18_2_1 gnd vdd FILL
XBUFX4_158 BUFX4_155/A gnd AOI22X1_7/C vdd BUFX4
XNOR2X1_229 MUX2X1_26/B NOR2X1_228/Y gnd NOR2X1_229/Y vdd NOR2X1
XNOR2X1_218 NOR2X1_218/A NOR2X1_216/B gnd NOR2X1_218/Y vdd NOR2X1
XOAI21X1_1004 INVX1_216/Y BUFX4_196/Y NAND2X1_438/Y gnd MUX2X1_158/A vdd OAI21X1
XOAI21X1_1015 INVX1_227/Y BUFX4_218/Y NAND2X1_450/Y gnd MUX2X1_167/B vdd OAI21X1
XDFFPOSX1_605 NAND2X1_518/B CLKBUF1_47/Y OAI21X1_338/Y gnd vdd DFFPOSX1
XOAI21X1_1037 INVX1_249/Y BUFX4_262/Y NAND2X1_473/Y gnd MUX2X1_184/B vdd OAI21X1
XOAI21X1_1026 INVX1_238/Y BUFX4_240/Y NAND2X1_462/Y gnd MUX2X1_175/A vdd OAI21X1
XDFFPOSX1_627 INVX1_164/A CLKBUF1_10/Y OAI21X1_382/Y gnd vdd DFFPOSX1
XDFFPOSX1_616 INVX1_483/A CLKBUF1_16/Y OAI21X1_360/Y gnd vdd DFFPOSX1
XDFFPOSX1_638 NAND2X1_589/B CLKBUF1_10/Y OAI21X1_404/Y gnd vdd DFFPOSX1
XOAI21X1_1059 INVX1_271/Y BUFX4_207/Y NAND2X1_498/Y gnd MUX2X1_200/B vdd OAI21X1
XOAI21X1_1048 INVX1_260/Y MUX2X1_9/S NAND2X1_486/Y gnd MUX2X1_191/A vdd OAI21X1
XDFFPOSX1_649 NOR2X1_73/A CLKBUF1_33/Y AOI21X1_57/Y gnd vdd DFFPOSX1
XINVX1_361 INVX1_361/A gnd INVX1_361/Y vdd INVX1
XINVX1_350 INVX1_350/A gnd INVX1_350/Y vdd INVX1
XNAND2X1_708 BUFX4_200/Y NAND2X1_708/B gnd NAND2X1_708/Y vdd NAND2X1
XINVX1_394 INVX1_394/A gnd INVX1_394/Y vdd INVX1
XINVX1_383 INVX1_383/A gnd INVX1_383/Y vdd INVX1
XNAND2X1_719 AOI22X1_72/Y AOI22X1_73/Y gnd AOI22X1_74/D vdd NAND2X1
XINVX1_372 INVX1_372/A gnd INVX1_372/Y vdd INVX1
XDFFPOSX1_20 NOR2X1_279/A CLKBUF1_44/Y AOI21X1_226/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 NOR2X1_267/A CLKBUF1_90/Y AOI21X1_216/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 INVX1_381/A CLKBUF1_23/Y DFFPOSX1_31/D gnd vdd DFFPOSX1
XDFFPOSX1_53 INVX1_256/A CLKBUF1_71/Y DFFPOSX1_53/D gnd vdd DFFPOSX1
XDFFPOSX1_75 DFFPOSX1_75/Q CLKBUF1_43/Y DFFPOSX1_75/D gnd vdd DFFPOSX1
XOAI21X1_1582 BUFX4_410/Y BUFX4_91/Y NAND2X1_632/B gnd OAI21X1_1583/C vdd OAI21X1
XOAI21X1_1571 BUFX4_128/Y NAND2X1_840/Y OAI21X1_1570/Y gnd OAI21X1_1571/Y vdd OAI21X1
XOAI21X1_1560 BUFX4_171/Y BUFX4_95/Y INVX1_204/A gnd OAI21X1_1561/C vdd OAI21X1
XDFFPOSX1_64 NOR2X1_293/A CLKBUF1_30/Y DFFPOSX1_64/D gnd vdd DFFPOSX1
XOAI21X1_1593 BUFX4_297/Y NAND2X1_842/Y OAI21X1_1592/Y gnd DFFPOSX1_260/D vdd OAI21X1
XDFFPOSX1_86 INVX1_322/A CLKBUF1_39/Y DFFPOSX1_86/D gnd vdd DFFPOSX1
XDFFPOSX1_97 INVX1_39/A CLKBUF1_55/Y DFFPOSX1_97/D gnd vdd DFFPOSX1
XFILL_42_0_1 gnd vdd FILL
XFILL_33_0_1 gnd vdd FILL
XDFFPOSX1_402 INVX1_86/A CLKBUF1_100/Y OAI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_413 OAI21X1_97/C CLKBUF1_4/Y OAI21X1_98/Y gnd vdd DFFPOSX1
XDFFPOSX1_424 INVX1_471/A CLKBUF1_41/Y OAI21X1_120/Y gnd vdd DFFPOSX1
XDFFPOSX1_446 OAI21X1_163/C CLKBUF1_82/Y OAI21X1_164/Y gnd vdd DFFPOSX1
XDFFPOSX1_435 INVX1_152/A CLKBUF1_11/Y OAI21X1_142/Y gnd vdd DFFPOSX1
XDFFPOSX1_457 NAND2X1_229/B CLKBUF1_87/Y OAI21X1_186/Y gnd vdd DFFPOSX1
XDFFPOSX1_468 INVX1_218/A CLKBUF1_3/Y OAI21X1_204/Y gnd vdd DFFPOSX1
XDFFPOSX1_479 NOR2X1_19/A CLKBUF1_23/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XINVX1_191 INVX1_191/A gnd INVX1_191/Y vdd INVX1
XNAND2X1_527 BUFX4_262/Y NOR2X1_97/A gnd NAND2X1_527/Y vdd NAND2X1
XNAND2X1_505 BUFX4_220/Y OAI21X1_97/C gnd NAND2X1_505/Y vdd NAND2X1
XNAND2X1_516 BUFX4_240/Y NAND2X1_516/B gnd NAND2X1_516/Y vdd NAND2X1
XNAND2X1_549 BUFX4_201/Y NOR2X1_271/A gnd NAND2X1_549/Y vdd NAND2X1
XNAND2X1_538 MUX2X1_5/S NAND2X1_538/B gnd NAND2X1_538/Y vdd NAND2X1
XFILL_24_0_1 gnd vdd FILL
XAOI21X1_151 BUFX4_375/Y NOR2X1_186/B NOR2X1_187/Y gnd AOI21X1_151/Y vdd AOI21X1
XAOI21X1_140 BUFX4_104/Y NOR2X1_173/B NOR2X1_174/Y gnd AOI21X1_140/Y vdd AOI21X1
XAOI21X1_162 BUFX4_131/Y NOR2X1_206/B NOR2X1_202/Y gnd AOI21X1_162/Y vdd AOI21X1
XAOI21X1_184 BUFX4_284/Y NOR2X1_222/B NOR2X1_226/Y gnd AOI21X1_184/Y vdd AOI21X1
XAOI21X1_173 BUFX4_298/Y NOR2X1_216/B NOR2X1_214/Y gnd AOI21X1_173/Y vdd AOI21X1
XAOI21X1_195 AOI21X1_195/A NOR2X1_246/Y BUFX4_92/Y gnd AOI21X1_195/Y vdd AOI21X1
XOAI21X1_1390 NAND2X1_811/Y BUFX4_286/Y OAI21X1_1389/Y gnd OAI21X1_1390/Y vdd OAI21X1
XDFFPOSX1_980 INVX1_250/A CLKBUF1_65/Y OAI21X1_767/Y gnd vdd DFFPOSX1
XDFFPOSX1_991 NOR2X1_217/A CLKBUF1_88/Y AOI21X1_176/Y gnd vdd DFFPOSX1
XFILL_7_1_1 gnd vdd FILL
XFILL_44_8_0 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XFILL_35_8_0 gnd vdd FILL
XOAI21X1_307 INVX1_161/Y NOR2X1_61/Y NAND2X1_71/Y gnd OAI21X1_307/Y vdd OAI21X1
XOAI21X1_329 BUFX4_87/Y BUFX4_386/Y NAND2X1_260/B gnd OAI21X1_330/C vdd OAI21X1
XOAI21X1_318 BUFX4_109/Y NAND2X1_77/Y OAI21X1_317/Y gnd OAI21X1_318/Y vdd OAI21X1
XDFFPOSX1_221 NOR2X1_346/A CLKBUF1_76/Y AOI21X1_275/Y gnd vdd DFFPOSX1
XDFFPOSX1_210 INVX1_74/A CLKBUF1_52/Y DFFPOSX1_210/D gnd vdd DFFPOSX1
XBUFX4_5 BUFX4_8/A gnd BUFX4_5/Y vdd BUFX4
XDFFPOSX1_243 INVX1_140/A CLKBUF1_5/Y OAI21X1_1559/Y gnd vdd DFFPOSX1
XDFFPOSX1_254 NAND2X1_563/B CLKBUF1_52/Y DFFPOSX1_254/D gnd vdd DFFPOSX1
XDFFPOSX1_232 INVX1_459/A CLKBUF1_64/Y DFFPOSX1_232/D gnd vdd DFFPOSX1
XNAND2X1_302 BUFX4_240/Y NOR2X1_14/A gnd OAI21X1_878/C vdd NAND2X1
XDFFPOSX1_276 INVX1_206/A CLKBUF1_30/Y DFFPOSX1_276/D gnd vdd DFFPOSX1
XDFFPOSX1_287 NOR2X1_366/A CLKBUF1_75/Y AOI21X1_292/Y gnd vdd DFFPOSX1
XDFFPOSX1_265 NAND2X1_217/B CLKBUF1_12/Y OAI21X1_1603/Y gnd vdd DFFPOSX1
XDFFPOSX1_298 NOR2X1_371/A CLKBUF1_68/Y AOI21X1_295/Y gnd vdd DFFPOSX1
XNAND2X1_313 BUFX4_260/Y NAND2X1_313/B gnd NAND2X1_313/Y vdd NAND2X1
XNAND2X1_335 BUFX4_203/Y NAND2X1_335/B gnd NAND2X1_335/Y vdd NAND2X1
XNAND2X1_324 MUX2X1_2/S NOR2X1_115/A gnd NAND2X1_324/Y vdd NAND2X1
XNAND2X1_346 BUFX4_221/Y NOR2X1_302/A gnd OAI21X1_918/C vdd NAND2X1
XNAND2X1_357 AOI22X1_20/Y AOI22X1_21/Y gnd AOI22X1_24/A vdd NAND2X1
XNAND2X1_368 BUFX4_263/Y NAND2X1_368/B gnd NAND2X1_368/Y vdd NAND2X1
XNAND2X1_379 MUX2X1_8/S NOR2X1_65/A gnd NAND2X1_379/Y vdd NAND2X1
XFILL_26_8_0 gnd vdd FILL
XFILL_1_8_0 gnd vdd FILL
XOAI21X1_841 INVX1_53/Y BUFX4_266/Y OAI21X1_841/C gnd MUX2X1_37/B vdd OAI21X1
XOAI21X1_830 INVX1_43/Y BUFX4_246/Y OAI21X1_830/C gnd NAND2X1_252/B vdd OAI21X1
XOAI21X1_863 INVX1_75/Y BUFX4_211/Y NAND2X1_286/Y gnd MUX2X1_53/B vdd OAI21X1
XOAI21X1_885 INVX1_97/Y BUFX4_255/Y NAND2X1_310/Y gnd MUX2X1_70/B vdd OAI21X1
XOAI21X1_852 INVX1_64/Y BUFX4_189/Y NAND2X1_275/Y gnd MUX2X1_44/A vdd OAI21X1
XOAI21X1_874 INVX1_86/Y BUFX4_233/Y OAI21X1_874/C gnd MUX2X1_61/A vdd OAI21X1
XOAI21X1_896 INVX1_108/Y BUFX4_277/Y OAI21X1_896/C gnd MUX2X1_77/A vdd OAI21X1
XMUX2X1_341 MUX2X1_341/A MUX2X1_341/B BUFX4_59/Y gnd MUX2X1_341/Y vdd MUX2X1
XMUX2X1_330 MUX2X1_329/Y MUX2X1_330/B MUX2X1_7/S gnd MUX2X1_330/Y vdd MUX2X1
XMUX2X1_363 MUX2X1_362/Y MUX2X1_361/Y MUX2X1_7/S gnd MUX2X1_363/Y vdd MUX2X1
XMUX2X1_374 MUX2X1_374/A MUX2X1_374/B BUFX4_52/Y gnd MUX2X1_375/A vdd MUX2X1
XMUX2X1_352 MUX2X1_352/A MUX2X1_352/B BUFX4_55/Y gnd MUX2X1_352/Y vdd MUX2X1
XFILL_17_8_0 gnd vdd FILL
XOAI21X1_104 BUFX4_374/Y OAI21X1_96/B OAI21X1_103/Y gnd OAI21X1_104/Y vdd OAI21X1
XOAI21X1_137 INVX4_3/A BUFX4_179/Y INVX1_25/A gnd OAI21X1_137/Y vdd OAI21X1
XOAI21X1_115 NOR2X1_91/B BUFX4_178/Y INVX1_343/A gnd OAI21X1_115/Y vdd OAI21X1
XOAI21X1_126 BUFX4_116/Y NAND2X1_17/Y OAI21X1_125/Y gnd OAI21X1_126/Y vdd OAI21X1
XOAI21X1_148 NAND2X1_18/Y AOI21X1_6/A OAI21X1_148/C gnd OAI21X1_148/Y vdd OAI21X1
XOAI21X1_159 BUFX4_411/Y BUFX4_178/Y OAI21X1_159/C gnd OAI21X1_160/C vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd q[1] vdd BUFX2
XNAND2X1_110 BUFX4_453/Y NOR2X1_91/Y gnd OAI21X1_554/C vdd NAND2X1
XNAND2X1_143 BUFX4_334/Y NOR2X1_133/Y gnd OAI21X1_616/C vdd NAND2X1
XNAND2X1_121 BUFX4_444/Y NOR2X1_101/Y gnd OAI21X1_565/C vdd NAND2X1
XNAND2X1_132 BUFX4_327/Y NOR2X1_111/Y gnd NAND2X1_132/Y vdd NAND2X1
XNAND2X1_165 BUFX4_427/Y NOR2X1_155/Y gnd OAI21X1_667/C vdd NAND2X1
XNAND2X1_176 INVX8_3/A NOR2X1_177/Y gnd OAI21X1_707/C vdd NAND2X1
XNAND2X1_187 BUFX4_329/Y NOR2X1_189/B gnd NAND2X1_187/Y vdd NAND2X1
XNAND2X1_154 BUFX4_145/Y NOR2X1_145/B gnd OAI21X1_656/C vdd NAND2X1
XNAND2X1_198 INVX8_10/A INVX2_5/Y gnd OAI21X1_729/B vdd NAND2X1
XFILL_41_6_0 gnd vdd FILL
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XOAI21X1_660 INVX1_498/Y NOR2X1_145/B OAI21X1_660/C gnd OAI21X1_660/Y vdd OAI21X1
XOAI21X1_693 BUFX4_147/Y BUFX4_64/Y OAI21X1_693/C gnd OAI21X1_693/Y vdd OAI21X1
XOAI21X1_682 BUFX4_301/Y NAND2X1_174/Y OAI21X1_682/C gnd OAI21X1_682/Y vdd OAI21X1
XAOI21X1_2 BUFX4_425/Y NOR2X1_2/Y NOR2X1_4/Y gnd AOI21X1_2/Y vdd AOI21X1
XOAI21X1_671 INVX1_308/Y NOR2X1_166/Y NAND2X1_169/Y gnd OAI21X1_671/Y vdd OAI21X1
XMUX2X1_182 MUX2X1_182/A MUX2X1_182/B MUX2X1_3/S gnd MUX2X1_182/Y vdd MUX2X1
XMUX2X1_160 MUX2X1_160/A MUX2X1_160/B BUFX4_43/Y gnd MUX2X1_160/Y vdd MUX2X1
XMUX2X1_171 MUX2X1_170/Y MUX2X1_171/B BUFX4_357/Y gnd MUX2X1_171/Y vdd MUX2X1
XMUX2X1_193 MUX2X1_193/A MUX2X1_193/B BUFX4_32/Y gnd MUX2X1_195/B vdd MUX2X1
XFILL_32_6_0 gnd vdd FILL
XFILL_23_6_0 gnd vdd FILL
XAOI21X1_10 BUFX4_423/Y NOR2X1_14/B NOR2X1_14/Y gnd AOI21X1_10/Y vdd AOI21X1
XAOI21X1_43 BUFX4_114/Y NOR2X1_55/B NOR2X1_55/Y gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_32 BUFX4_374/Y NOR2X1_38/B NOR2X1_40/Y gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_21 BUFX4_395/Y NOR2X1_27/B NOR2X1_27/Y gnd AOI21X1_21/Y vdd AOI21X1
XAOI21X1_54 BUFX4_101/Y NOR2X1_67/B NOR2X1_68/Y gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_76 BUFX4_298/Y NOR2X1_96/B NOR2X1_96/Y gnd AOI21X1_76/Y vdd AOI21X1
XAOI21X1_65 BUFX4_127/Y NOR2X1_90/B NOR2X1_83/Y gnd AOI21X1_65/Y vdd AOI21X1
XOAI21X1_5 BUFX4_310/Y OAI21X1_5/B INVX1_147/A gnd OAI21X1_6/C vdd OAI21X1
XAOI21X1_98 BUFX4_130/Y NOR2X1_122/Y NOR2X1_123/Y gnd AOI21X1_98/Y vdd AOI21X1
XAOI21X1_87 BUFX4_280/Y NOR2X1_103/B NOR2X1_109/Y gnd AOI21X1_87/Y vdd AOI21X1
XFILL_6_7_0 gnd vdd FILL
XBUFX4_307 INVX8_14/Y gnd BUFX4_307/Y vdd BUFX4
XBUFX4_318 BUFX4_316/A gnd OAI21X1_7/B vdd BUFX4
XBUFX4_329 d[5] gnd BUFX4_329/Y vdd BUFX4
XFILL_14_6_0 gnd vdd FILL
XOAI21X1_1208 INVX1_420/Y BUFX4_208/Y NAND2X1_658/Y gnd MUX2X1_311/A vdd OAI21X1
XOAI21X1_1219 INVX1_431/Y BUFX4_230/Y NAND2X1_670/Y gnd MUX2X1_320/B vdd OAI21X1
XOAI21X1_490 NAND2X1_96/Y BUFX4_400/Y OAI21X1_489/Y gnd OAI21X1_490/Y vdd OAI21X1
XDFFPOSX1_809 MUX2X1_4/A CLKBUF1_74/Y AOI21X1_99/Y gnd vdd DFFPOSX1
XFILL_45_2 gnd vdd FILL
XFILL_38_1 gnd vdd FILL
XMUX2X1_9 MUX2X1_9/A MUX2X1_9/B MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XBUFX4_115 INVX8_4/Y gnd BUFX4_115/Y vdd BUFX4
XBUFX4_137 d[6] gnd BUFX4_137/Y vdd BUFX4
XBUFX4_104 INVX8_7/Y gnd BUFX4_104/Y vdd BUFX4
XBUFX4_126 INVX8_2/Y gnd BUFX4_126/Y vdd BUFX4
XFILL_46_5_0 gnd vdd FILL
XBUFX4_159 BUFX4_155/A gnd BUFX4_159/Y vdd BUFX4
XBUFX4_148 INVX8_11/Y gnd BUFX4_148/Y vdd BUFX4
XNOR2X1_208 NOR2X1_208/A NOR2X1_206/B gnd NOR2X1_208/Y vdd NOR2X1
XNOR2X1_219 BUFX4_438/Y BUFX4_370/Y gnd NOR2X1_222/B vdd NOR2X1
XOAI21X1_1016 INVX1_228/Y BUFX4_220/Y NAND2X1_451/Y gnd MUX2X1_167/A vdd OAI21X1
XOAI21X1_1005 INVX1_217/Y INVX8_1/A NAND2X1_439/Y gnd MUX2X1_160/B vdd OAI21X1
XOAI21X1_1027 INVX1_239/Y BUFX4_242/Y NAND2X1_463/Y gnd MUX2X1_176/B vdd OAI21X1
XDFFPOSX1_617 NAND2X1_261/B CLKBUF1_6/Y OAI21X1_362/Y gnd vdd DFFPOSX1
XDFFPOSX1_628 INVX1_228/A CLKBUF1_6/Y OAI21X1_384/Y gnd vdd DFFPOSX1
XDFFPOSX1_606 OAI21X1_339/C CLKBUF1_60/Y OAI21X1_340/Y gnd vdd DFFPOSX1
XDFFPOSX1_639 NAND2X1_658/B CLKBUF1_60/Y OAI21X1_406/Y gnd vdd DFFPOSX1
XOAI21X1_1038 INVX1_250/Y BUFX4_264/Y NAND2X1_474/Y gnd MUX2X1_184/A vdd OAI21X1
XOAI21X1_1049 INVX1_261/Y MUX2X1_12/S NAND2X1_487/Y gnd MUX2X1_193/B vdd OAI21X1
XINVX1_340 INVX1_340/A gnd INVX1_340/Y vdd INVX1
XINVX1_362 INVX1_362/A gnd INVX1_362/Y vdd INVX1
XINVX1_351 INVX1_351/A gnd INVX1_351/Y vdd INVX1
XNAND2X1_709 BUFX4_202/Y OAI21X1_31/C gnd NAND2X1_709/Y vdd NAND2X1
XINVX1_373 INVX1_373/A gnd INVX1_373/Y vdd INVX1
XINVX1_395 INVX1_395/A gnd INVX1_395/Y vdd INVX1
XINVX1_384 INVX1_384/A gnd INVX1_384/Y vdd INVX1
XFILL_37_5_0 gnd vdd FILL
XAOI21X1_300 BUFX4_279/Y NOR2X1_373/B NOR2X1_376/Y gnd AOI21X1_300/Y vdd AOI21X1
XFILL_20_4_0 gnd vdd FILL
XDFFPOSX1_10 NOR2X1_257/A CLKBUF1_5/Y AOI21X1_208/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 NOR2X1_268/A CLKBUF1_76/Y DFFPOSX1_43/D gnd vdd DFFPOSX1
XOAI21X1_1550 NAND2X1_837/Y BUFX4_282/Y OAI21X1_1550/C gnd OAI21X1_1550/Y vdd OAI21X1
XDFFPOSX1_54 INVX1_320/A CLKBUF1_3/Y DFFPOSX1_54/D gnd vdd DFFPOSX1
XDFFPOSX1_32 INVX1_445/A CLKBUF1_56/Y DFFPOSX1_32/D gnd vdd DFFPOSX1
XDFFPOSX1_21 NOR2X1_280/A CLKBUF1_37/Y AOI21X1_227/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 DFFPOSX1_76/Q CLKBUF1_42/Y DFFPOSX1_76/D gnd vdd DFFPOSX1
XDFFPOSX1_65 INVX1_37/A CLKBUF1_84/Y DFFPOSX1_65/D gnd vdd DFFPOSX1
XOAI21X1_1583 BUFX4_282/Y NAND2X1_840/Y OAI21X1_1583/C gnd DFFPOSX1_255/D vdd OAI21X1
XOAI21X1_1561 NAND2X1_839/Y BUFX4_303/Y OAI21X1_1561/C gnd DFFPOSX1_244/D vdd OAI21X1
XOAI21X1_1572 BUFX4_410/Y BUFX4_95/Y NAND2X1_287/B gnd OAI21X1_1573/C vdd OAI21X1
XDFFPOSX1_87 INVX1_386/A CLKBUF1_20/Y DFFPOSX1_87/D gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX1_67/A CLKBUF1_75/Y DFFPOSX1_98/D gnd vdd DFFPOSX1
XOAI21X1_1594 BUFX4_454/Y BUFX4_348/Y INVX1_269/A gnd OAI21X1_1595/C vdd OAI21X1
XFILL_3_5_0 gnd vdd FILL
XFILL_28_5_0 gnd vdd FILL
XFILL_11_4_0 gnd vdd FILL
XFILL_19_5_0 gnd vdd FILL
XDFFPOSX1_403 INVX1_150/A CLKBUF1_29/Y OAI21X1_78/Y gnd vdd DFFPOSX1
XDFFPOSX1_414 OAI21X1_99/C CLKBUF1_29/Y OAI21X1_100/Y gnd vdd DFFPOSX1
XDFFPOSX1_425 OAI21X1_121/C CLKBUF1_77/Y OAI21X1_122/Y gnd vdd DFFPOSX1
XDFFPOSX1_447 NAND2X1_645/B CLKBUF1_77/Y OAI21X1_166/Y gnd vdd DFFPOSX1
XDFFPOSX1_436 INVX1_216/A CLKBUF1_27/Y OAI21X1_144/Y gnd vdd DFFPOSX1
XDFFPOSX1_458 OAI21X1_187/C CLKBUF1_50/Y OAI21X1_188/Y gnd vdd DFFPOSX1
XDFFPOSX1_469 INVX1_282/A CLKBUF1_18/Y OAI21X1_205/Y gnd vdd DFFPOSX1
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XNAND2X1_517 BUFX4_242/Y NOR2X1_67/A gnd NAND2X1_517/Y vdd NAND2X1
XINVX1_192 INVX1_192/A gnd INVX1_192/Y vdd INVX1
XNAND2X1_506 BUFX4_222/Y NAND2X1_506/B gnd NAND2X1_506/Y vdd NAND2X1
XNAND2X1_539 MUX2X1_9/S NOR2X1_184/A gnd NAND2X1_539/Y vdd NAND2X1
XNAND2X1_528 BUFX4_264/Y NOR2X1_107/A gnd NAND2X1_528/Y vdd NAND2X1
XAOI21X1_130 BUFX4_394/Y NOR2X1_158/B NOR2X1_162/Y gnd AOI21X1_130/Y vdd AOI21X1
XAOI21X1_141 BUFX4_286/Y NOR2X1_173/B NOR2X1_175/Y gnd AOI21X1_141/Y vdd AOI21X1
XAOI21X1_152 BUFX4_131/Y NOR2X1_189/B NOR2X1_189/Y gnd AOI21X1_152/Y vdd AOI21X1
XAOI21X1_163 BUFX4_426/Y NOR2X1_206/B NOR2X1_203/Y gnd AOI21X1_163/Y vdd AOI21X1
XAOI21X1_185 BUFX4_378/Y NOR2X1_222/B NOR2X1_227/Y gnd AOI21X1_185/Y vdd AOI21X1
XAOI21X1_174 BUFX4_400/Y NOR2X1_216/B NOR2X1_215/Y gnd AOI21X1_174/Y vdd AOI21X1
XAOI21X1_196 INVX8_1/Y INVX1_17/Y OR2X2_1/A gnd AOI21X1_196/Y vdd AOI21X1
XOAI21X1_1380 NAND2X1_811/Y BUFX4_422/Y OAI21X1_1380/C gnd DFFPOSX1_114/D vdd OAI21X1
XOAI21X1_1391 BUFX4_167/Y INVX2_7/A INVX1_452/A gnd OAI21X1_1392/C vdd OAI21X1
XDFFPOSX1_992 NOR2X1_218/A CLKBUF1_73/Y AOI21X1_177/Y gnd vdd DFFPOSX1
XDFFPOSX1_981 INVX1_314/A CLKBUF1_67/Y OAI21X1_769/Y gnd vdd DFFPOSX1
XDFFPOSX1_970 NAND2X1_335/B CLKBUF1_59/Y OAI21X1_747/Y gnd vdd DFFPOSX1
XFILL_44_8_1 gnd vdd FILL
XFILL_43_3_0 gnd vdd FILL
XFILL_35_8_1 gnd vdd FILL
XFILL_34_3_0 gnd vdd FILL
XOAI21X1_319 BUFX4_404/Y INVX2_3/A INVX1_226/A gnd OAI21X1_320/C vdd OAI21X1
XOAI21X1_308 INVX1_225/Y NOR2X1_61/Y NAND2X1_72/Y gnd OAI21X1_308/Y vdd OAI21X1
XDFFPOSX1_211 INVX1_138/A CLKBUF1_76/Y DFFPOSX1_211/D gnd vdd DFFPOSX1
XDFFPOSX1_222 NOR2X1_347/A CLKBUF1_35/Y AOI21X1_276/Y gnd vdd DFFPOSX1
XDFFPOSX1_200 INVX1_457/A CLKBUF1_36/Y OAI21X1_1504/Y gnd vdd DFFPOSX1
XBUFX4_6 BUFX4_8/A gnd BUFX4_6/Y vdd BUFX4
XDFFPOSX1_255 NAND2X1_632/B CLKBUF1_52/Y DFFPOSX1_255/D gnd vdd DFFPOSX1
XDFFPOSX1_244 INVX1_204/A CLKBUF1_64/Y DFFPOSX1_244/D gnd vdd DFFPOSX1
XDFFPOSX1_233 INVX1_14/A CLKBUF1_10/Y OAI21X1_1553/Y gnd vdd DFFPOSX1
XDFFPOSX1_266 NAND2X1_289/B CLKBUF1_93/Y OAI21X1_1605/Y gnd vdd DFFPOSX1
XDFFPOSX1_277 INVX1_270/A CLKBUF1_89/Y OAI21X1_1622/Y gnd vdd DFFPOSX1
XDFFPOSX1_288 NOR2X1_367/A CLKBUF1_48/Y AOI21X1_293/Y gnd vdd DFFPOSX1
XNAND2X1_303 BUFX4_242/Y NOR2X1_24/A gnd OAI21X1_879/C vdd NAND2X1
XNAND2X1_336 BUFX4_205/Y NOR2X1_212/A gnd OAI21X1_910/C vdd NAND2X1
XNAND2X1_314 BUFX4_262/Y NOR2X1_74/A gnd OAI21X1_889/C vdd NAND2X1
XNAND2X1_325 MUX2X1_5/S NOR2X1_126/A gnd OAI21X1_899/C vdd NAND2X1
XDFFPOSX1_299 NOR2X1_372/A CLKBUF1_39/Y AOI21X1_296/Y gnd vdd DFFPOSX1
XNAND2X1_358 BUFX4_243/Y NAND2X1_358/B gnd NAND2X1_358/Y vdd NAND2X1
XNAND2X1_347 BUFX4_223/Y NOR2X1_314/A gnd NAND2X1_347/Y vdd NAND2X1
XNAND2X1_369 BUFX4_265/Y OAI21X1_157/C gnd OAI21X1_940/C vdd NAND2X1
XFILL_26_8_1 gnd vdd FILL
XFILL_0_3_0 gnd vdd FILL
XFILL_1_8_1 gnd vdd FILL
XFILL_25_3_0 gnd vdd FILL
XNOR2X1_380 NOR2X1_380/A NOR2X1_387/B gnd NOR2X1_380/Y vdd NOR2X1
XOAI21X1_842 INVX1_54/Y BUFX4_268/Y NAND2X1_264/Y gnd MUX2X1_37/A vdd OAI21X1
XOAI21X1_820 INVX1_35/Y BUFX4_230/Y NAND2X1_235/Y gnd NAND2X1_236/B vdd OAI21X1
XOAI21X1_831 INVX1_44/Y BUFX4_248/Y OAI21X1_831/C gnd NAND2X1_254/B vdd OAI21X1
XOAI21X1_864 INVX1_76/Y BUFX4_213/Y NAND2X1_287/Y gnd MUX2X1_53/A vdd OAI21X1
XOAI21X1_875 INVX1_87/Y BUFX4_235/Y OAI21X1_875/C gnd MUX2X1_62/B vdd OAI21X1
XOAI21X1_853 INVX1_65/Y BUFX4_191/Y NAND2X1_276/Y gnd MUX2X1_46/B vdd OAI21X1
XOAI21X1_886 INVX1_98/Y BUFX4_257/Y NAND2X1_311/Y gnd MUX2X1_70/A vdd OAI21X1
XOAI21X1_897 INVX1_109/Y MUX2X1_1/S OAI21X1_897/C gnd MUX2X1_79/B vdd OAI21X1
XMUX2X1_331 MUX2X1_331/A MUX2X1_331/B BUFX4_7/Y gnd MUX2X1_333/B vdd MUX2X1
XMUX2X1_320 MUX2X1_320/A MUX2X1_320/B BUFX4_21/Y gnd MUX2X1_320/Y vdd MUX2X1
XMUX2X1_342 MUX2X1_341/Y MUX2X1_340/Y INVX2_6/A gnd MUX2X1_342/Y vdd MUX2X1
XMUX2X1_375 MUX2X1_375/A MUX2X1_373/Y INVX2_6/A gnd MUX2X1_375/Y vdd MUX2X1
XMUX2X1_353 MUX2X1_353/A MUX2X1_353/B BUFX4_8/Y gnd MUX2X1_354/A vdd MUX2X1
XMUX2X1_364 MUX2X1_364/A MUX2X1_364/B BUFX4_56/Y gnd MUX2X1_364/Y vdd MUX2X1
XFILL_8_4_0 gnd vdd FILL
XNAND2X1_870 INVX8_9/A NOR2X1_378/Y gnd NAND2X1_870/Y vdd NAND2X1
XFILL_16_3_0 gnd vdd FILL
XFILL_17_8_1 gnd vdd FILL
XOAI21X1_105 NOR2X1_21/B INVX2_1/A INVX1_26/A gnd OAI21X1_105/Y vdd OAI21X1
XOAI21X1_138 NAND2X1_18/Y BUFX4_127/Y OAI21X1_137/Y gnd OAI21X1_138/Y vdd OAI21X1
XOAI21X1_116 AOI21X1_6/A NAND2X1_16/Y OAI21X1_115/Y gnd OAI21X1_116/Y vdd OAI21X1
XOAI21X1_127 NOR2X1_52/B BUFX4_178/Y OAI21X1_127/C gnd OAI21X1_128/C vdd OAI21X1
XOAI21X1_149 INVX4_3/A BUFX4_173/Y INVX1_408/A gnd OAI21X1_150/C vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd q[2] vdd BUFX2
XNAND2X1_100 INVX8_11/A INVX1_2/Y gnd OAI21X1_544/B vdd NAND2X1
XNAND2X1_144 BUFX4_144/Y NOR2X1_133/Y gnd NAND2X1_144/Y vdd NAND2X1
XNAND2X1_122 BUFX4_326/Y NOR2X1_101/Y gnd NAND2X1_122/Y vdd NAND2X1
XNAND2X1_111 BUFX4_335/Y NOR2X1_91/Y gnd NAND2X1_111/Y vdd NAND2X1
XNAND2X1_133 BUFX4_137/Y NOR2X1_111/Y gnd OAI21X1_606/C vdd NAND2X1
XNAND2X1_155 BUFX4_448/Y NOR2X1_145/B gnd NAND2X1_155/Y vdd NAND2X1
XNAND2X1_177 INVX8_4/A NOR2X1_177/Y gnd OAI21X1_708/C vdd NAND2X1
XNAND2X1_166 BUFX4_450/Y NOR2X1_166/Y gnd OAI21X1_668/C vdd NAND2X1
XNAND2X1_199 INVX8_11/A INVX2_5/Y gnd OAI21X1_757/B vdd NAND2X1
XNAND2X1_188 BUFX4_139/Y NOR2X1_189/B gnd OAI21X1_719/C vdd NAND2X1
XFILL_41_6_1 gnd vdd FILL
XFILL_40_1_0 gnd vdd FILL
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XOAI21X1_650 BUFX4_153/Y BUFX4_121/Y NAND2X1_672/B gnd OAI21X1_651/C vdd OAI21X1
XOAI21X1_683 BUFX4_462/Y BUFX4_66/Y INVX1_309/A gnd OAI21X1_684/C vdd OAI21X1
XAOI21X1_3 AOI21X1_3/A NOR2X1_2/Y NOR2X1_5/Y gnd AOI21X1_3/Y vdd AOI21X1
XOAI21X1_661 INVX1_115/Y NOR2X1_155/Y OAI21X1_661/C gnd OAI21X1_661/Y vdd OAI21X1
XOAI21X1_672 INVX1_372/Y NOR2X1_166/Y NAND2X1_170/Y gnd OAI21X1_672/Y vdd OAI21X1
XOAI21X1_694 BUFX4_426/Y OAI21X1_704/B OAI21X1_693/Y gnd OAI21X1_694/Y vdd OAI21X1
XMUX2X1_150 MUX2X1_149/Y MUX2X1_150/B MUX2X1_84/S gnd MUX2X1_150/Y vdd MUX2X1
XMUX2X1_183 MUX2X1_182/Y MUX2X1_181/Y MUX2X1_84/S gnd MUX2X1_183/Y vdd MUX2X1
XMUX2X1_161 MUX2X1_161/A MUX2X1_161/B BUFX4_59/Y gnd MUX2X1_162/A vdd MUX2X1
XMUX2X1_172 MUX2X1_172/A MUX2X1_172/B BUFX4_55/Y gnd MUX2X1_174/B vdd MUX2X1
XMUX2X1_194 MUX2X1_194/A MUX2X1_194/B BUFX4_52/Y gnd MUX2X1_195/A vdd MUX2X1
XFILL_48_2_0 gnd vdd FILL
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XFILL_32_6_1 gnd vdd FILL
XFILL_31_1_0 gnd vdd FILL
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XFILL_39_2_0 gnd vdd FILL
XFILL_23_6_1 gnd vdd FILL
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_33 BUFX4_129/Y NOR2X1_43/B NOR2X1_43/Y gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_44 BUFX4_299/Y NOR2X1_55/B NOR2X1_56/Y gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_11 AOI21X1_3/A NOR2X1_14/B NOR2X1_15/Y gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_22 BUFX4_97/Y NOR2X1_27/B NOR2X1_28/Y gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_55 BUFX4_283/Y NOR2X1_67/B NOR2X1_69/Y gnd AOI21X1_55/Y vdd AOI21X1
XAOI21X1_66 BUFX4_425/Y NOR2X1_90/B NOR2X1_84/Y gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_77 BUFX4_396/Y NOR2X1_96/B NOR2X1_97/Y gnd AOI21X1_77/Y vdd AOI21X1
XOAI21X1_6 BUFX4_109/Y NAND2X1_1/Y OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_99 BUFX4_130/Y NOR2X1_126/B NOR2X1_125/Y gnd AOI21X1_99/Y vdd AOI21X1
XAOI21X1_88 BUFX4_372/Y NOR2X1_103/B NOR2X1_110/Y gnd AOI21X1_88/Y vdd AOI21X1
XFILL_6_7_1 gnd vdd FILL
XFILL_5_2_0 gnd vdd FILL
XBUFX4_319 BUFX4_316/A gnd BUFX4_319/Y vdd BUFX4
XBUFX4_308 INVX8_14/Y gnd BUFX4_308/Y vdd BUFX4
XFILL_13_1_0 gnd vdd FILL
XFILL_14_6_1 gnd vdd FILL
XOAI21X1_1209 INVX1_421/Y BUFX4_210/Y NAND2X1_659/Y gnd MUX2X1_313/B vdd OAI21X1
XOAI21X1_480 BUFX4_377/Y NAND2X1_95/Y OAI21X1_479/Y gnd OAI21X1_480/Y vdd OAI21X1
XOAI21X1_491 BUFX4_169/Y BUFX4_340/Y INVX1_360/A gnd OAI21X1_492/C vdd OAI21X1
XINVX1_500 INVX1_500/A gnd INVX1_500/Y vdd INVX1
XBUFX4_105 BUFX4_105/A gnd BUFX4_105/Y vdd BUFX4
XBUFX4_127 INVX8_2/Y gnd BUFX4_127/Y vdd BUFX4
XBUFX4_116 INVX8_4/Y gnd BUFX4_116/Y vdd BUFX4
XFILL_46_5_1 gnd vdd FILL
XBUFX4_149 INVX8_11/Y gnd NOR2X1_72/B vdd BUFX4
XBUFX4_138 d[6] gnd INVX8_8/A vdd BUFX4
XFILL_45_0_0 gnd vdd FILL
XNOR2X1_209 NOR2X1_209/A NOR2X1_206/B gnd NOR2X1_209/Y vdd NOR2X1
XOAI21X1_1006 INVX1_218/Y BUFX4_200/Y NAND2X1_440/Y gnd MUX2X1_160/A vdd OAI21X1
XOAI21X1_1017 INVX1_229/Y BUFX4_222/Y NAND2X1_452/Y gnd MUX2X1_169/B vdd OAI21X1
XOAI21X1_1028 INVX1_240/Y BUFX4_244/Y NAND2X1_464/Y gnd MUX2X1_176/A vdd OAI21X1
XDFFPOSX1_607 NAND2X1_656/B CLKBUF1_70/Y OAI21X1_342/Y gnd vdd DFFPOSX1
XDFFPOSX1_618 NAND2X1_312/B CLKBUF1_79/Y OAI21X1_364/Y gnd vdd DFFPOSX1
XDFFPOSX1_629 INVX1_292/A CLKBUF1_6/Y OAI21X1_386/Y gnd vdd DFFPOSX1
XOAI21X1_1039 INVX1_251/Y BUFX4_266/Y NAND2X1_475/Y gnd MUX2X1_185/B vdd OAI21X1
XINVX1_330 INVX1_330/A gnd INVX1_330/Y vdd INVX1
XINVX1_341 INVX1_341/A gnd INVX1_341/Y vdd INVX1
XINVX1_352 INVX1_352/A gnd INVX1_352/Y vdd INVX1
XINVX1_396 INVX1_396/A gnd INVX1_396/Y vdd INVX1
XINVX1_374 INVX1_374/A gnd INVX1_374/Y vdd INVX1
XINVX1_363 INVX1_363/A gnd INVX1_363/Y vdd INVX1
XINVX1_385 INVX1_385/A gnd INVX1_385/Y vdd INVX1
XFILL_37_5_1 gnd vdd FILL
XFILL_36_0_0 gnd vdd FILL
XFILL_20_4_1 gnd vdd FILL
XAOI21X1_301 BUFX4_376/Y NOR2X1_373/B NOR2X1_377/Y gnd AOI21X1_301/Y vdd AOI21X1
XDFFPOSX1_11 NOR2X1_258/A CLKBUF1_5/Y AOI21X1_209/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 NOR2X1_269/A CLKBUF1_14/Y DFFPOSX1_44/D gnd vdd DFFPOSX1
XOAI21X1_1540 NAND2X1_837/Y BUFX4_424/Y OAI21X1_1540/C gnd DFFPOSX1_226/D vdd OAI21X1
XDFFPOSX1_22 NOR2X1_281/A CLKBUF1_56/Y DFFPOSX1_22/D gnd vdd DFFPOSX1
XDFFPOSX1_33 INVX1_35/A CLKBUF1_44/Y DFFPOSX1_33/D gnd vdd DFFPOSX1
XDFFPOSX1_77 NAND2X1_483/B CLKBUF1_43/Y DFFPOSX1_77/D gnd vdd DFFPOSX1
XOAI21X1_1562 BUFX4_171/Y INVX2_9/A INVX1_268/A gnd OAI21X1_1562/Y vdd OAI21X1
XOAI21X1_1584 BUFX4_410/Y BUFX4_93/Y NAND2X1_701/B gnd OAI21X1_1585/C vdd OAI21X1
XOAI21X1_1573 BUFX4_424/Y NAND2X1_840/Y OAI21X1_1573/C gnd DFFPOSX1_250/D vdd OAI21X1
XOAI21X1_1551 BUFX4_312/Y BUFX4_95/Y INVX1_459/A gnd OAI21X1_1551/Y vdd OAI21X1
XDFFPOSX1_55 INVX1_384/A CLKBUF1_56/Y DFFPOSX1_55/D gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX1_65/A CLKBUF1_43/Y DFFPOSX1_66/D gnd vdd DFFPOSX1
XDFFPOSX1_99 INVX1_131/A CLKBUF1_12/Y DFFPOSX1_99/D gnd vdd DFFPOSX1
XOAI21X1_1595 BUFX4_399/Y NAND2X1_842/Y OAI21X1_1595/C gnd OAI21X1_1595/Y vdd OAI21X1
XDFFPOSX1_88 INVX1_450/A CLKBUF1_53/Y DFFPOSX1_88/D gnd vdd DFFPOSX1
XFILL_28_5_1 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XFILL_11_4_1 gnd vdd FILL
XFILL_19_5_1 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XDFFPOSX1_404 INVX1_214/A CLKBUF1_26/Y OAI21X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_415 NAND2X1_643/B CLKBUF1_49/Y OAI21X1_102/Y gnd vdd DFFPOSX1
XDFFPOSX1_426 NAND2X1_299/B CLKBUF1_49/Y OAI21X1_124/Y gnd vdd DFFPOSX1
XDFFPOSX1_437 INVX1_280/A CLKBUF1_27/Y OAI21X1_146/Y gnd vdd DFFPOSX1
XDFFPOSX1_459 OAI21X1_189/C CLKBUF1_5/Y OAI21X1_190/Y gnd vdd DFFPOSX1
XDFFPOSX1_448 NAND2X1_714/B CLKBUF1_72/Y OAI21X1_168/Y gnd vdd DFFPOSX1
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XNAND2X1_518 BUFX4_244/Y NAND2X1_518/B gnd NAND2X1_518/Y vdd NAND2X1
XINVX1_182 INVX1_182/A gnd INVX1_182/Y vdd INVX1
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XNAND2X1_507 BUFX4_224/Y NAND2X1_507/B gnd NAND2X1_507/Y vdd NAND2X1
XNAND2X1_529 AOI22X1_45/Y AOI22X1_46/Y gnd AOI22X1_49/A vdd NAND2X1
XAOI21X1_120 BUFX4_299/Y NOR2X1_153/B NOR2X1_150/Y gnd AOI21X1_120/Y vdd AOI21X1
XAOI21X1_131 BUFX4_104/Y NOR2X1_158/B NOR2X1_163/Y gnd AOI21X1_131/Y vdd AOI21X1
XAOI21X1_142 BUFX4_372/Y NOR2X1_173/B NOR2X1_176/Y gnd AOI21X1_142/Y vdd AOI21X1
XAOI21X1_164 BUFX4_115/Y NOR2X1_206/B NOR2X1_204/Y gnd AOI21X1_164/Y vdd AOI21X1
XAOI21X1_153 BUFX4_131/Y NOR2X1_197/B NOR2X1_191/Y gnd AOI21X1_153/Y vdd AOI21X1
XAOI21X1_175 BUFX4_103/Y NOR2X1_216/B NOR2X1_216/Y gnd AOI21X1_175/Y vdd AOI21X1
XAOI21X1_186 BUFX4_123/Y NOR2X1_228/Y NOR2X1_229/Y gnd AOI21X1_186/Y vdd AOI21X1
XAOI21X1_197 INVX8_1/Y INVX1_21/Y OR2X2_1/A gnd OAI21X1_806/C vdd AOI21X1
XOAI21X1_1381 BUFX4_167/Y BUFX4_465/Y INVX1_132/A gnd OAI21X1_1382/C vdd OAI21X1
XOAI21X1_1392 NAND2X1_811/Y BUFX4_373/Y OAI21X1_1392/C gnd DFFPOSX1_120/D vdd OAI21X1
XDFFPOSX1_960 NOR2X1_209/A CLKBUF1_87/Y AOI21X1_169/Y gnd vdd DFFPOSX1
XOAI21X1_1370 INVX1_67/Y NOR2X1_309/Y NAND2X1_803/Y gnd DFFPOSX1_98/D vdd OAI21X1
XDFFPOSX1_993 MUX2X1_25/B CLKBUF1_97/Y OAI21X1_777/Y gnd vdd DFFPOSX1
XDFFPOSX1_971 NAND2X1_404/B CLKBUF1_67/Y OAI21X1_749/Y gnd vdd DFFPOSX1
XDFFPOSX1_982 INVX1_378/A CLKBUF1_59/Y OAI21X1_771/Y gnd vdd DFFPOSX1
XFILL_43_3_1 gnd vdd FILL
XFILL_34_3_1 gnd vdd FILL
XFILL_13_1 gnd vdd FILL
XOAI21X1_309 INVX1_289/Y NOR2X1_61/Y NAND2X1_73/Y gnd OAI21X1_309/Y vdd OAI21X1
XDFFPOSX1_212 INVX1_202/A CLKBUF1_76/Y OAI21X1_1528/Y gnd vdd DFFPOSX1
XDFFPOSX1_201 MUX2X1_29/A CLKBUF1_36/Y OAI21X1_1506/Y gnd vdd DFFPOSX1
XBUFX4_7 BUFX4_8/A gnd BUFX4_7/Y vdd BUFX4
XDFFPOSX1_234 NOR2X1_351/A CLKBUF1_66/Y AOI21X1_279/Y gnd vdd DFFPOSX1
XDFFPOSX1_245 INVX1_268/A CLKBUF1_66/Y OAI21X1_1563/Y gnd vdd DFFPOSX1
XDFFPOSX1_223 NOR2X1_348/A CLKBUF1_35/Y AOI21X1_277/Y gnd vdd DFFPOSX1
XDFFPOSX1_256 NAND2X1_701/B CLKBUF1_64/Y DFFPOSX1_256/D gnd vdd DFFPOSX1
XDFFPOSX1_267 NAND2X1_358/B CLKBUF1_12/Y OAI21X1_1607/Y gnd vdd DFFPOSX1
XDFFPOSX1_289 INVX1_18/A CLKBUF1_63/Y OAI21X1_1626/Y gnd vdd DFFPOSX1
XDFFPOSX1_278 INVX1_334/A CLKBUF1_75/Y DFFPOSX1_278/D gnd vdd DFFPOSX1
XNAND2X1_326 MUX2X1_9/S NOR2X1_137/A gnd NAND2X1_326/Y vdd NAND2X1
XNAND2X1_315 BUFX4_264/Y NAND2X1_315/B gnd OAI21X1_890/C vdd NAND2X1
XNAND2X1_304 BUFX4_244/Y NOR2X1_34/A gnd OAI21X1_880/C vdd NAND2X1
XNAND2X1_337 BUFX4_207/Y NOR2X1_221/A gnd OAI21X1_911/C vdd NAND2X1
XNAND2X1_359 BUFX4_245/Y NOR2X1_362/A gnd NAND2X1_359/Y vdd NAND2X1
XNAND2X1_348 BUFX4_225/Y NAND2X1_348/B gnd NAND2X1_348/Y vdd NAND2X1
XFILL_25_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XNOR2X1_370 NOR2X1_370/A NOR2X1_373/B gnd NOR2X1_370/Y vdd NOR2X1
XNOR2X1_381 NOR2X1_381/A NOR2X1_387/B gnd NOR2X1_381/Y vdd NOR2X1
XOAI21X1_821 INVX1_36/Y BUFX4_232/Y OAI21X1_821/C gnd NAND2X1_238/B vdd OAI21X1
XOAI21X1_810 INVX8_1/Y OAI21X1_153/C OAI21X1_810/C gnd NAND3X1_3/A vdd OAI21X1
XOAI21X1_832 OAI21X1_832/A OAI21X1_832/B BUFX4_321/Y gnd NAND3X1_5/C vdd OAI21X1
XOAI21X1_843 INVX1_55/Y BUFX4_270/Y NAND2X1_265/Y gnd MUX2X1_38/B vdd OAI21X1
XOAI21X1_865 INVX1_77/Y BUFX4_215/Y OAI21X1_865/C gnd MUX2X1_55/B vdd OAI21X1
XOAI21X1_876 INVX1_88/Y BUFX4_237/Y NAND2X1_300/Y gnd MUX2X1_62/A vdd OAI21X1
XOAI21X1_854 INVX1_66/Y BUFX4_193/Y OAI21X1_854/C gnd MUX2X1_46/A vdd OAI21X1
XOAI21X1_887 INVX1_99/Y BUFX4_259/Y NAND2X1_312/Y gnd MUX2X1_71/B vdd OAI21X1
XOAI21X1_898 INVX1_110/Y MUX2X1_4/S NAND2X1_324/Y gnd MUX2X1_79/A vdd OAI21X1
XMUX2X1_310 MUX2X1_310/A MUX2X1_310/B BUFX4_37/Y gnd MUX2X1_312/B vdd MUX2X1
XMUX2X1_332 MUX2X1_332/A MUX2X1_332/B BUFX4_38/Y gnd MUX2X1_333/A vdd MUX2X1
XMUX2X1_321 MUX2X1_320/Y MUX2X1_321/B BUFX4_363/Y gnd AOI22X1_67/A vdd MUX2X1
XMUX2X1_354 MUX2X1_354/A MUX2X1_352/Y BUFX4_363/Y gnd AOI22X1_73/D vdd MUX2X1
XMUX2X1_343 MUX2X1_343/A MUX2X1_343/B BUFX4_22/Y gnd MUX2X1_345/B vdd MUX2X1
XMUX2X1_365 MUX2X1_365/A MUX2X1_365/B BUFX4_19/Y gnd MUX2X1_365/Y vdd MUX2X1
XMUX2X1_376 MUX2X1_376/A MUX2X1_376/B BUFX4_5/Y gnd MUX2X1_376/Y vdd MUX2X1
XDFFPOSX1_790 INVX1_366/A CLKBUF1_92/Y OAI21X1_605/Y gnd vdd DFFPOSX1
XFILL_8_4_1 gnd vdd FILL
XNAND2X1_871 INVX2_11/Y INVX8_12/A gnd NAND2X1_871/Y vdd NAND2X1
XNAND2X1_860 INVX2_10/Y INVX4_3/Y gnd NAND2X1_860/Y vdd NAND2X1
XFILL_16_3_1 gnd vdd FILL
XOAI21X1_106 BUFX4_127/Y NAND2X1_16/Y OAI21X1_105/Y gnd OAI21X1_106/Y vdd OAI21X1
XOAI21X1_117 NOR2X1_51/B BUFX4_179/Y INVX1_407/A gnd OAI21X1_118/C vdd OAI21X1
XOAI21X1_128 BUFX4_297/Y NAND2X1_17/Y OAI21X1_128/C gnd OAI21X1_128/Y vdd OAI21X1
XOAI21X1_139 INVX4_3/A BUFX4_173/Y INVX1_88/A gnd OAI21X1_139/Y vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd q[3] vdd BUFX2
XNAND2X1_101 INVX8_2/A NOR2X1_81/Y gnd OAI21X1_545/C vdd NAND2X1
XNAND2X1_123 BUFX4_136/Y NOR2X1_101/Y gnd NAND2X1_123/Y vdd NAND2X1
XNAND2X1_112 BUFX4_145/Y NOR2X1_91/Y gnd OAI21X1_556/C vdd NAND2X1
XNAND2X1_134 BUFX4_428/Y NOR2X1_111/Y gnd OAI21X1_607/C vdd NAND2X1
XNAND2X1_167 BUFX4_332/Y NOR2X1_166/Y gnd NAND2X1_167/Y vdd NAND2X1
XNAND2X1_145 BUFX4_447/Y NOR2X1_133/Y gnd OAI21X1_618/C vdd NAND2X1
XNAND2X1_178 INVX8_5/A NOR2X1_177/Y gnd OAI21X1_709/C vdd NAND2X1
XNAND2X1_156 BUFX4_330/Y NOR2X1_145/B gnd NAND2X1_156/Y vdd NAND2X1
XNAND2X1_189 BUFX4_430/Y NOR2X1_189/B gnd OAI21X1_720/C vdd NAND2X1
XFILL_40_1_1 gnd vdd FILL
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XOAI21X1_651 BUFX4_287/Y OAI21X1_651/B OAI21X1_651/C gnd OAI21X1_651/Y vdd OAI21X1
XOAI21X1_640 BUFX4_153/Y INVX1_4/A NAND2X1_327/B gnd OAI21X1_640/Y vdd OAI21X1
XOAI21X1_662 INVX1_179/Y NOR2X1_155/Y OAI21X1_662/C gnd OAI21X1_662/Y vdd OAI21X1
XOAI21X1_684 BUFX4_402/Y NAND2X1_174/Y OAI21X1_684/C gnd OAI21X1_684/Y vdd OAI21X1
XAOI21X1_4 BUFX4_298/Y NOR2X1_2/Y NOR2X1_6/Y gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_673 INVX1_436/Y NOR2X1_166/Y NAND2X1_171/Y gnd OAI21X1_673/Y vdd OAI21X1
XOAI21X1_695 BUFX4_146/Y INVX1_5/A NAND2X1_400/B gnd OAI21X1_695/Y vdd OAI21X1
XMUX2X1_140 MUX2X1_140/A MUX2X1_140/B BUFX4_21/Y gnd MUX2X1_140/Y vdd MUX2X1
XMUX2X1_162 MUX2X1_162/A MUX2X1_160/Y MUX2X1_96/S gnd MUX2X1_162/Y vdd MUX2X1
XMUX2X1_151 MUX2X1_151/A MUX2X1_151/B BUFX4_7/Y gnd MUX2X1_153/B vdd MUX2X1
XMUX2X1_173 MUX2X1_173/A MUX2X1_173/B BUFX4_8/Y gnd MUX2X1_174/A vdd MUX2X1
XMUX2X1_184 MUX2X1_184/A MUX2X1_184/B BUFX4_56/Y gnd MUX2X1_186/B vdd MUX2X1
XMUX2X1_195 MUX2X1_195/A MUX2X1_195/B MUX2X1_96/S gnd AOI22X1_41/A vdd MUX2X1
XFILL_48_2_1 gnd vdd FILL
XNAND2X1_690 BUFX4_265/Y NAND2X1_690/B gnd NAND2X1_690/Y vdd NAND2X1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XFILL_31_1_1 gnd vdd FILL
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XFILL_39_2_1 gnd vdd FILL
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_34 BUFX4_422/Y NOR2X1_43/B NOR2X1_44/Y gnd AOI21X1_34/Y vdd AOI21X1
XAOI21X1_12 BUFX4_304/Y NOR2X1_14/B NOR2X1_16/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_23 BUFX4_285/Y NOR2X1_27/B NOR2X1_29/Y gnd AOI21X1_23/Y vdd AOI21X1
XAOI21X1_56 BUFX4_377/Y NOR2X1_67/B NOR2X1_70/Y gnd AOI21X1_56/Y vdd AOI21X1
XAOI21X1_67 BUFX4_110/Y NOR2X1_90/B NOR2X1_85/Y gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_45 BUFX4_394/Y NOR2X1_55/B NOR2X1_57/Y gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_89 BUFX4_130/Y NOR2X1_111/Y NOR2X1_112/Y gnd AOI21X1_89/Y vdd AOI21X1
XAOI21X1_78 BUFX4_104/Y NOR2X1_96/B NOR2X1_98/Y gnd AOI21X1_78/Y vdd AOI21X1
XOAI21X1_7 BUFX4_307/Y OAI21X1_7/B INVX1_211/A gnd OAI21X1_7/Y vdd OAI21X1
XFILL_5_2_1 gnd vdd FILL
XBUFX4_309 INVX8_14/Y gnd NOR2X1_51/B vdd BUFX4
XFILL_13_1_1 gnd vdd FILL
XOAI21X1_470 BUFX4_109/Y NAND2X1_95/Y OAI21X1_470/C gnd OAI21X1_470/Y vdd OAI21X1
XINVX1_501 INVX1_501/A gnd INVX1_501/Y vdd INVX1
XOAI21X1_492 NAND2X1_96/Y BUFX4_101/Y OAI21X1_492/C gnd OAI21X1_492/Y vdd OAI21X1
XOAI21X1_481 BUFX4_169/Y BUFX4_336/Y INVX1_56/A gnd OAI21X1_482/C vdd OAI21X1
XOAI21X1_1700 BUFX4_85/Y OAI21X1_5/B NAND2X1_570/B gnd OAI21X1_1701/C vdd OAI21X1
XBUFX4_128 INVX8_2/Y gnd BUFX4_128/Y vdd BUFX4
XBUFX4_117 INVX8_4/Y gnd BUFX4_117/Y vdd BUFX4
XBUFX4_106 BUFX4_105/A gnd INVX1_3/A vdd BUFX4
XBUFX4_139 d[6] gnd BUFX4_139/Y vdd BUFX4
XFILL_45_0_1 gnd vdd FILL
XOAI21X1_1018 INVX1_230/Y BUFX4_224/Y NAND2X1_453/Y gnd MUX2X1_169/A vdd OAI21X1
XOAI21X1_1007 INVX1_219/Y BUFX4_202/Y NAND2X1_441/Y gnd MUX2X1_161/B vdd OAI21X1
XOAI21X1_1029 INVX1_241/Y BUFX4_246/Y NAND2X1_465/Y gnd MUX2X1_178/B vdd OAI21X1
XDFFPOSX1_619 NAND2X1_381/B CLKBUF1_34/Y OAI21X1_366/Y gnd vdd DFFPOSX1
XDFFPOSX1_608 NAND2X1_725/B CLKBUF1_69/Y OAI21X1_344/Y gnd vdd DFFPOSX1
XINVX1_331 INVX1_331/A gnd INVX1_331/Y vdd INVX1
XINVX1_320 INVX1_320/A gnd INVX1_320/Y vdd INVX1
XINVX1_353 INVX1_353/A gnd INVX1_353/Y vdd INVX1
XINVX1_342 INVX1_342/A gnd INVX1_342/Y vdd INVX1
XINVX1_375 INVX1_375/A gnd INVX1_375/Y vdd INVX1
XINVX1_364 INVX1_364/A gnd INVX1_364/Y vdd INVX1
XINVX1_386 INVX1_386/A gnd INVX1_386/Y vdd INVX1
XINVX1_397 INVX1_397/A gnd INVX1_397/Y vdd INVX1
XFILL_1_1 gnd vdd FILL
XFILL_36_0_1 gnd vdd FILL
XFILL_43_1 gnd vdd FILL
XAOI21X1_302 BUFX4_123/Y NOR2X1_387/B NOR2X1_380/Y gnd AOI21X1_302/Y vdd AOI21X1
XOAI21X1_1541 NOR2X1_21/B INVX2_9/A INVX1_139/A gnd OAI21X1_1542/C vdd OAI21X1
XOAI21X1_1530 NAND2X1_836/Y BUFX4_402/Y OAI21X1_1530/C gnd DFFPOSX1_213/D vdd OAI21X1
XDFFPOSX1_45 NOR2X1_270/A CLKBUF1_21/Y AOI21X1_219/Y gnd vdd DFFPOSX1
XDFFPOSX1_12 NOR2X1_259/A CLKBUF1_14/Y AOI21X1_210/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 NOR2X1_282/A CLKBUF1_50/Y DFFPOSX1_23/D gnd vdd DFFPOSX1
XDFFPOSX1_34 INVX1_63/A CLKBUF1_50/Y DFFPOSX1_34/D gnd vdd DFFPOSX1
XDFFPOSX1_67 INVX1_129/A CLKBUF1_84/Y DFFPOSX1_67/D gnd vdd DFFPOSX1
XOAI21X1_1574 BUFX4_410/Y INVX2_9/A NAND2X1_356/B gnd OAI21X1_1575/C vdd OAI21X1
XOAI21X1_1563 NAND2X1_839/Y BUFX4_398/Y OAI21X1_1562/Y gnd OAI21X1_1563/Y vdd OAI21X1
XOAI21X1_1552 NAND2X1_837/Y BUFX4_380/Y OAI21X1_1551/Y gnd DFFPOSX1_232/D vdd OAI21X1
XDFFPOSX1_56 INVX1_448/A CLKBUF1_40/Y DFFPOSX1_56/D gnd vdd DFFPOSX1
XDFFPOSX1_78 NAND2X1_552/B CLKBUF1_17/Y DFFPOSX1_78/D gnd vdd DFFPOSX1
XDFFPOSX1_89 NOR2X1_300/A CLKBUF1_42/Y AOI21X1_239/Y gnd vdd DFFPOSX1
XOAI21X1_1585 BUFX4_380/Y NAND2X1_840/Y OAI21X1_1585/C gnd DFFPOSX1_256/D vdd OAI21X1
XOAI21X1_1596 BUFX4_454/Y BUFX4_348/Y INVX1_333/A gnd OAI21X1_1596/Y vdd OAI21X1
XFILL_2_0_1 gnd vdd FILL
XFILL_27_0_1 gnd vdd FILL
XFILL_47_8_0 gnd vdd FILL
XFILL_18_0_1 gnd vdd FILL
XFILL_30_7_0 gnd vdd FILL
XDFFPOSX1_416 NAND2X1_712/B CLKBUF1_94/Y OAI21X1_104/Y gnd vdd DFFPOSX1
XDFFPOSX1_405 INVX1_278/A CLKBUF1_75/Y OAI21X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_438 INVX1_344/A CLKBUF1_41/Y OAI21X1_148/Y gnd vdd DFFPOSX1
XDFFPOSX1_427 NAND2X1_368/B CLKBUF1_41/Y OAI21X1_126/Y gnd vdd DFFPOSX1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XDFFPOSX1_449 INVX1_32/A CLKBUF1_71/Y OAI21X1_170/Y gnd vdd DFFPOSX1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XINVX1_194 INVX1_194/A gnd INVX1_194/Y vdd INVX1
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XNAND2X1_508 BUFX4_226/Y NAND2X1_508/B gnd NAND2X1_508/Y vdd NAND2X1
XINVX1_172 INVX1_172/A gnd INVX1_172/Y vdd INVX1
XNAND2X1_519 BUFX4_246/Y NAND2X1_519/B gnd NAND2X1_519/Y vdd NAND2X1
XFILL_38_8_0 gnd vdd FILL
XFILL_21_7_0 gnd vdd FILL
XAOI21X1_132 BUFX4_287/Y NOR2X1_158/B NOR2X1_164/Y gnd AOI21X1_132/Y vdd AOI21X1
XAOI21X1_121 BUFX4_396/Y NOR2X1_153/B NOR2X1_151/Y gnd AOI21X1_121/Y vdd AOI21X1
XAOI21X1_110 BUFX4_117/Y NOR2X1_139/B NOR2X1_138/Y gnd AOI21X1_110/Y vdd AOI21X1
XAOI21X1_154 BUFX4_426/Y NOR2X1_197/B NOR2X1_192/Y gnd AOI21X1_154/Y vdd AOI21X1
XAOI21X1_165 BUFX4_301/Y NOR2X1_206/B NOR2X1_205/Y gnd AOI21X1_165/Y vdd AOI21X1
XAOI21X1_143 BUFX4_131/Y NOR2X1_177/Y NOR2X1_178/Y gnd AOI21X1_143/Y vdd AOI21X1
XAOI21X1_176 BUFX4_281/Y NOR2X1_216/B NOR2X1_217/Y gnd AOI21X1_176/Y vdd AOI21X1
XAOI21X1_187 BUFX4_123/Y NOR2X1_236/B NOR2X1_231/Y gnd AOI21X1_187/Y vdd AOI21X1
XAOI21X1_198 INVX8_1/Y INVX1_25/Y OR2X2_1/A gnd OAI21X1_810/C vdd AOI21X1
XOAI21X1_1360 BUFX4_373/Y NAND2X1_793/Y OAI21X1_1359/Y gnd DFFPOSX1_80/D vdd OAI21X1
XOAI21X1_1382 NAND2X1_811/Y BUFX4_112/Y OAI21X1_1382/C gnd OAI21X1_1382/Y vdd OAI21X1
XDFFPOSX1_950 INVX1_376/A CLKBUF1_14/Y OAI21X1_725/Y gnd vdd DFFPOSX1
XOAI21X1_1371 INVX1_131/Y NOR2X1_309/Y NAND2X1_804/Y gnd DFFPOSX1_99/D vdd OAI21X1
XDFFPOSX1_994 INVX1_123/A CLKBUF1_73/Y OAI21X1_779/Y gnd vdd DFFPOSX1
XDFFPOSX1_972 NAND2X1_473/B CLKBUF1_67/Y OAI21X1_751/Y gnd vdd DFFPOSX1
XDFFPOSX1_983 INVX1_442/A CLKBUF1_67/Y OAI21X1_773/Y gnd vdd DFFPOSX1
XDFFPOSX1_961 MUX2X1_22/B CLKBUF1_88/Y OAI21X1_729/Y gnd vdd DFFPOSX1
XOAI21X1_1393 BUFX4_416/Y BUFX4_463/Y NAND2X1_245/B gnd OAI21X1_1393/Y vdd OAI21X1
XFILL_29_8_0 gnd vdd FILL
XFILL_4_8_0 gnd vdd FILL
XFILL_12_7_0 gnd vdd FILL
XDFFPOSX1_213 INVX1_266/A CLKBUF1_76/Y DFFPOSX1_213/D gnd vdd DFFPOSX1
XDFFPOSX1_202 NAND2X1_284/B CLKBUF1_35/Y DFFPOSX1_202/D gnd vdd DFFPOSX1
XDFFPOSX1_246 INVX1_332/A CLKBUF1_64/Y DFFPOSX1_246/D gnd vdd DFFPOSX1
XDFFPOSX1_224 NOR2X1_349/A CLKBUF1_36/Y AOI21X1_278/Y gnd vdd DFFPOSX1
XDFFPOSX1_235 NOR2X1_352/A CLKBUF1_10/Y AOI21X1_280/Y gnd vdd DFFPOSX1
XBUFX4_8 BUFX4_8/A gnd BUFX4_8/Y vdd BUFX4
XDFFPOSX1_279 INVX1_398/A CLKBUF1_89/Y OAI21X1_1624/Y gnd vdd DFFPOSX1
XDFFPOSX1_268 NAND2X1_427/B CLKBUF1_49/Y DFFPOSX1_268/D gnd vdd DFFPOSX1
XDFFPOSX1_257 INVX1_20/A CLKBUF1_25/Y DFFPOSX1_257/D gnd vdd DFFPOSX1
XNAND2X1_316 BUFX4_266/Y NAND2X1_316/B gnd NAND2X1_316/Y vdd NAND2X1
XNAND2X1_305 AOI22X1_12/Y AOI22X1_13/Y gnd AOI22X1_14/D vdd NAND2X1
XNAND2X1_327 MUX2X1_12/S NAND2X1_327/B gnd OAI21X1_901/C vdd NAND2X1
XNAND2X1_338 BUFX4_209/Y NOR2X1_232/A gnd NAND2X1_338/Y vdd NAND2X1
XNAND2X1_349 BUFX4_227/Y NAND2X1_349/B gnd NAND2X1_349/Y vdd NAND2X1
XNOR2X1_360 NOR2X1_360/A NOR2X1_367/B gnd NOR2X1_360/Y vdd NOR2X1
XNOR2X1_382 NOR2X1_382/A NOR2X1_387/B gnd NOR2X1_382/Y vdd NOR2X1
XNOR2X1_371 NOR2X1_371/A NOR2X1_373/B gnd NOR2X1_371/Y vdd NOR2X1
XOAI21X1_800 NOR2X1_275/B INVX1_14/Y OAI21X1_800/C gnd NOR2X1_246/A vdd OAI21X1
XOAI21X1_833 INVX1_45/Y BUFX4_250/Y OAI21X1_833/C gnd MUX2X1_31/B vdd OAI21X1
XOAI21X1_822 AOI21X1_201/Y OAI21X1_822/B BUFX4_354/Y gnd NAND3X1_5/A vdd OAI21X1
XOAI21X1_811 INVX1_26/Y BUFX4_214/Y OAI21X1_811/C gnd NAND2X1_223/B vdd OAI21X1
XOAI21X1_844 INVX1_56/Y BUFX4_272/Y NAND2X1_266/Y gnd MUX2X1_38/A vdd OAI21X1
XOAI21X1_866 INVX1_78/Y BUFX4_217/Y OAI21X1_866/C gnd MUX2X1_55/A vdd OAI21X1
XOAI21X1_855 INVX1_67/Y BUFX4_195/Y OAI21X1_855/C gnd MUX2X1_47/B vdd OAI21X1
XOAI21X1_888 INVX1_100/Y BUFX4_261/Y NAND2X1_313/Y gnd MUX2X1_71/A vdd OAI21X1
XOAI21X1_877 INVX1_89/Y BUFX4_239/Y NAND2X1_301/Y gnd MUX2X1_64/B vdd OAI21X1
XOAI21X1_899 INVX1_111/Y MUX2X1_8/S OAI21X1_899/C gnd MUX2X1_80/B vdd OAI21X1
XMUX2X1_322 MUX2X1_322/A MUX2X1_322/B BUFX4_46/Y gnd MUX2X1_324/B vdd MUX2X1
XMUX2X1_311 MUX2X1_311/A MUX2X1_311/B INVX4_1/A gnd MUX2X1_311/Y vdd MUX2X1
XMUX2X1_300 MUX2X1_299/Y MUX2X1_298/Y MUX2X1_69/S gnd MUX2X1_300/Y vdd MUX2X1
XOAI21X1_1190 INVX1_402/Y BUFX4_271/Y NAND2X1_639/Y gnd MUX2X1_298/A vdd OAI21X1
XMUX2X1_333 MUX2X1_333/A MUX2X1_333/B MUX2X1_69/S gnd MUX2X1_333/Y vdd MUX2X1
XMUX2X1_355 MUX2X1_355/A MUX2X1_355/B BUFX4_39/Y gnd MUX2X1_355/Y vdd MUX2X1
XMUX2X1_344 MUX2X1_344/A MUX2X1_344/B BUFX4_47/Y gnd MUX2X1_345/A vdd MUX2X1
XMUX2X1_366 MUX2X1_365/Y MUX2X1_364/Y MUX2X1_69/S gnd AOI22X1_76/D vdd MUX2X1
XMUX2X1_377 MUX2X1_377/A MUX2X1_377/B BUFX4_36/Y gnd MUX2X1_377/Y vdd MUX2X1
XDFFPOSX1_780 NAND2X1_461/B CLKBUF1_26/Y OAI21X1_592/Y gnd vdd DFFPOSX1
XDFFPOSX1_791 INVX1_430/A CLKBUF1_82/Y OAI21X1_606/Y gnd vdd DFFPOSX1
XNAND2X1_872 INVX2_11/Y INVX8_13/A gnd NAND2X1_872/Y vdd NAND2X1
XNAND2X1_850 BUFX4_136/Y NOR2X1_358/Y gnd NAND2X1_850/Y vdd NAND2X1
XNAND2X1_861 INVX8_16/A INVX2_10/Y gnd NAND2X1_861/Y vdd NAND2X1
XFILL_44_6_0 gnd vdd FILL
XFILL_35_6_0 gnd vdd FILL
XOAI21X1_118 BUFX4_280/Y NAND2X1_16/Y OAI21X1_118/C gnd OAI21X1_118/Y vdd OAI21X1
XOAI21X1_107 NOR2X1_51/B BUFX4_175/Y INVX1_87/A gnd OAI21X1_108/C vdd OAI21X1
XOAI21X1_129 BUFX4_371/Y BUFX4_179/Y NAND2X1_506/B gnd OAI21X1_130/C vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd q[4] vdd BUFX2
XNAND2X1_102 BUFX4_452/Y NOR2X1_81/Y gnd NAND2X1_102/Y vdd NAND2X1
XNAND2X1_135 INVX8_3/A NOR2X1_122/Y gnd OAI21X1_608/C vdd NAND2X1
XNAND2X1_113 BUFX4_448/Y NOR2X1_91/Y gnd OAI21X1_557/C vdd NAND2X1
XNAND2X1_124 BUFX4_427/Y NOR2X1_101/Y gnd OAI21X1_568/C vdd NAND2X1
XNAND2X1_168 BUFX4_142/Y NOR2X1_166/Y gnd NAND2X1_168/Y vdd NAND2X1
XNAND2X1_146 BUFX4_329/Y NOR2X1_133/Y gnd OAI21X1_619/C vdd NAND2X1
XNAND2X1_157 BUFX4_140/Y NOR2X1_145/B gnd NAND2X1_157/Y vdd NAND2X1
XNAND2X1_179 INVX8_6/A NOR2X1_177/Y gnd OAI21X1_710/C vdd NAND2X1
XFILL_26_6_0 gnd vdd FILL
XFILL_1_6_0 gnd vdd FILL
XNOR2X1_190 BUFX4_64/Y NOR2X1_22/B gnd NOR2X1_197/B vdd NOR2X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XOAI21X1_630 BUFX4_456/Y BUFX4_121/Y INVX1_305/A gnd OAI21X1_631/C vdd OAI21X1
XOAI21X1_641 BUFX4_418/Y OAI21X1_651/B OAI21X1_640/Y gnd OAI21X1_641/Y vdd OAI21X1
XOAI21X1_652 BUFX4_153/Y BUFX4_120/Y NAND2X1_741/B gnd OAI21X1_653/C vdd OAI21X1
XOAI21X1_663 INVX1_243/Y NOR2X1_155/Y OAI21X1_663/C gnd OAI21X1_663/Y vdd OAI21X1
XAOI21X1_5 BUFX4_399/Y NOR2X1_2/Y NOR2X1_7/Y gnd AOI21X1_5/Y vdd AOI21X1
XOAI21X1_674 INVX1_500/Y NOR2X1_166/Y NAND2X1_172/Y gnd OAI21X1_674/Y vdd OAI21X1
XOAI21X1_685 BUFX4_462/Y INVX1_5/A INVX1_373/A gnd OAI21X1_685/Y vdd OAI21X1
XOAI21X1_696 BUFX4_115/Y OAI21X1_704/B OAI21X1_695/Y gnd OAI21X1_696/Y vdd OAI21X1
XMUX2X1_141 MUX2X1_140/Y MUX2X1_139/Y MUX2X1_42/S gnd MUX2X1_141/Y vdd MUX2X1
XMUX2X1_130 MUX2X1_130/A MUX2X1_130/B BUFX4_37/Y gnd MUX2X1_130/Y vdd MUX2X1
XMUX2X1_174 MUX2X1_174/A MUX2X1_174/B MUX2X1_42/S gnd AOI22X1_36/D vdd MUX2X1
XMUX2X1_152 MUX2X1_152/A MUX2X1_152/B BUFX4_38/Y gnd MUX2X1_153/A vdd MUX2X1
XMUX2X1_163 MUX2X1_163/A MUX2X1_163/B BUFX4_22/Y gnd MUX2X1_165/B vdd MUX2X1
XFILL_9_7_0 gnd vdd FILL
XMUX2X1_196 MUX2X1_196/A MUX2X1_196/B BUFX4_5/Y gnd MUX2X1_196/Y vdd MUX2X1
XMUX2X1_185 MUX2X1_185/A MUX2X1_185/B BUFX4_19/Y gnd MUX2X1_185/Y vdd MUX2X1
XNAND2X1_680 BUFX4_249/Y NAND2X1_680/B gnd NAND2X1_680/Y vdd NAND2X1
XNAND2X1_691 BUFX4_267/Y NOR2X1_307/A gnd NAND2X1_691/Y vdd NAND2X1
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XFILL_17_6_0 gnd vdd FILL
XNOR2X1_3 NOR2X1_3/A NOR2X1_2/Y gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_35 BUFX4_114/Y NOR2X1_43/B NOR2X1_45/Y gnd AOI21X1_35/Y vdd AOI21X1
XAOI21X1_13 BUFX4_395/Y NOR2X1_14/B NOR2X1_17/Y gnd AOI21X1_13/Y vdd AOI21X1
XAOI21X1_24 BUFX4_376/Y NOR2X1_27/B NOR2X1_30/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_57 BUFX4_127/Y NOR2X1_77/B NOR2X1_73/Y gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_68 BUFX4_298/Y NOR2X1_90/B NOR2X1_86/Y gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_46 AOI21X1_6/A NOR2X1_55/B NOR2X1_58/Y gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_79 BUFX4_280/Y NOR2X1_96/B NOR2X1_99/Y gnd AOI21X1_79/Y vdd AOI21X1
XOAI21X1_8 BUFX4_300/Y NAND2X1_1/Y OAI21X1_7/Y gnd OAI21X1_8/Y vdd OAI21X1
XFILL_41_4_0 gnd vdd FILL
XINVX1_502 INVX1_502/A gnd INVX1_502/Y vdd INVX1
XOAI21X1_493 BUFX4_169/Y BUFX4_341/Y INVX1_424/A gnd OAI21X1_494/C vdd OAI21X1
XOAI21X1_471 BUFX4_368/Y BUFX4_340/Y NAND2X1_454/B gnd OAI21X1_471/Y vdd OAI21X1
XOAI21X1_460 BUFX4_101/Y NAND2X1_94/Y OAI21X1_460/C gnd OAI21X1_460/Y vdd OAI21X1
XOAI21X1_482 NAND2X1_96/Y BUFX4_124/Y OAI21X1_482/C gnd OAI21X1_482/Y vdd OAI21X1
XFILL_32_4_0 gnd vdd FILL
XOAI21X1_1701 BUFX4_101/Y NAND2X1_872/Y OAI21X1_1701/C gnd DFFPOSX1_350/D vdd OAI21X1
XFILL_23_4_0 gnd vdd FILL
XFILL_6_5_0 gnd vdd FILL
XBUFX4_107 BUFX4_105/A gnd BUFX4_107/Y vdd BUFX4
XBUFX4_118 BUFX4_121/A gnd BUFX4_118/Y vdd BUFX4
XBUFX4_129 INVX8_2/Y gnd BUFX4_129/Y vdd BUFX4
XFILL_14_4_0 gnd vdd FILL
XOAI21X1_1019 INVX1_231/Y BUFX4_226/Y NAND2X1_454/Y gnd MUX2X1_170/B vdd OAI21X1
XOAI21X1_1008 INVX1_220/Y BUFX4_204/Y NAND2X1_442/Y gnd MUX2X1_161/A vdd OAI21X1
XOAI21X1_290 BUFX4_126/Y NAND2X1_67/Y OAI21X1_290/C gnd OAI21X1_290/Y vdd OAI21X1
XDFFPOSX1_609 INVX1_51/A CLKBUF1_22/Y OAI21X1_346/Y gnd vdd DFFPOSX1
XINVX1_310 INVX1_310/A gnd INVX1_310/Y vdd INVX1
XINVX1_321 INVX1_321/A gnd INVX1_321/Y vdd INVX1
XINVX1_332 INVX1_332/A gnd INVX1_332/Y vdd INVX1
XINVX1_343 INVX1_343/A gnd INVX1_343/Y vdd INVX1
XINVX1_354 INVX1_354/A gnd INVX1_354/Y vdd INVX1
XINVX1_376 INVX1_376/A gnd INVX1_376/Y vdd INVX1
XINVX1_387 INVX1_387/A gnd INVX1_387/Y vdd INVX1
XINVX1_365 INVX1_365/A gnd INVX1_365/Y vdd INVX1
XINVX1_398 INVX1_398/A gnd INVX1_398/Y vdd INVX1
XFILL_36_1 gnd vdd FILL
XAOI21X1_303 BUFX4_419/Y NOR2X1_387/B NOR2X1_381/Y gnd AOI21X1_303/Y vdd AOI21X1
XOAI21X1_1531 BUFX4_405/Y BUFX4_91/Y INVX1_330/A gnd OAI21X1_1532/C vdd OAI21X1
XOAI21X1_1520 BUFX4_375/Y NAND2X1_835/Y OAI21X1_1519/Y gnd DFFPOSX1_208/D vdd OAI21X1
XDFFPOSX1_13 NOR2X1_260/A CLKBUF1_18/Y DFFPOSX1_13/D gnd vdd DFFPOSX1
XDFFPOSX1_35 INVX1_127/A CLKBUF1_71/Y DFFPOSX1_35/D gnd vdd DFFPOSX1
XDFFPOSX1_24 NOR2X1_283/A CLKBUF1_40/Y AOI21X1_230/Y gnd vdd DFFPOSX1
XDFFPOSX1_57 NOR2X1_286/A CLKBUF1_37/Y AOI21X1_231/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 INVX1_193/A CLKBUF1_17/Y DFFPOSX1_68/D gnd vdd DFFPOSX1
XOAI21X1_1542 NAND2X1_837/Y BUFX4_113/Y OAI21X1_1542/C gnd DFFPOSX1_227/D vdd OAI21X1
XOAI21X1_1575 BUFX4_113/Y NAND2X1_840/Y OAI21X1_1575/C gnd OAI21X1_1575/Y vdd OAI21X1
XDFFPOSX1_46 NOR2X1_271/A CLKBUF1_9/Y AOI21X1_220/Y gnd vdd DFFPOSX1
XOAI21X1_1564 BUFX4_171/Y BUFX4_95/Y INVX1_332/A gnd OAI21X1_1565/C vdd OAI21X1
XOAI21X1_1553 INVX1_14/Y NOR2X1_352/B NAND2X1_838/Y gnd OAI21X1_1553/Y vdd OAI21X1
XOAI21X1_1597 BUFX4_97/Y NAND2X1_842/Y OAI21X1_1596/Y gnd OAI21X1_1597/Y vdd OAI21X1
XOAI21X1_1586 BUFX4_454/Y INVX2_10/A INVX1_20/A gnd OAI21X1_1587/C vdd OAI21X1
XDFFPOSX1_79 NAND2X1_621/B CLKBUF1_17/Y DFFPOSX1_79/D gnd vdd DFFPOSX1
XFILL_47_8_1 gnd vdd FILL
XFILL_46_3_0 gnd vdd FILL
XFILL_30_7_1 gnd vdd FILL
XDFFPOSX1_417 INVX1_26/A CLKBUF1_30/Y OAI21X1_106/Y gnd vdd DFFPOSX1
XDFFPOSX1_406 INVX1_342/A CLKBUF1_29/Y OAI21X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_428 OAI21X1_127/C CLKBUF1_82/Y OAI21X1_128/Y gnd vdd DFFPOSX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XDFFPOSX1_439 INVX1_408/A CLKBUF1_49/Y OAI21X1_150/Y gnd vdd DFFPOSX1
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XNAND2X1_509 BUFX4_228/Y NOR2X1_17/A gnd NAND2X1_509/Y vdd NAND2X1
XINVX1_173 INVX1_173/A gnd INVX1_173/Y vdd INVX1
XINVX1_195 INVX1_195/A gnd INVX1_195/Y vdd INVX1
XFILL_37_3_0 gnd vdd FILL
XFILL_38_8_1 gnd vdd FILL
XBUFX4_460 INVX8_10/Y gnd BUFX4_460/Y vdd BUFX4
XAOI21X1_100 BUFX4_425/Y NOR2X1_126/B NOR2X1_126/Y gnd AOI21X1_100/Y vdd AOI21X1
XAOI21X1_133 BUFX4_372/Y NOR2X1_158/B NOR2X1_165/Y gnd AOI21X1_133/Y vdd AOI21X1
XFILL_20_2_0 gnd vdd FILL
XFILL_21_7_1 gnd vdd FILL
XAOI21X1_111 BUFX4_304/Y NOR2X1_139/B NOR2X1_139/Y gnd AOI21X1_111/Y vdd AOI21X1
XAOI21X1_122 BUFX4_104/Y NOR2X1_153/B NOR2X1_152/Y gnd AOI21X1_122/Y vdd AOI21X1
XAOI21X1_155 BUFX4_115/Y NOR2X1_197/B NOR2X1_193/Y gnd AOI21X1_155/Y vdd AOI21X1
XAOI21X1_144 BUFX4_131/Y NOR2X1_186/B NOR2X1_180/Y gnd AOI21X1_144/Y vdd AOI21X1
XAOI21X1_166 BUFX4_395/Y NOR2X1_206/B NOR2X1_206/Y gnd AOI21X1_166/Y vdd AOI21X1
XAOI21X1_188 BUFX4_419/Y NOR2X1_236/B NOR2X1_232/Y gnd AOI21X1_188/Y vdd AOI21X1
XAOI21X1_177 BUFX4_378/Y NOR2X1_216/B NOR2X1_218/Y gnd AOI21X1_177/Y vdd AOI21X1
XAOI21X1_199 INVX8_1/Y INVX1_29/Y OR2X2_1/A gnd OAI21X1_814/C vdd AOI21X1
XOAI21X1_1350 BUFX4_112/Y NAND2X1_793/Y OAI21X1_1349/Y gnd DFFPOSX1_75/D vdd OAI21X1
XOAI21X1_1383 BUFX4_168/Y BUFX4_468/Y INVX1_196/A gnd OAI21X1_1383/Y vdd OAI21X1
XOAI21X1_1361 INVX1_38/Y NOR2X1_297/Y NAND2X1_794/Y gnd DFFPOSX1_81/D vdd OAI21X1
XDFFPOSX1_940 NOR2X1_194/A CLKBUF1_18/Y AOI21X1_156/Y gnd vdd DFFPOSX1
XDFFPOSX1_951 INVX1_440/A CLKBUF1_71/Y OAI21X1_726/Y gnd vdd DFFPOSX1
XOAI21X1_1372 INVX1_195/Y NOR2X1_309/Y NAND2X1_805/Y gnd DFFPOSX1_100/D vdd OAI21X1
XDFFPOSX1_984 INVX1_506/A CLKBUF1_73/Y OAI21X1_775/Y gnd vdd DFFPOSX1
XDFFPOSX1_973 NAND2X1_542/B CLKBUF1_59/Y OAI21X1_753/Y gnd vdd DFFPOSX1
XDFFPOSX1_962 INVX1_121/A CLKBUF1_59/Y OAI21X1_731/Y gnd vdd DFFPOSX1
XOAI21X1_1394 BUFX4_125/Y NAND2X1_812/Y OAI21X1_1393/Y gnd OAI21X1_1394/Y vdd OAI21X1
XDFFPOSX1_995 INVX1_187/A CLKBUF1_97/Y OAI21X1_781/Y gnd vdd DFFPOSX1
XFILL_4_8_1 gnd vdd FILL
XFILL_28_3_0 gnd vdd FILL
XFILL_29_8_1 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_12_7_1 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XDFFPOSX1_203 NAND2X1_353/B CLKBUF1_51/Y OAI21X1_1510/Y gnd vdd DFFPOSX1
XDFFPOSX1_236 NOR2X1_353/A CLKBUF1_52/Y AOI21X1_281/Y gnd vdd DFFPOSX1
XDFFPOSX1_214 INVX1_330/A CLKBUF1_52/Y DFFPOSX1_214/D gnd vdd DFFPOSX1
XDFFPOSX1_225 INVX1_15/A CLKBUF1_35/Y DFFPOSX1_225/D gnd vdd DFFPOSX1
XBUFX4_9 clk gnd BUFX4_9/Y vdd BUFX4
XDFFPOSX1_247 INVX1_396/A CLKBUF1_66/Y DFFPOSX1_247/D gnd vdd DFFPOSX1
XDFFPOSX1_269 NAND2X1_496/B CLKBUF1_89/Y DFFPOSX1_269/D gnd vdd DFFPOSX1
XDFFPOSX1_258 INVX1_77/A CLKBUF1_25/Y OAI21X1_1589/Y gnd vdd DFFPOSX1
XNAND2X1_306 BUFX4_246/Y NAND2X1_306/B gnd OAI21X1_881/C vdd NAND2X1
XNAND2X1_317 BUFX4_268/Y OAI21X1_499/C gnd NAND2X1_317/Y vdd NAND2X1
XNAND2X1_339 AOI22X1_17/Y AOI22X1_18/Y gnd AOI22X1_19/D vdd NAND2X1
XNAND2X1_328 BUFX4_189/Y NOR2X1_148/A gnd OAI21X1_902/C vdd NAND2X1
XBUFX4_290 BUFX4_288/A gnd BUFX4_290/Y vdd BUFX4
XNOR2X1_350 BUFX4_92/Y NOR2X1_22/B gnd NOR2X1_352/B vdd NOR2X1
XNOR2X1_361 NOR2X1_361/A NOR2X1_367/B gnd NOR2X1_361/Y vdd NOR2X1
XNOR2X1_383 NOR2X1_383/A NOR2X1_387/B gnd NOR2X1_383/Y vdd NOR2X1
XNOR2X1_372 NOR2X1_372/A NOR2X1_373/B gnd NOR2X1_372/Y vdd NOR2X1
XOAI21X1_823 INVX1_37/Y BUFX4_234/Y OAI21X1_823/C gnd NAND2X1_240/B vdd OAI21X1
XOAI21X1_801 NOR2X1_247/Y NOR2X1_248/Y INVX2_6/Y gnd AOI21X1_195/A vdd OAI21X1
XOAI21X1_812 INVX1_27/Y BUFX4_216/Y OAI21X1_812/C gnd AOI22X1_4/A vdd OAI21X1
XOAI21X1_834 INVX1_46/Y BUFX4_252/Y OAI21X1_834/C gnd MUX2X1_31/A vdd OAI21X1
XOAI21X1_867 INVX1_79/Y BUFX4_219/Y OAI21X1_867/C gnd MUX2X1_56/B vdd OAI21X1
XOAI21X1_845 INVX1_57/Y BUFX4_274/Y OAI21X1_845/C gnd MUX2X1_40/B vdd OAI21X1
XOAI21X1_856 INVX1_68/Y BUFX4_197/Y OAI21X1_856/C gnd MUX2X1_47/A vdd OAI21X1
XOAI21X1_878 INVX1_90/Y BUFX4_241/Y OAI21X1_878/C gnd MUX2X1_64/A vdd OAI21X1
XOAI21X1_889 INVX1_101/Y BUFX4_263/Y OAI21X1_889/C gnd MUX2X1_73/B vdd OAI21X1
XMUX2X1_312 MUX2X1_311/Y MUX2X1_312/B MUX2X1_48/S gnd MUX2X1_312/Y vdd MUX2X1
XMUX2X1_301 MUX2X1_301/A MUX2X1_301/B BUFX4_61/Y gnd MUX2X1_303/B vdd MUX2X1
XMUX2X1_323 MUX2X1_323/A MUX2X1_323/B BUFX4_62/Y gnd MUX2X1_324/A vdd MUX2X1
XOAI21X1_1180 INVX1_392/Y BUFX4_251/Y NAND2X1_628/Y gnd MUX2X1_290/A vdd OAI21X1
XOAI21X1_1191 INVX1_403/Y BUFX4_273/Y NAND2X1_640/Y gnd MUX2X1_299/B vdd OAI21X1
XMUX2X1_345 MUX2X1_345/A MUX2X1_345/B MUX2X1_48/S gnd AOI22X1_72/A vdd MUX2X1
XMUX2X1_356 MUX2X1_356/A MUX2X1_356/B INVX4_1/A gnd MUX2X1_357/A vdd MUX2X1
XMUX2X1_334 MUX2X1_334/A MUX2X1_334/B INVX4_1/A gnd MUX2X1_336/B vdd MUX2X1
XMUX2X1_378 MUX2X1_377/Y MUX2X1_376/Y MUX2X1_48/S gnd MUX2X1_378/Y vdd MUX2X1
XDFFPOSX1_770 INVX1_109/A CLKBUF1_74/Y OAI21X1_572/Y gnd vdd DFFPOSX1
XMUX2X1_367 MUX2X1_367/A MUX2X1_367/B BUFX4_44/Y gnd MUX2X1_369/B vdd MUX2X1
XDFFPOSX1_781 OAI21X1_593/C CLKBUF1_62/Y OAI21X1_594/Y gnd vdd DFFPOSX1
XDFFPOSX1_792 INVX1_494/A CLKBUF1_92/Y OAI21X1_607/Y gnd vdd DFFPOSX1
XNAND2X1_840 INVX8_16/A INVX2_9/Y gnd NAND2X1_840/Y vdd NAND2X1
XNAND2X1_862 BUFX4_157/Y NAND2X1_5/B gnd BUFX4_316/A vdd NAND2X1
XNAND2X1_851 BUFX4_427/Y NOR2X1_358/Y gnd NAND2X1_851/Y vdd NAND2X1
XFILL_44_6_1 gnd vdd FILL
XFILL_43_1_0 gnd vdd FILL
XFILL_34_1_0 gnd vdd FILL
XFILL_35_6_1 gnd vdd FILL
XNOR2X1_90 NOR2X1_90/A NOR2X1_90/B gnd NOR2X1_90/Y vdd NOR2X1
XOAI21X1_119 NOR2X1_51/B BUFX4_175/Y INVX1_471/A gnd OAI21X1_120/C vdd OAI21X1
XOAI21X1_108 BUFX4_422/Y NAND2X1_16/Y OAI21X1_108/C gnd OAI21X1_108/Y vdd OAI21X1
XBUFX2_6 BUFX2_6/A gnd q[5] vdd BUFX2
XNAND2X1_103 BUFX4_334/Y NOR2X1_81/Y gnd OAI21X1_547/C vdd NAND2X1
XNAND2X1_114 BUFX4_330/Y NOR2X1_91/Y gnd OAI21X1_558/C vdd NAND2X1
XNAND2X1_125 INVX1_6/A AOI22X1_69/C gnd BUFX4_105/A vdd NAND2X1
XNAND2X1_147 BUFX4_139/Y NOR2X1_133/Y gnd OAI21X1_620/C vdd NAND2X1
XNAND2X1_136 INVX8_4/A NOR2X1_122/Y gnd OAI21X1_609/C vdd NAND2X1
XNAND2X1_158 BUFX4_431/Y NOR2X1_145/B gnd OAI21X1_660/C vdd NAND2X1
XNAND2X1_169 BUFX4_445/Y NOR2X1_166/Y gnd NAND2X1_169/Y vdd NAND2X1
XNAND2X1_1 INVX2_11/Y INVX8_14/A gnd NAND2X1_1/Y vdd NAND2X1
XFILL_0_1_0 gnd vdd FILL
XFILL_1_6_1 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XFILL_26_6_1 gnd vdd FILL
XNOR2X1_180 MUX2X1_16/A NOR2X1_186/B gnd NOR2X1_180/Y vdd NOR2X1
XNOR2X1_191 MUX2X1_18/A NOR2X1_197/B gnd NOR2X1_191/Y vdd NOR2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XOAI21X1_631 BUFX4_396/Y OAI21X1_635/B OAI21X1_631/C gnd OAI21X1_631/Y vdd OAI21X1
XOAI21X1_620 INVX1_432/Y NOR2X1_133/Y OAI21X1_620/C gnd OAI21X1_620/Y vdd OAI21X1
XOAI21X1_642 BUFX4_153/Y INVX1_4/A OAI21X1_642/C gnd OAI21X1_642/Y vdd OAI21X1
XOAI21X1_653 BUFX4_372/Y OAI21X1_651/B OAI21X1_653/C gnd OAI21X1_653/Y vdd OAI21X1
XOAI21X1_664 INVX1_307/Y NOR2X1_155/Y NAND2X1_162/Y gnd OAI21X1_664/Y vdd OAI21X1
XOAI21X1_675 BUFX4_462/Y BUFX4_66/Y MUX2X1_15/B gnd OAI21X1_675/Y vdd OAI21X1
XAOI21X1_6 AOI21X1_6/A NOR2X1_2/Y NOR2X1_8/Y gnd AOI21X1_6/Y vdd AOI21X1
XOAI21X1_686 BUFX4_98/Y NAND2X1_174/Y OAI21X1_685/Y gnd OAI21X1_686/Y vdd OAI21X1
XOAI21X1_697 BUFX4_146/Y BUFX4_67/Y NAND2X1_469/B gnd OAI21X1_697/Y vdd OAI21X1
XMUX2X1_120 MUX2X1_119/Y MUX2X1_120/B BUFX4_362/Y gnd MUX2X1_120/Y vdd MUX2X1
XMUX2X1_131 MUX2X1_131/A MUX2X1_131/B INVX4_1/A gnd MUX2X1_132/A vdd MUX2X1
XMUX2X1_142 MUX2X1_142/A MUX2X1_142/B BUFX4_46/Y gnd MUX2X1_144/B vdd MUX2X1
XMUX2X1_153 MUX2X1_153/A MUX2X1_153/B BUFX4_362/Y gnd AOI22X1_32/A vdd MUX2X1
XMUX2X1_164 MUX2X1_164/A MUX2X1_164/B BUFX4_47/Y gnd MUX2X1_164/Y vdd MUX2X1
XFILL_9_7_1 gnd vdd FILL
XMUX2X1_197 MUX2X1_197/A MUX2X1_197/B BUFX4_36/Y gnd MUX2X1_197/Y vdd MUX2X1
XFILL_8_2_0 gnd vdd FILL
XMUX2X1_186 MUX2X1_185/Y MUX2X1_186/B BUFX4_362/Y gnd AOI22X1_38/D vdd MUX2X1
XMUX2X1_175 MUX2X1_175/A MUX2X1_175/B BUFX4_39/Y gnd MUX2X1_177/B vdd MUX2X1
XNAND2X1_681 BUFX4_251/Y NOR2X1_217/A gnd NAND2X1_681/Y vdd NAND2X1
XNAND2X1_670 BUFX4_229/Y NOR2X1_131/A gnd NAND2X1_670/Y vdd NAND2X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XNAND2X1_692 BUFX4_269/Y NOR2X1_319/A gnd NAND2X1_692/Y vdd NAND2X1
XFILL_16_1_0 gnd vdd FILL
XFILL_17_6_1 gnd vdd FILL
XDFFPOSX1_1 INVX1_34/A CLKBUF1_71/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XNOR2X1_4 NOR2X1_4/A NOR2X1_2/Y gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_14 BUFX4_96/Y NOR2X1_14/B NOR2X1_18/Y gnd AOI21X1_14/Y vdd AOI21X1
XAOI21X1_25 AOI21X1_1/A NOR2X1_38/B NOR2X1_33/Y gnd AOI21X1_25/Y vdd AOI21X1
XAOI21X1_36 BUFX4_299/Y NOR2X1_43/B NOR2X1_46/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_58 BUFX4_425/Y NOR2X1_77/B NOR2X1_74/Y gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_47 BUFX4_280/Y NOR2X1_55/B NOR2X1_59/Y gnd AOI21X1_47/Y vdd AOI21X1
XAOI21X1_69 BUFX4_399/Y NOR2X1_90/B NOR2X1_87/Y gnd AOI21X1_69/Y vdd AOI21X1
XOAI21X1_9 BUFX4_307/Y BUFX4_319/Y INVX1_275/A gnd OAI21X1_9/Y vdd OAI21X1
XFILL_41_4_1 gnd vdd FILL
XOAI21X1_450 BUFX4_124/Y NAND2X1_94/Y OAI21X1_450/C gnd OAI21X1_450/Y vdd OAI21X1
XOAI21X1_483 BUFX4_172/Y BUFX4_337/Y INVX1_104/A gnd OAI21X1_483/Y vdd OAI21X1
XOAI21X1_472 BUFX4_300/Y NAND2X1_95/Y OAI21X1_471/Y gnd OAI21X1_472/Y vdd OAI21X1
XOAI21X1_461 BUFX4_310/Y BUFX4_336/Y INVX1_423/A gnd OAI21X1_462/C vdd OAI21X1
XINVX1_503 INVX1_503/A gnd INVX1_503/Y vdd INVX1
XOAI21X1_494 NAND2X1_96/Y BUFX4_284/Y OAI21X1_494/C gnd OAI21X1_494/Y vdd OAI21X1
XFILL_48_0_0 gnd vdd FILL
XFILL_32_4_1 gnd vdd FILL
XOAI21X1_1702 BUFX4_87/Y OAI21X1_1/B NAND2X1_639/B gnd OAI21X1_1703/C vdd OAI21X1
XFILL_39_0_0 gnd vdd FILL
XFILL_23_4_1 gnd vdd FILL
XBUFX4_119 BUFX4_121/A gnd INVX1_4/A vdd BUFX4
XFILL_6_5_1 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XBUFX4_108 BUFX4_105/A gnd BUFX4_108/Y vdd BUFX4
XFILL_14_4_1 gnd vdd FILL
XOAI21X1_1009 INVX1_221/Y BUFX4_206/Y NAND2X1_444/Y gnd MUX2X1_163/B vdd OAI21X1
XOAI21X1_291 BUFX4_411/Y BUFX4_433/Y NAND2X1_309/B gnd OAI21X1_291/Y vdd OAI21X1
XINVX1_300 INVX1_300/A gnd INVX1_300/Y vdd INVX1
XOAI21X1_280 NAND2X1_66/Y BUFX4_299/Y OAI21X1_279/Y gnd OAI21X1_280/Y vdd OAI21X1
XINVX1_311 INVX1_311/A gnd INVX1_311/Y vdd INVX1
XINVX1_333 INVX1_333/A gnd INVX1_333/Y vdd INVX1
XINVX1_344 INVX1_344/A gnd INVX1_344/Y vdd INVX1
XINVX1_322 INVX1_322/A gnd INVX1_322/Y vdd INVX1
XINVX1_355 INVX1_355/A gnd INVX1_355/Y vdd INVX1
XINVX1_377 INVX1_377/A gnd INVX1_377/Y vdd INVX1
XINVX1_366 INVX1_366/A gnd INVX1_366/Y vdd INVX1
XINVX1_399 INVX1_399/A gnd INVX1_399/Y vdd INVX1
XINVX1_388 INVX1_388/A gnd INVX1_388/Y vdd INVX1
XFILL_36_2 gnd vdd FILL
XFILL_29_1 gnd vdd FILL
XAOI21X1_304 BUFX4_117/Y NOR2X1_387/B NOR2X1_382/Y gnd AOI21X1_304/Y vdd AOI21X1
XDFFPOSX1_14 NOR2X1_261/A CLKBUF1_90/Y DFFPOSX1_14/D gnd vdd DFFPOSX1
XOAI21X1_1521 BUFX4_405/Y BUFX4_91/Y MUX2X1_30/B gnd OAI21X1_1521/Y vdd OAI21X1
XOAI21X1_1532 NAND2X1_836/Y BUFX4_96/Y OAI21X1_1532/C gnd DFFPOSX1_214/D vdd OAI21X1
XOAI21X1_1510 BUFX4_115/Y NAND2X1_835/Y OAI21X1_1510/C gnd OAI21X1_1510/Y vdd OAI21X1
XDFFPOSX1_36 INVX1_191/A CLKBUF1_44/Y DFFPOSX1_36/D gnd vdd DFFPOSX1
XDFFPOSX1_25 INVX1_33/A CLKBUF1_71/Y DFFPOSX1_25/D gnd vdd DFFPOSX1
XDFFPOSX1_69 INVX1_257/A CLKBUF1_43/Y DFFPOSX1_69/D gnd vdd DFFPOSX1
XDFFPOSX1_47 NOR2X1_272/A CLKBUF1_86/Y AOI21X1_221/Y gnd vdd DFFPOSX1
XOAI21X1_1554 BUFX4_166/Y INVX2_9/A NAND2X1_211/A gnd OAI21X1_1554/Y vdd OAI21X1
XOAI21X1_1543 BUFX4_312/Y BUFX4_93/Y INVX1_203/A gnd OAI21X1_1544/C vdd OAI21X1
XOAI21X1_1565 NAND2X1_839/Y BUFX4_96/Y OAI21X1_1565/C gnd DFFPOSX1_246/D vdd OAI21X1
XDFFPOSX1_58 NOR2X1_287/A CLKBUF1_50/Y DFFPOSX1_58/D gnd vdd DFFPOSX1
XOAI21X1_1576 BUFX4_410/Y BUFX4_95/Y NAND2X1_425/B gnd OAI21X1_1576/Y vdd OAI21X1
XOAI21X1_1598 BUFX4_454/Y BUFX4_348/Y INVX1_397/A gnd OAI21X1_1598/Y vdd OAI21X1
XOAI21X1_1587 BUFX4_129/Y NAND2X1_842/Y OAI21X1_1587/C gnd DFFPOSX1_257/D vdd OAI21X1
XFILL_46_3_1 gnd vdd FILL
XDFFPOSX1_407 INVX1_406/A CLKBUF1_75/Y OAI21X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_418 INVX1_87/A CLKBUF1_41/Y OAI21X1_108/Y gnd vdd DFFPOSX1
XDFFPOSX1_429 NAND2X1_506/B CLKBUF1_48/Y OAI21X1_130/Y gnd vdd DFFPOSX1
XINVX1_130 INVX1_130/A gnd INVX1_130/Y vdd INVX1
XINVX1_141 INVX1_141/A gnd INVX1_141/Y vdd INVX1
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XINVX1_185 INVX1_185/A gnd INVX1_185/Y vdd INVX1
XINVX1_174 INVX1_174/A gnd INVX1_174/Y vdd INVX1
XINVX1_196 INVX1_196/A gnd INVX1_196/Y vdd INVX1
XCLKBUF1_100 BUFX4_9/Y gnd CLKBUF1_100/Y vdd CLKBUF1
XFILL_37_3_1 gnd vdd FILL
XBUFX4_450 d[1] gnd BUFX4_450/Y vdd BUFX4
XBUFX4_461 INVX8_10/Y gnd BUFX4_461/Y vdd BUFX4
XAOI21X1_123 BUFX4_287/Y NOR2X1_153/B NOR2X1_153/Y gnd AOI21X1_123/Y vdd AOI21X1
XAOI21X1_112 BUFX4_402/Y NOR2X1_139/B NOR2X1_140/Y gnd AOI21X1_112/Y vdd AOI21X1
XAOI21X1_101 BUFX4_110/Y NOR2X1_126/B NOR2X1_127/Y gnd AOI21X1_101/Y vdd AOI21X1
XAOI21X1_167 BUFX4_98/Y NOR2X1_206/B NOR2X1_207/Y gnd AOI21X1_167/Y vdd AOI21X1
XAOI21X1_145 BUFX4_426/Y NOR2X1_186/B NOR2X1_181/Y gnd AOI21X1_145/Y vdd AOI21X1
XAOI21X1_156 BUFX4_301/Y NOR2X1_197/B NOR2X1_194/Y gnd AOI21X1_156/Y vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_134 BUFX4_129/Y NOR2X1_166/Y NOR2X1_167/Y gnd AOI21X1_134/Y vdd AOI21X1
XAOI21X1_178 BUFX4_123/Y NOR2X1_222/B NOR2X1_220/Y gnd AOI21X1_178/Y vdd AOI21X1
XAOI21X1_189 BUFX4_113/Y NOR2X1_236/B NOR2X1_233/Y gnd AOI21X1_189/Y vdd AOI21X1
XOAI21X1_1340 BUFX4_99/Y NAND2X1_792/Y OAI21X1_1339/Y gnd DFFPOSX1_70/D vdd OAI21X1
XOAI21X1_1351 BUFX4_154/Y BUFX4_467/Y DFFPOSX1_76/Q gnd OAI21X1_1351/Y vdd OAI21X1
XDFFPOSX1_930 INVX1_119/A CLKBUF1_14/Y OAI21X1_714/Y gnd vdd DFFPOSX1
XDFFPOSX1_941 NOR2X1_195/A CLKBUF1_9/Y AOI21X1_157/Y gnd vdd DFFPOSX1
XOAI21X1_1373 INVX1_259/Y NOR2X1_309/Y NAND2X1_806/Y gnd OAI21X1_1373/Y vdd OAI21X1
XOAI21X1_1362 INVX1_66/Y NOR2X1_297/Y NAND2X1_795/Y gnd DFFPOSX1_82/D vdd OAI21X1
XOAI21X1_1384 NAND2X1_811/Y BUFX4_305/Y OAI21X1_1383/Y gnd OAI21X1_1384/Y vdd OAI21X1
XDFFPOSX1_952 INVX1_504/A CLKBUF1_50/Y OAI21X1_727/Y gnd vdd DFFPOSX1
XDFFPOSX1_974 NAND2X1_611/B CLKBUF1_69/Y OAI21X1_755/Y gnd vdd DFFPOSX1
XDFFPOSX1_963 INVX1_185/A CLKBUF1_59/Y OAI21X1_733/Y gnd vdd DFFPOSX1
XDFFPOSX1_985 MUX2X1_23/A CLKBUF1_65/Y AOI21X1_170/Y gnd vdd DFFPOSX1
XOAI21X1_1395 BUFX4_417/Y INVX2_7/A NAND2X1_279/B gnd OAI21X1_1396/C vdd OAI21X1
XDFFPOSX1_996 INVX1_251/A CLKBUF1_73/Y OAI21X1_783/Y gnd vdd DFFPOSX1
XFILL_28_3_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XDFFPOSX1_204 NAND2X1_422/B CLKBUF1_5/Y DFFPOSX1_204/D gnd vdd DFFPOSX1
XDFFPOSX1_237 NOR2X1_354/A CLKBUF1_66/Y AOI21X1_282/Y gnd vdd DFFPOSX1
XDFFPOSX1_226 INVX1_75/A CLKBUF1_66/Y DFFPOSX1_226/D gnd vdd DFFPOSX1
XDFFPOSX1_215 INVX1_394/A CLKBUF1_35/Y DFFPOSX1_215/D gnd vdd DFFPOSX1
XDFFPOSX1_248 INVX1_460/A CLKBUF1_64/Y DFFPOSX1_248/D gnd vdd DFFPOSX1
XDFFPOSX1_259 INVX1_141/A CLKBUF1_25/Y OAI21X1_1591/Y gnd vdd DFFPOSX1
XNAND2X1_307 BUFX4_248/Y NOR2X1_44/A gnd OAI21X1_882/C vdd NAND2X1
XNAND2X1_318 BUFX4_270/Y NAND2X1_318/B gnd OAI21X1_893/C vdd NAND2X1
XNAND2X1_329 BUFX4_191/Y NOR2X1_159/A gnd OAI21X1_903/C vdd NAND2X1
XBUFX4_291 BUFX4_288/A gnd AOI22X1_6/C vdd BUFX4
XBUFX4_280 INVX8_8/Y gnd BUFX4_280/Y vdd BUFX4
XNOR2X1_351 NOR2X1_351/A NOR2X1_352/B gnd NOR2X1_351/Y vdd NOR2X1
XNOR2X1_340 NOR2X1_340/A NOR2X1_338/B gnd NOR2X1_340/Y vdd NOR2X1
XNOR2X1_384 NOR2X1_384/A NOR2X1_387/B gnd NOR2X1_384/Y vdd NOR2X1
XNOR2X1_362 NOR2X1_362/A NOR2X1_367/B gnd NOR2X1_362/Y vdd NOR2X1
XNOR2X1_373 NOR2X1_373/A NOR2X1_373/B gnd NOR2X1_373/Y vdd NOR2X1
XOAI21X1_824 INVX1_38/Y BUFX4_236/Y OAI21X1_824/C gnd NAND2X1_242/B vdd OAI21X1
XOAI21X1_813 INVX1_28/Y BUFX4_218/Y OAI21X1_813/C gnd AOI22X1_4/D vdd OAI21X1
XOAI21X1_802 INVX8_1/Y OAI21X1_802/B AOI21X1_196/Y gnd NAND3X1_1/A vdd OAI21X1
XOAI21X1_857 INVX1_69/Y BUFX4_199/Y NAND2X1_280/Y gnd MUX2X1_49/B vdd OAI21X1
XOAI21X1_846 INVX1_58/Y BUFX4_276/Y OAI21X1_846/C gnd MUX2X1_40/A vdd OAI21X1
XOAI21X1_835 INVX1_47/Y BUFX4_254/Y OAI21X1_835/C gnd MUX2X1_32/B vdd OAI21X1
XOAI21X1_879 INVX1_91/Y BUFX4_243/Y OAI21X1_879/C gnd MUX2X1_65/B vdd OAI21X1
XOAI21X1_868 INVX1_80/Y BUFX4_221/Y OAI21X1_868/C gnd MUX2X1_56/A vdd OAI21X1
XMUX2X1_313 MUX2X1_313/A MUX2X1_313/B BUFX4_80/Y gnd MUX2X1_315/B vdd MUX2X1
XMUX2X1_302 MUX2X1_302/A MUX2X1_302/B BUFX4_49/Y gnd MUX2X1_303/A vdd MUX2X1
XOAI21X1_1181 INVX1_393/Y BUFX4_253/Y NAND2X1_629/Y gnd MUX2X1_292/B vdd OAI21X1
XOAI21X1_1192 INVX1_404/Y BUFX4_275/Y NAND2X1_641/Y gnd MUX2X1_299/A vdd OAI21X1
XOAI21X1_1170 INVX1_382/Y BUFX4_231/Y NAND2X1_618/Y gnd MUX2X1_283/A vdd OAI21X1
XMUX2X1_346 MUX2X1_346/A MUX2X1_346/B BUFX4_63/Y gnd MUX2X1_348/B vdd MUX2X1
XMUX2X1_335 MUX2X1_335/A MUX2X1_335/B BUFX4_80/Y gnd MUX2X1_336/A vdd MUX2X1
XMUX2X1_357 MUX2X1_357/A MUX2X1_355/Y BUFX4_364/Y gnd AOI22X1_75/A vdd MUX2X1
XMUX2X1_324 MUX2X1_324/A MUX2X1_324/B BUFX4_364/Y gnd AOI22X1_67/D vdd MUX2X1
XMUX2X1_368 MUX2X1_368/A MUX2X1_368/B BUFX4_60/Y gnd MUX2X1_368/Y vdd MUX2X1
XDFFPOSX1_793 MUX2X1_2/A CLKBUF1_74/Y AOI21X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_782 OAI21X1_595/C CLKBUF1_26/Y OAI21X1_596/Y gnd vdd DFFPOSX1
XDFFPOSX1_771 INVX1_173/A CLKBUF1_62/Y OAI21X1_574/Y gnd vdd DFFPOSX1
XDFFPOSX1_760 INVX1_492/A CLKBUF1_7/Y OAI21X1_568/Y gnd vdd DFFPOSX1
XNAND2X1_830 BUFX4_140/Y NOR2X1_331/Y gnd NAND2X1_830/Y vdd NAND2X1
XNAND2X1_863 BUFX4_164/Y NOR2X1_378/Y gnd NAND2X1_863/Y vdd NAND2X1
XNAND2X1_841 BUFX4_354/Y NAND2X1_5/B gnd BUFX4_344/A vdd NAND2X1
XNAND2X1_852 BUFX4_163/Y NOR2X1_368/Y gnd NAND2X1_852/Y vdd NAND2X1
XFILL_43_1_1 gnd vdd FILL
XNOR2X1_80 NOR2X1_80/A NOR2X1_77/B gnd NOR2X1_80/Y vdd NOR2X1
XFILL_34_1_1 gnd vdd FILL
XNOR2X1_91 NOR2X1_91/A NOR2X1_91/B gnd NOR2X1_91/Y vdd NOR2X1
XFILL_11_1 gnd vdd FILL
XOAI21X1_109 NOR2X1_51/B BUFX4_173/Y INVX1_151/A gnd OAI21X1_110/C vdd OAI21X1
XBUFX2_7 BUFX2_7/A gnd q[6] vdd BUFX2
XNAND2X1_104 BUFX4_144/Y NOR2X1_81/Y gnd NAND2X1_104/Y vdd NAND2X1
XNAND2X1_115 BUFX4_140/Y NOR2X1_91/Y gnd OAI21X1_559/C vdd NAND2X1
XNAND2X1_126 INVX8_10/A INVX1_3/Y gnd OAI21X1_584/B vdd NAND2X1
XNAND2X1_148 BUFX4_430/Y NOR2X1_133/Y gnd OAI21X1_621/C vdd NAND2X1
XNAND2X1_137 INVX8_5/A NOR2X1_122/Y gnd NAND2X1_137/Y vdd NAND2X1
XNAND2X1_159 BUFX4_449/Y NOR2X1_155/Y gnd OAI21X1_661/C vdd NAND2X1
XNAND2X1_2 INVX2_11/Y INVX8_15/A gnd NAND2X1_2/Y vdd NAND2X1
XFILL_25_1_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_170 NOR2X1_170/A NOR2X1_173/B gnd NOR2X1_170/Y vdd NOR2X1
XNOR2X1_192 NOR2X1_192/A NOR2X1_197/B gnd NOR2X1_192/Y vdd NOR2X1
XNOR2X1_181 NOR2X1_181/A NOR2X1_186/B gnd NOR2X1_181/Y vdd NOR2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XOAI21X1_632 BUFX4_456/Y BUFX4_120/Y INVX1_369/A gnd OAI21X1_633/C vdd OAI21X1
XOAI21X1_621 INVX1_496/Y NOR2X1_133/Y OAI21X1_621/C gnd OAI21X1_621/Y vdd OAI21X1
XOAI21X1_610 INVX1_239/Y NOR2X1_122/Y NAND2X1_137/Y gnd OAI21X1_610/Y vdd OAI21X1
XAOI21X1_7 BUFX4_279/Y NOR2X1_2/Y NOR2X1_9/Y gnd AOI21X1_7/Y vdd AOI21X1
XOAI21X1_654 INVX1_114/Y NOR2X1_145/B OAI21X1_654/C gnd OAI21X1_654/Y vdd OAI21X1
XOAI21X1_665 INVX1_371/Y NOR2X1_155/Y OAI21X1_665/C gnd OAI21X1_665/Y vdd OAI21X1
XOAI21X1_643 BUFX4_116/Y OAI21X1_651/B OAI21X1_642/Y gnd OAI21X1_643/Y vdd OAI21X1
XOAI21X1_676 BUFX4_131/Y NAND2X1_174/Y OAI21X1_675/Y gnd OAI21X1_676/Y vdd OAI21X1
XOAI21X1_698 BUFX4_301/Y OAI21X1_704/B OAI21X1_697/Y gnd OAI21X1_698/Y vdd OAI21X1
XOAI21X1_687 BUFX4_462/Y INVX1_5/A INVX1_437/A gnd OAI21X1_687/Y vdd OAI21X1
XMUX2X1_121 MUX2X1_121/A MUX2X1_121/B BUFX4_61/Y gnd MUX2X1_123/B vdd MUX2X1
XMUX2X1_132 MUX2X1_132/A MUX2X1_130/Y MUX2X1_7/S gnd AOI22X1_27/D vdd MUX2X1
XMUX2X1_110 MUX2X1_110/A MUX2X1_110/B BUFX4_80/Y gnd MUX2X1_111/A vdd MUX2X1
XMUX2X1_154 MUX2X1_154/A MUX2X1_154/B INVX4_1/A gnd MUX2X1_154/Y vdd MUX2X1
XMUX2X1_165 MUX2X1_164/Y MUX2X1_165/B MUX2X1_7/S gnd AOI22X1_35/A vdd MUX2X1
XMUX2X1_143 MUX2X1_143/A MUX2X1_143/B BUFX4_62/Y gnd MUX2X1_143/Y vdd MUX2X1
XDFFPOSX1_590 NOR2X1_68/A CLKBUF1_16/Y AOI21X1_54/Y gnd vdd DFFPOSX1
XMUX2X1_198 MUX2X1_197/Y MUX2X1_196/Y MUX2X1_7/S gnd MUX2X1_198/Y vdd MUX2X1
XMUX2X1_187 MUX2X1_187/A MUX2X1_187/B BUFX4_44/Y gnd MUX2X1_187/Y vdd MUX2X1
XMUX2X1_176 MUX2X1_176/A MUX2X1_176/B INVX4_1/A gnd MUX2X1_177/A vdd MUX2X1
XFILL_8_2_1 gnd vdd FILL
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XNAND2X1_660 BUFX4_211/Y OAI21X1_445/C gnd NAND2X1_660/Y vdd NAND2X1
XNAND2X1_682 BUFX4_253/Y NOR2X1_226/A gnd NAND2X1_682/Y vdd NAND2X1
XNAND2X1_671 BUFX4_231/Y NOR2X1_142/A gnd NAND2X1_671/Y vdd NAND2X1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XNAND2X1_693 BUFX4_271/Y NAND2X1_693/B gnd NAND2X1_693/Y vdd NAND2X1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XDFFPOSX1_2 INVX1_62/A CLKBUF1_90/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_2/Y gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_15 BUFX4_285/Y NOR2X1_14/B NOR2X1_19/Y gnd AOI21X1_15/Y vdd AOI21X1
XAOI21X1_26 BUFX4_423/Y NOR2X1_38/B NOR2X1_34/Y gnd AOI21X1_26/Y vdd AOI21X1
XAOI21X1_37 BUFX4_394/Y NOR2X1_43/B NOR2X1_47/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_59 BUFX4_110/Y NOR2X1_77/B NOR2X1_75/Y gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_48 BUFX4_379/Y NOR2X1_55/B NOR2X1_60/Y gnd AOI21X1_48/Y vdd AOI21X1
XFILL_10_8_0 gnd vdd FILL
XOAI21X1_440 BUFX4_302/Y NAND2X1_93/Y OAI21X1_440/C gnd OAI21X1_440/Y vdd OAI21X1
XOAI21X1_484 NAND2X1_96/Y BUFX4_421/Y OAI21X1_483/Y gnd OAI21X1_484/Y vdd OAI21X1
XOAI21X1_451 BUFX4_308/Y BUFX4_342/Y INVX1_103/A gnd OAI21X1_452/C vdd OAI21X1
XOAI21X1_473 BUFX4_368/Y BUFX4_340/Y NAND2X1_523/B gnd OAI21X1_474/C vdd OAI21X1
XOAI21X1_462 BUFX4_284/Y NAND2X1_94/Y OAI21X1_462/C gnd OAI21X1_462/Y vdd OAI21X1
XOAI21X1_495 BUFX4_172/Y BUFX4_337/Y INVX1_488/A gnd OAI21X1_495/Y vdd OAI21X1
XINVX1_504 INVX1_504/A gnd INVX1_504/Y vdd INVX1
XFILL_48_0_1 gnd vdd FILL
XNAND2X1_490 BUFX4_192/Y NAND2X1_490/B gnd NAND2X1_490/Y vdd NAND2X1
XOAI21X1_1703 BUFX4_283/Y NAND2X1_872/Y OAI21X1_1703/C gnd OAI21X1_1703/Y vdd OAI21X1
XFILL_39_0_1 gnd vdd FILL
XBUFX4_109 INVX8_4/Y gnd BUFX4_109/Y vdd BUFX4
XFILL_5_0_1 gnd vdd FILL
XFILL_42_7_0 gnd vdd FILL
XOAI21X1_281 BUFX4_165/Y BUFX4_437/Y INVX1_288/A gnd OAI21X1_281/Y vdd OAI21X1
XOAI21X1_292 BUFX4_418/Y NAND2X1_67/Y OAI21X1_291/Y gnd OAI21X1_292/Y vdd OAI21X1
XINVX1_301 INVX1_301/A gnd INVX1_301/Y vdd INVX1
XOAI21X1_270 INVX1_351/Y NOR2X1_51/Y NAND2X1_63/Y gnd OAI21X1_270/Y vdd OAI21X1
XINVX1_312 INVX1_312/A gnd INVX1_312/Y vdd INVX1
XINVX1_323 INVX1_323/A gnd INVX1_323/Y vdd INVX1
XINVX1_334 INVX1_334/A gnd INVX1_334/Y vdd INVX1
XINVX1_356 INVX1_356/A gnd INVX1_356/Y vdd INVX1
XINVX1_345 INVX1_345/A gnd INVX1_345/Y vdd INVX1
XINVX1_378 INVX1_378/A gnd INVX1_378/Y vdd INVX1
XINVX1_367 INVX1_367/A gnd INVX1_367/Y vdd INVX1
XINVX1_389 INVX1_389/A gnd INVX1_389/Y vdd INVX1
XFILL_36_3 gnd vdd FILL
XFILL_29_2 gnd vdd FILL
XFILL_33_7_0 gnd vdd FILL
XAOI21X1_305 BUFX4_302/Y NOR2X1_387/B NOR2X1_383/Y gnd AOI21X1_305/Y vdd AOI21X1
XOAI21X1_1522 NAND2X1_836/Y BUFX4_128/Y OAI21X1_1521/Y gnd DFFPOSX1_209/D vdd OAI21X1
XOAI21X1_1500 BUFX4_98/Y NAND2X1_834/Y OAI21X1_1499/Y gnd DFFPOSX1_198/D vdd OAI21X1
XOAI21X1_1511 BUFX4_147/Y BUFX4_92/Y NAND2X1_422/B gnd OAI21X1_1512/C vdd OAI21X1
XDFFPOSX1_15 NOR2X1_262/A CLKBUF1_14/Y DFFPOSX1_15/D gnd vdd DFFPOSX1
XDFFPOSX1_26 INVX1_61/A CLKBUF1_5/Y DFFPOSX1_26/D gnd vdd DFFPOSX1
XOAI21X1_1566 BUFX4_166/Y BUFX4_92/Y INVX1_396/A gnd OAI21X1_1567/C vdd OAI21X1
XDFFPOSX1_48 NOR2X1_273/A CLKBUF1_90/Y DFFPOSX1_48/D gnd vdd DFFPOSX1
XOAI21X1_1555 NAND2X1_839/Y BUFX4_128/Y OAI21X1_1554/Y gnd DFFPOSX1_241/D vdd OAI21X1
XOAI21X1_1533 BUFX4_405/Y BUFX4_89/Y INVX1_394/A gnd OAI21X1_1534/C vdd OAI21X1
XOAI21X1_1544 NAND2X1_837/Y BUFX4_303/Y OAI21X1_1544/C gnd DFFPOSX1_228/D vdd OAI21X1
XDFFPOSX1_59 NOR2X1_288/A CLKBUF1_2/Y DFFPOSX1_59/D gnd vdd DFFPOSX1
XDFFPOSX1_37 INVX1_255/A CLKBUF1_71/Y DFFPOSX1_37/D gnd vdd DFFPOSX1
XOAI21X1_1577 BUFX4_303/Y NAND2X1_840/Y OAI21X1_1576/Y gnd DFFPOSX1_252/D vdd OAI21X1
XOAI21X1_1599 BUFX4_279/Y NAND2X1_842/Y OAI21X1_1598/Y gnd OAI21X1_1599/Y vdd OAI21X1
XOAI21X1_1588 BUFX4_454/Y BUFX4_344/Y INVX1_77/A gnd OAI21X1_1589/C vdd OAI21X1
XFILL_24_7_0 gnd vdd FILL
XFILL_7_8_0 gnd vdd FILL
XCLKBUF1_90 BUFX4_16/Y gnd CLKBUF1_90/Y vdd CLKBUF1
XFILL_15_7_0 gnd vdd FILL
XDFFPOSX1_408 INVX1_470/A CLKBUF1_72/Y OAI21X1_88/Y gnd vdd DFFPOSX1
XDFFPOSX1_419 INVX1_151/A CLKBUF1_27/Y OAI21X1_110/Y gnd vdd DFFPOSX1
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XINVX1_186 INVX1_186/A gnd INVX1_186/Y vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XINVX1_197 INVX1_197/A gnd INVX1_197/Y vdd INVX1
XCLKBUF1_101 BUFX4_16/Y gnd CLKBUF1_101/Y vdd CLKBUF1
XBUFX4_440 BUFX4_439/A gnd BUFX4_440/Y vdd BUFX4
XBUFX4_462 INVX8_10/Y gnd BUFX4_462/Y vdd BUFX4
XBUFX4_451 d[1] gnd INVX8_3/A vdd BUFX4
XFILL_41_1 gnd vdd FILL
XAOI21X1_124 BUFX4_372/Y NOR2X1_153/B NOR2X1_154/Y gnd AOI21X1_124/Y vdd AOI21X1
XAOI21X1_113 BUFX4_96/Y NOR2X1_139/B NOR2X1_141/Y gnd AOI21X1_113/Y vdd AOI21X1
XAOI21X1_102 BUFX4_304/Y NOR2X1_126/B NOR2X1_128/Y gnd AOI21X1_102/Y vdd AOI21X1
XAOI21X1_146 BUFX4_115/Y NOR2X1_186/B NOR2X1_182/Y gnd AOI21X1_146/Y vdd AOI21X1
XAOI21X1_157 BUFX4_402/Y NOR2X1_197/B NOR2X1_195/Y gnd AOI21X1_157/Y vdd AOI21X1
XAOI21X1_135 BUFX4_129/Y NOR2X1_173/B NOR2X1_169/Y gnd AOI21X1_135/Y vdd AOI21X1
XAOI21X1_168 BUFX4_285/Y NOR2X1_206/B NOR2X1_208/Y gnd AOI21X1_168/Y vdd AOI21X1
XAOI21X1_179 BUFX4_419/Y NOR2X1_222/B NOR2X1_221/Y gnd AOI21X1_179/Y vdd AOI21X1
XOAI21X1_1330 BUFX4_125/Y NAND2X1_792/Y OAI21X1_1329/Y gnd DFFPOSX1_65/D vdd OAI21X1
XOAI21X1_1341 BUFX4_460/Y BUFX4_465/Y INVX1_385/A gnd OAI21X1_1341/Y vdd OAI21X1
XOAI21X1_1363 INVX1_130/Y NOR2X1_297/Y NAND2X1_796/Y gnd DFFPOSX1_83/D vdd OAI21X1
XOAI21X1_1352 BUFX4_305/Y NAND2X1_793/Y OAI21X1_1351/Y gnd DFFPOSX1_76/D vdd OAI21X1
XDFFPOSX1_931 INVX1_183/A CLKBUF1_86/Y OAI21X1_715/Y gnd vdd DFFPOSX1
XDFFPOSX1_920 INVX1_502/A CLKBUF1_21/Y OAI21X1_713/Y gnd vdd DFFPOSX1
XDFFPOSX1_942 NOR2X1_196/A CLKBUF1_21/Y AOI21X1_158/Y gnd vdd DFFPOSX1
XOAI21X1_1374 INVX1_323/Y NOR2X1_309/Y NAND2X1_807/Y gnd DFFPOSX1_102/D vdd OAI21X1
XOAI21X1_1385 BUFX4_168/Y BUFX4_467/Y INVX1_260/A gnd OAI21X1_1385/Y vdd OAI21X1
XDFFPOSX1_953 MUX2X1_19/A CLKBUF1_9/Y AOI21X1_162/Y gnd vdd DFFPOSX1
XDFFPOSX1_964 INVX1_249/A CLKBUF1_67/Y OAI21X1_735/Y gnd vdd DFFPOSX1
XDFFPOSX1_975 NAND2X1_680/B CLKBUF1_59/Y OAI21X1_757/Y gnd vdd DFFPOSX1
XOAI21X1_1396 BUFX4_420/Y NAND2X1_812/Y OAI21X1_1396/C gnd DFFPOSX1_122/D vdd OAI21X1
XDFFPOSX1_997 INVX1_315/A CLKBUF1_73/Y OAI21X1_785/Y gnd vdd DFFPOSX1
XDFFPOSX1_986 NOR2X1_212/A CLKBUF1_33/Y AOI21X1_171/Y gnd vdd DFFPOSX1
XFILL_47_6_0 gnd vdd FILL
XFILL_30_5_0 gnd vdd FILL
XDFFPOSX1_205 NAND2X1_491/B CLKBUF1_76/Y OAI21X1_1514/Y gnd vdd DFFPOSX1
XDFFPOSX1_227 INVX1_139/A CLKBUF1_66/Y DFFPOSX1_227/D gnd vdd DFFPOSX1
XDFFPOSX1_216 INVX1_458/A CLKBUF1_35/Y DFFPOSX1_216/D gnd vdd DFFPOSX1
XDFFPOSX1_238 NOR2X1_355/A CLKBUF1_52/Y AOI21X1_283/Y gnd vdd DFFPOSX1
XDFFPOSX1_249 INVX1_16/A CLKBUF1_35/Y OAI21X1_1571/Y gnd vdd DFFPOSX1
XNAND2X1_308 BUFX4_250/Y NOR2X1_54/A gnd OAI21X1_883/C vdd NAND2X1
XNAND2X1_319 BUFX4_272/Y NOR2X1_84/A gnd NAND2X1_319/Y vdd NAND2X1
XFILL_38_6_0 gnd vdd FILL
XBUFX4_281 INVX8_8/Y gnd BUFX4_281/Y vdd BUFX4
XBUFX4_270 BUFX4_28/Y gnd BUFX4_270/Y vdd BUFX4
XNOR2X1_341 BUFX4_91/Y BUFX4_87/Y gnd NOR2X1_342/B vdd NOR2X1
XNOR2X1_352 NOR2X1_352/A NOR2X1_352/B gnd NOR2X1_352/Y vdd NOR2X1
XBUFX4_292 BUFX4_288/A gnd BUFX4_292/Y vdd BUFX4
XNOR2X1_330 NOR2X1_330/A NOR2X1_325/B gnd NOR2X1_330/Y vdd NOR2X1
XNOR2X1_385 NOR2X1_385/A NOR2X1_387/B gnd NOR2X1_385/Y vdd NOR2X1
XNOR2X1_363 NOR2X1_363/A NOR2X1_367/B gnd NOR2X1_363/Y vdd NOR2X1
XNOR2X1_374 NOR2X1_374/A NOR2X1_373/B gnd NOR2X1_374/Y vdd NOR2X1
XFILL_21_5_0 gnd vdd FILL
XOAI21X1_814 INVX8_1/Y NOR2X1_33/A OAI21X1_814/C gnd NAND3X1_4/A vdd OAI21X1
XOAI21X1_803 INVX1_18/Y BUFX4_202/Y OAI21X1_803/C gnd NAND2X1_215/B vdd OAI21X1
XOAI21X1_858 INVX1_70/Y BUFX4_201/Y OAI21X1_858/C gnd MUX2X1_49/A vdd OAI21X1
XOAI21X1_825 INVX1_39/Y BUFX4_238/Y OAI21X1_825/C gnd NAND2X1_244/B vdd OAI21X1
XOAI21X1_847 INVX1_59/Y BUFX4_278/Y OAI21X1_847/C gnd MUX2X1_41/B vdd OAI21X1
XOAI21X1_836 INVX1_48/Y BUFX4_256/Y NAND2X1_258/Y gnd MUX2X1_32/A vdd OAI21X1
XOAI21X1_869 INVX1_81/Y BUFX4_223/Y OAI21X1_869/C gnd MUX2X1_58/B vdd OAI21X1
XMUX2X1_314 MUX2X1_314/A MUX2X1_314/B BUFX4_81/Y gnd MUX2X1_314/Y vdd MUX2X1
XMUX2X1_303 MUX2X1_303/A MUX2X1_303/B BUFX4_357/Y gnd AOI22X1_63/A vdd MUX2X1
XOAI21X1_1182 INVX1_394/Y BUFX4_255/Y NAND2X1_630/Y gnd MUX2X1_292/A vdd OAI21X1
XMUX2X1_325 MUX2X1_325/A MUX2X1_325/B BUFX4_50/Y gnd MUX2X1_325/Y vdd MUX2X1
XMUX2X1_347 MUX2X1_347/A MUX2X1_347/B BUFX4_51/Y gnd MUX2X1_347/Y vdd MUX2X1
XOAI21X1_1171 INVX1_383/Y BUFX4_233/Y NAND2X1_619/Y gnd MUX2X1_284/B vdd OAI21X1
XDFFPOSX1_750 NOR2X1_98/A CLKBUF1_100/Y AOI21X1_78/Y gnd vdd DFFPOSX1
XMUX2X1_336 MUX2X1_336/A MUX2X1_336/B BUFX4_357/Y gnd AOI22X1_70/D vdd MUX2X1
XOAI21X1_1160 INVX1_372/Y BUFX4_211/Y NAND2X1_606/Y gnd MUX2X1_275/A vdd OAI21X1
XMUX2X1_358 MUX2X1_358/A MUX2X1_358/B BUFX4_80/Y gnd MUX2X1_358/Y vdd MUX2X1
XMUX2X1_369 MUX2X1_368/Y MUX2X1_369/B BUFX4_357/Y gnd AOI22X1_77/A vdd MUX2X1
XDFFPOSX1_783 OAI21X1_597/C CLKBUF1_26/Y OAI21X1_598/Y gnd vdd DFFPOSX1
XOAI21X1_1193 INVX1_405/Y BUFX4_277/Y NAND2X1_642/Y gnd MUX2X1_301/B vdd OAI21X1
XDFFPOSX1_772 INVX1_237/A CLKBUF1_62/Y OAI21X1_576/Y gnd vdd DFFPOSX1
XDFFPOSX1_761 NOR2X1_103/A CLKBUF1_11/Y AOI21X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_794 NOR2X1_115/A CLKBUF1_74/Y AOI21X1_91/Y gnd vdd DFFPOSX1
XNAND2X1_820 BUFX4_447/Y NOR2X1_321/Y gnd NAND2X1_820/Y vdd NAND2X1
XNAND2X1_831 BUFX4_431/Y NOR2X1_331/Y gnd NAND2X1_831/Y vdd NAND2X1
XNAND2X1_864 INVX8_3/A NOR2X1_378/Y gnd NAND2X1_864/Y vdd NAND2X1
XNAND2X1_853 BUFX4_450/Y NOR2X1_368/Y gnd NAND2X1_853/Y vdd NAND2X1
XNAND2X1_842 INVX8_10/A INVX2_10/Y gnd NAND2X1_842/Y vdd NAND2X1
XFILL_4_6_0 gnd vdd FILL
XFILL_29_6_0 gnd vdd FILL
XFILL_12_5_0 gnd vdd FILL
XNOR2X1_70 NOR2X1_70/A NOR2X1_67/B gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_81 BUFX4_295/Y NOR2X1_81/B gnd NOR2X1_81/Y vdd NOR2X1
XNOR2X1_92 BUFX4_295/Y NOR2X1_52/B gnd NOR2X1_96/B vdd NOR2X1
XFILL_11_2 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd q[7] vdd BUFX2
XNAND2X1_105 BUFX4_447/Y NOR2X1_81/Y gnd OAI21X1_549/C vdd NAND2X1
XNAND2X1_116 BUFX4_431/Y NOR2X1_91/Y gnd NAND2X1_116/Y vdd NAND2X1
XNAND2X1_138 INVX8_6/A NOR2X1_122/Y gnd NAND2X1_138/Y vdd NAND2X1
XNAND2X1_149 INVX1_8/A AOI22X1_69/C gnd BUFX4_121/A vdd NAND2X1
XNAND2X1_127 INVX8_11/A INVX1_3/Y gnd OAI21X1_590/B vdd NAND2X1
XNAND2X1_3 INVX2_11/Y INVX4_3/Y gnd NAND2X1_3/Y vdd NAND2X1
XNOR2X1_160 NOR2X1_160/A NOR2X1_158/B gnd NOR2X1_160/Y vdd NOR2X1
XNOR2X1_171 NOR2X1_171/A NOR2X1_173/B gnd NOR2X1_171/Y vdd NOR2X1
XNOR2X1_182 NOR2X1_182/A NOR2X1_186/B gnd NOR2X1_182/Y vdd NOR2X1
XNOR2X1_193 NOR2X1_193/A NOR2X1_197/B gnd NOR2X1_193/Y vdd NOR2X1
XOAI21X1_622 BUFX4_456/Y INVX1_4/A MUX2X1_8/B gnd OAI21X1_622/Y vdd OAI21X1
XOAI21X1_633 BUFX4_104/Y OAI21X1_635/B OAI21X1_633/C gnd OAI21X1_633/Y vdd OAI21X1
XOAI21X1_611 INVX1_303/Y NOR2X1_122/Y NAND2X1_138/Y gnd OAI21X1_611/Y vdd OAI21X1
XOAI21X1_600 BUFX4_374/Y OAI21X1_590/B OAI21X1_599/Y gnd OAI21X1_600/Y vdd OAI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XOAI21X1_644 BUFX4_153/Y BUFX4_121/Y NAND2X1_465/B gnd OAI21X1_645/C vdd OAI21X1
XAOI21X1_8 BUFX4_374/Y NOR2X1_2/Y NOR2X1_10/Y gnd AOI21X1_8/Y vdd AOI21X1
XOAI21X1_655 INVX1_178/Y NOR2X1_145/B OAI21X1_655/C gnd OAI21X1_655/Y vdd OAI21X1
XOAI21X1_666 INVX1_435/Y NOR2X1_155/Y NAND2X1_164/Y gnd OAI21X1_666/Y vdd OAI21X1
XOAI21X1_677 BUFX4_462/Y BUFX4_67/Y INVX1_117/A gnd OAI21X1_677/Y vdd OAI21X1
XOAI21X1_699 BUFX4_146/Y BUFX4_67/Y NAND2X1_538/B gnd OAI21X1_699/Y vdd OAI21X1
XOAI21X1_688 BUFX4_285/Y NAND2X1_174/Y OAI21X1_687/Y gnd OAI21X1_688/Y vdd OAI21X1
XMUX2X1_100 MUX2X1_100/A MUX2X1_100/B BUFX4_48/Y gnd MUX2X1_100/Y vdd MUX2X1
XMUX2X1_122 MUX2X1_122/A MUX2X1_122/B BUFX4_49/Y gnd MUX2X1_122/Y vdd MUX2X1
XMUX2X1_111 MUX2X1_111/A MUX2X1_111/B INVX2_6/A gnd AOI22X1_23/A vdd MUX2X1
XMUX2X1_133 MUX2X1_133/A MUX2X1_133/B BUFX4_80/Y gnd MUX2X1_133/Y vdd MUX2X1
XMUX2X1_155 MUX2X1_155/A MUX2X1_155/B BUFX4_80/Y gnd MUX2X1_155/Y vdd MUX2X1
XMUX2X1_144 MUX2X1_143/Y MUX2X1_144/B INVX2_6/A gnd AOI22X1_30/D vdd MUX2X1
XDFFPOSX1_591 NOR2X1_69/A CLKBUF1_6/Y AOI21X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_580 INVX1_225/A CLKBUF1_83/Y OAI21X1_308/Y gnd vdd DFFPOSX1
XMUX2X1_166 MUX2X1_166/A MUX2X1_166/B BUFX4_63/Y gnd MUX2X1_166/Y vdd MUX2X1
XMUX2X1_188 MUX2X1_188/A MUX2X1_188/B BUFX4_60/Y gnd MUX2X1_189/A vdd MUX2X1
XMUX2X1_177 MUX2X1_177/A MUX2X1_177/B INVX2_6/A gnd MUX2X1_177/Y vdd MUX2X1
XMUX2X1_199 MUX2X1_199/A MUX2X1_199/B INVX4_1/A gnd MUX2X1_201/B vdd MUX2X1
XNAND2X1_672 BUFX4_233/Y NAND2X1_672/B gnd NAND2X1_672/Y vdd NAND2X1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XNAND2X1_661 BUFX4_213/Y NAND2X1_661/B gnd NAND2X1_661/Y vdd NAND2X1
XNAND2X1_650 AOI22X1_62/Y AOI22X1_63/Y gnd AOI22X1_64/D vdd NAND2X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XNAND2X1_683 BUFX4_255/Y NOR2X1_237/A gnd NAND2X1_683/Y vdd NAND2X1
XNAND2X1_694 BUFX4_273/Y NAND2X1_694/B gnd NAND2X1_694/Y vdd NAND2X1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XFILL_44_4_0 gnd vdd FILL
XDFFPOSX1_3 INVX1_126/A CLKBUF1_87/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XNOR2X1_6 NOR2X1_6/A NOR2X1_2/Y gnd NOR2X1_6/Y vdd NOR2X1
XFILL_35_4_0 gnd vdd FILL
XAOI21X1_16 BUFX4_376/Y NOR2X1_14/B NOR2X1_20/Y gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_49 BUFX4_123/Y NOR2X1_67/B NOR2X1_63/Y gnd AOI21X1_49/Y vdd AOI21X1
XAOI21X1_27 AOI21X1_3/A NOR2X1_38/B NOR2X1_35/Y gnd AOI21X1_27/Y vdd AOI21X1
XAOI21X1_38 AOI21X1_6/A NOR2X1_43/B NOR2X1_48/Y gnd AOI21X1_38/Y vdd AOI21X1
XFILL_1_4_0 gnd vdd FILL
XFILL_26_4_0 gnd vdd FILL
XOAI21X1_441 BUFX4_83/Y INVX2_4/A NAND2X1_522/B gnd OAI21X1_442/C vdd OAI21X1
XFILL_10_8_1 gnd vdd FILL
XOAI21X1_430 BUFX4_284/Y NAND2X1_92/Y OAI21X1_430/C gnd OAI21X1_430/Y vdd OAI21X1
XOAI21X1_463 BUFX4_308/Y INVX2_4/A INVX1_487/A gnd OAI21X1_464/C vdd OAI21X1
XOAI21X1_452 BUFX4_421/Y NAND2X1_94/Y OAI21X1_452/C gnd OAI21X1_452/Y vdd OAI21X1
XOAI21X1_474 BUFX4_401/Y NAND2X1_95/Y OAI21X1_474/C gnd OAI21X1_474/Y vdd OAI21X1
XOAI21X1_485 BUFX4_172/Y BUFX4_337/Y INVX1_168/A gnd OAI21X1_486/C vdd OAI21X1
XOAI21X1_496 NAND2X1_96/Y BUFX4_377/Y OAI21X1_495/Y gnd OAI21X1_496/Y vdd OAI21X1
XINVX1_505 INVX1_505/A gnd INVX1_505/Y vdd INVX1
XFILL_9_5_0 gnd vdd FILL
XNAND2X1_480 BUFX4_271/Y NOR2X1_270/A gnd NAND2X1_480/Y vdd NAND2X1
XNAND2X1_491 BUFX4_194/Y NAND2X1_491/B gnd NAND2X1_491/Y vdd NAND2X1
XFILL_17_4_0 gnd vdd FILL
XOAI21X1_1704 BUFX4_85/Y BUFX4_319/Y NAND2X1_708/B gnd OAI21X1_1705/C vdd OAI21X1
XOAI21X1_90 BUFX4_127/Y OAI21X1_96/B OAI21X1_90/C gnd OAI21X1_90/Y vdd OAI21X1
XFILL_41_2_0 gnd vdd FILL
XFILL_42_7_1 gnd vdd FILL
XOAI21X1_282 NAND2X1_66/Y BUFX4_394/Y OAI21X1_281/Y gnd OAI21X1_282/Y vdd OAI21X1
XOAI21X1_271 INVX1_415/Y NOR2X1_51/Y NAND2X1_64/Y gnd OAI21X1_271/Y vdd OAI21X1
XOAI21X1_260 INVX1_222/Y NOR2X1_41/Y NAND2X1_53/Y gnd OAI21X1_260/Y vdd OAI21X1
XOAI21X1_293 BUFX4_412/Y BUFX4_436/Y NAND2X1_378/B gnd OAI21X1_294/C vdd OAI21X1
XINVX1_313 INVX1_313/A gnd INVX1_313/Y vdd INVX1
XINVX1_324 INVX1_324/A gnd INVX1_324/Y vdd INVX1
XINVX1_302 INVX1_302/A gnd INVX1_302/Y vdd INVX1
XINVX1_335 INVX1_335/A gnd INVX1_335/Y vdd INVX1
XINVX1_346 INVX1_346/A gnd INVX1_346/Y vdd INVX1
XINVX1_368 INVX1_368/A gnd INVX1_368/Y vdd INVX1
XINVX1_357 INVX1_357/A gnd INVX1_357/Y vdd INVX1
XINVX1_379 INVX1_379/A gnd INVX1_379/Y vdd INVX1
XFILL_32_2_0 gnd vdd FILL
XFILL_33_7_1 gnd vdd FILL
XAOI21X1_306 BUFX4_400/Y NOR2X1_387/B NOR2X1_384/Y gnd AOI21X1_306/Y vdd AOI21X1
XOAI21X1_1523 BUFX4_404/Y BUFX4_93/Y INVX1_74/A gnd OAI21X1_1524/C vdd OAI21X1
XOAI21X1_1501 NOR2X1_61/B BUFX4_89/Y INVX1_393/A gnd OAI21X1_1501/Y vdd OAI21X1
XOAI21X1_1512 BUFX4_303/Y NAND2X1_835/Y OAI21X1_1512/C gnd DFFPOSX1_204/D vdd OAI21X1
XDFFPOSX1_27 INVX1_125/A CLKBUF1_87/Y DFFPOSX1_27/D gnd vdd DFFPOSX1
XDFFPOSX1_16 NOR2X1_263/A CLKBUF1_56/Y DFFPOSX1_16/D gnd vdd DFFPOSX1
XOAI21X1_1545 NOR2X1_21/B INVX2_9/A INVX1_267/A gnd OAI21X1_1546/C vdd OAI21X1
XOAI21X1_1556 BUFX4_166/Y INVX2_9/A INVX1_76/A gnd OAI21X1_1557/C vdd OAI21X1
XOAI21X1_1534 NAND2X1_836/Y BUFX4_282/Y OAI21X1_1534/C gnd DFFPOSX1_215/D vdd OAI21X1
XDFFPOSX1_38 INVX1_319/A CLKBUF1_10/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XDFFPOSX1_49 INVX1_36/A CLKBUF1_37/Y DFFPOSX1_49/D gnd vdd DFFPOSX1
XOAI21X1_1567 NAND2X1_839/Y BUFX4_282/Y OAI21X1_1567/C gnd DFFPOSX1_247/D vdd OAI21X1
XOAI21X1_1578 BUFX4_410/Y BUFX4_93/Y NAND2X1_494/B gnd OAI21X1_1578/Y vdd OAI21X1
XOAI21X1_1589 BUFX4_422/Y NAND2X1_842/Y OAI21X1_1589/C gnd OAI21X1_1589/Y vdd OAI21X1
XFILL_23_2_0 gnd vdd FILL
XFILL_24_7_1 gnd vdd FILL
XFILL_7_8_1 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XCLKBUF1_91 BUFX4_14/Y gnd CLKBUF1_91/Y vdd CLKBUF1
XCLKBUF1_80 BUFX4_18/Y gnd CLKBUF1_80/Y vdd CLKBUF1
XFILL_15_7_1 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XDFFPOSX1_409 OAI21X1_89/C CLKBUF1_4/Y OAI21X1_90/Y gnd vdd DFFPOSX1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XINVX1_132 INVX1_132/A gnd INVX1_132/Y vdd INVX1
XINVX1_176 INVX1_176/A gnd INVX1_176/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_165 INVX1_165/A gnd INVX1_165/Y vdd INVX1
XINVX1_187 INVX1_187/A gnd INVX1_187/Y vdd INVX1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XCLKBUF1_102 BUFX4_12/Y gnd CLKBUF1_102/Y vdd CLKBUF1
XBUFX4_430 d[7] gnd BUFX4_430/Y vdd BUFX4
XBUFX4_441 BUFX4_439/A gnd BUFX4_441/Y vdd BUFX4
XBUFX4_452 d[1] gnd BUFX4_452/Y vdd BUFX4
XBUFX4_463 BUFX4_467/A gnd BUFX4_463/Y vdd BUFX4
XFILL_34_1 gnd vdd FILL
XAOI21X1_103 BUFX4_395/Y NOR2X1_126/B NOR2X1_129/Y gnd AOI21X1_103/Y vdd AOI21X1
XAOI21X1_114 BUFX4_279/Y NOR2X1_139/B NOR2X1_142/Y gnd AOI21X1_114/Y vdd AOI21X1
XAOI21X1_147 BUFX4_301/Y NOR2X1_186/B NOR2X1_183/Y gnd AOI21X1_147/Y vdd AOI21X1
XAOI21X1_158 BUFX4_98/Y NOR2X1_197/B NOR2X1_196/Y gnd AOI21X1_158/Y vdd AOI21X1
XAOI21X1_125 BUFX4_127/Y NOR2X1_155/Y NOR2X1_156/Y gnd AOI21X1_125/Y vdd AOI21X1
XAOI21X1_136 BUFX4_418/Y NOR2X1_173/B NOR2X1_170/Y gnd AOI21X1_136/Y vdd AOI21X1
XAOI21X1_169 BUFX4_375/Y NOR2X1_206/B NOR2X1_209/Y gnd AOI21X1_169/Y vdd AOI21X1
XOAI21X1_1320 INVX1_447/Y NOR2X1_274/Y NAND2X1_782/Y gnd DFFPOSX1_40/D vdd OAI21X1
XOAI21X1_1331 BUFX4_460/Y BUFX4_465/Y INVX1_65/A gnd OAI21X1_1331/Y vdd OAI21X1
XOAI21X1_1364 INVX1_194/Y NOR2X1_297/Y NAND2X1_797/Y gnd DFFPOSX1_84/D vdd OAI21X1
XOAI21X1_1353 BUFX4_154/Y BUFX4_467/Y NAND2X1_483/B gnd OAI21X1_1353/Y vdd OAI21X1
XDFFPOSX1_910 NAND2X1_607/B CLKBUF1_51/Y OAI21X1_702/Y gnd vdd DFFPOSX1
XDFFPOSX1_921 MUX2X1_16/A CLKBUF1_101/Y AOI21X1_144/Y gnd vdd DFFPOSX1
XDFFPOSX1_932 INVX1_247/A CLKBUF1_18/Y OAI21X1_716/Y gnd vdd DFFPOSX1
XOAI21X1_1342 BUFX4_286/Y NAND2X1_792/Y OAI21X1_1341/Y gnd DFFPOSX1_71/D vdd OAI21X1
XOAI21X1_1386 NAND2X1_811/Y BUFX4_397/Y OAI21X1_1385/Y gnd OAI21X1_1386/Y vdd OAI21X1
XDFFPOSX1_954 NOR2X1_203/A CLKBUF1_14/Y AOI21X1_163/Y gnd vdd DFFPOSX1
XDFFPOSX1_943 NOR2X1_197/A CLKBUF1_23/Y AOI21X1_159/Y gnd vdd DFFPOSX1
XDFFPOSX1_965 INVX1_313/A CLKBUF1_67/Y OAI21X1_737/Y gnd vdd DFFPOSX1
XDFFPOSX1_976 NAND2X1_749/B CLKBUF1_67/Y OAI21X1_759/Y gnd vdd DFFPOSX1
XOAI21X1_1375 INVX1_387/Y NOR2X1_309/Y NAND2X1_808/Y gnd OAI21X1_1375/Y vdd OAI21X1
XOAI21X1_1397 BUFX4_416/Y BUFX4_463/Y NAND2X1_348/B gnd OAI21X1_1398/C vdd OAI21X1
XDFFPOSX1_998 INVX1_379/A CLKBUF1_83/Y OAI21X1_787/Y gnd vdd DFFPOSX1
XDFFPOSX1_987 NOR2X1_213/A CLKBUF1_65/Y AOI21X1_172/Y gnd vdd DFFPOSX1
XFILL_47_6_1 gnd vdd FILL
XFILL_46_1_0 gnd vdd FILL
XFILL_30_5_1 gnd vdd FILL
XDFFPOSX1_206 NAND2X1_560/B CLKBUF1_36/Y DFFPOSX1_206/D gnd vdd DFFPOSX1
XDFFPOSX1_228 INVX1_203/A CLKBUF1_52/Y DFFPOSX1_228/D gnd vdd DFFPOSX1
XDFFPOSX1_217 MUX2X1_30/A CLKBUF1_51/Y AOI21X1_271/Y gnd vdd DFFPOSX1
XDFFPOSX1_239 NOR2X1_356/A CLKBUF1_36/Y AOI21X1_284/Y gnd vdd DFFPOSX1
XNAND2X1_309 BUFX4_252/Y NAND2X1_309/B gnd OAI21X1_884/C vdd NAND2X1
XFILL_37_1_0 gnd vdd FILL
XFILL_38_6_1 gnd vdd FILL
XBUFX4_260 BUFX4_24/Y gnd BUFX4_260/Y vdd BUFX4
XBUFX4_282 INVX8_8/Y gnd BUFX4_282/Y vdd BUFX4
XBUFX4_271 BUFX4_29/Y gnd BUFX4_271/Y vdd BUFX4
XNOR2X1_342 MUX2X1_30/A NOR2X1_342/B gnd NOR2X1_342/Y vdd NOR2X1
XNOR2X1_320 INVX4_2/Y OR2X2_1/Y gnd INVX8_16/A vdd NOR2X1
XNOR2X1_331 BUFX4_390/Y NOR2X1_21/B gnd NOR2X1_331/Y vdd NOR2X1
XBUFX4_293 BUFX4_294/A gnd BUFX4_293/Y vdd BUFX4
XNOR2X1_353 NOR2X1_353/A NOR2X1_352/B gnd NOR2X1_353/Y vdd NOR2X1
XNOR2X1_386 NOR2X1_386/A NOR2X1_387/B gnd NOR2X1_386/Y vdd NOR2X1
XNOR2X1_364 NOR2X1_364/A NOR2X1_367/B gnd NOR2X1_364/Y vdd NOR2X1
XNOR2X1_375 NOR2X1_375/A NOR2X1_373/B gnd NOR2X1_375/Y vdd NOR2X1
XFILL_20_0_0 gnd vdd FILL
XFILL_21_5_1 gnd vdd FILL
XOAI21X1_815 INVX1_30/Y BUFX4_220/Y OAI21X1_815/C gnd NAND2X1_227/B vdd OAI21X1
XOAI21X1_804 INVX1_19/Y BUFX4_204/Y OAI21X1_804/C gnd AOI22X1_1/A vdd OAI21X1
XOAI21X1_837 INVX1_49/Y BUFX4_258/Y OAI21X1_837/C gnd MUX2X1_34/B vdd OAI21X1
XOAI21X1_848 INVX1_60/Y MUX2X1_2/S OAI21X1_848/C gnd MUX2X1_41/A vdd OAI21X1
XOAI21X1_826 INVX1_40/Y BUFX4_240/Y OAI21X1_826/C gnd NAND2X1_246/B vdd OAI21X1
XOAI21X1_859 INVX1_71/Y BUFX4_203/Y OAI21X1_859/C gnd MUX2X1_50/B vdd OAI21X1
XMUX2X1_304 MUX2X1_304/A MUX2X1_304/B BUFX4_2/Y gnd MUX2X1_304/Y vdd MUX2X1
XOAI21X1_1161 INVX1_373/Y BUFX4_213/Y NAND2X1_607/Y gnd MUX2X1_277/B vdd OAI21X1
XOAI21X1_1183 INVX1_395/Y BUFX4_257/Y NAND2X1_631/Y gnd MUX2X1_293/B vdd OAI21X1
XMUX2X1_348 MUX2X1_347/Y MUX2X1_348/B MUX2X1_84/S gnd MUX2X1_348/Y vdd MUX2X1
XOAI21X1_1172 INVX1_384/Y BUFX4_235/Y NAND2X1_620/Y gnd MUX2X1_284/A vdd OAI21X1
XMUX2X1_326 MUX2X1_326/A MUX2X1_326/B BUFX4_3/Y gnd MUX2X1_327/A vdd MUX2X1
XMUX2X1_315 MUX2X1_314/Y MUX2X1_315/B MUX2X1_84/S gnd MUX2X1_315/Y vdd MUX2X1
XOAI21X1_1150 INVX1_362/Y BUFX4_191/Y NAND2X1_595/Y gnd MUX2X1_268/A vdd OAI21X1
XDFFPOSX1_740 INVX1_235/A CLKBUF1_26/Y OAI21X1_556/Y gnd vdd DFFPOSX1
XMUX2X1_337 MUX2X1_337/A MUX2X1_337/B BUFX4_81/Y gnd MUX2X1_339/B vdd MUX2X1
XMUX2X1_359 MUX2X1_359/A MUX2X1_359/B BUFX4_81/Y gnd MUX2X1_359/Y vdd MUX2X1
XDFFPOSX1_751 NOR2X1_99/A CLKBUF1_4/Y AOI21X1_79/Y gnd vdd DFFPOSX1
XOAI21X1_1194 INVX1_406/Y MUX2X1_1/S NAND2X1_643/Y gnd MUX2X1_301/A vdd OAI21X1
XDFFPOSX1_773 INVX1_301/A CLKBUF1_62/Y OAI21X1_578/Y gnd vdd DFFPOSX1
XDFFPOSX1_784 NAND2X1_737/B CLKBUF1_26/Y OAI21X1_600/Y gnd vdd DFFPOSX1
XDFFPOSX1_762 NOR2X1_104/A CLKBUF1_27/Y AOI21X1_82/Y gnd vdd DFFPOSX1
XNAND2X1_810 we INVX1_509/A gnd BUFX4_168/A vdd NAND2X1
XNAND2X1_821 BUFX4_329/Y NOR2X1_321/Y gnd NAND2X1_821/Y vdd NAND2X1
XDFFPOSX1_795 NOR2X1_116/A CLKBUF1_62/Y AOI21X1_92/Y gnd vdd DFFPOSX1
XNAND2X1_843 INVX8_11/A INVX2_10/Y gnd NAND2X1_843/Y vdd NAND2X1
XNAND2X1_854 BUFX4_332/Y NOR2X1_368/Y gnd NAND2X1_854/Y vdd NAND2X1
XNAND2X1_832 INVX2_8/Y INVX4_3/Y gnd NAND2X1_832/Y vdd NAND2X1
XNAND2X1_865 INVX8_4/A NOR2X1_378/Y gnd NAND2X1_865/Y vdd NAND2X1
XFILL_4_6_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_29_6_1 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_71 NOR2X1_72/A BUFX4_455/Y gnd NOR2X1_71/Y vdd NOR2X1
XNOR2X1_82 BUFX4_295/Y BUFX4_86/Y gnd NOR2X1_90/B vdd NOR2X1
XNOR2X1_60 NOR2X1_60/A NOR2X1_55/B gnd NOR2X1_60/Y vdd NOR2X1
XNOR2X1_93 NOR2X1_93/A NOR2X1_96/B gnd NOR2X1_93/Y vdd NOR2X1
XNAND2X1_106 BUFX4_329/Y NOR2X1_81/Y gnd OAI21X1_550/C vdd NAND2X1
XNAND2X1_117 BUFX4_163/Y NOR2X1_101/Y gnd NAND2X1_117/Y vdd NAND2X1
XNAND2X1_139 INVX8_7/A NOR2X1_122/Y gnd OAI21X1_612/C vdd NAND2X1
XNAND2X1_128 BUFX4_450/Y NOR2X1_111/Y gnd OAI21X1_601/C vdd NAND2X1
XNAND2X1_4 INVX8_16/A INVX2_11/Y gnd NAND2X1_4/Y vdd NAND2X1
XNOR2X1_150 NOR2X1_150/A NOR2X1_153/B gnd NOR2X1_150/Y vdd NOR2X1
XNOR2X1_161 NOR2X1_161/A NOR2X1_158/B gnd NOR2X1_161/Y vdd NOR2X1
XNOR2X1_172 NOR2X1_172/A NOR2X1_173/B gnd NOR2X1_172/Y vdd NOR2X1
XNOR2X1_183 NOR2X1_183/A NOR2X1_186/B gnd NOR2X1_183/Y vdd NOR2X1
XNOR2X1_194 NOR2X1_194/A NOR2X1_197/B gnd NOR2X1_194/Y vdd NOR2X1
XOAI21X1_623 BUFX4_126/Y OAI21X1_635/B OAI21X1_622/Y gnd OAI21X1_623/Y vdd OAI21X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XOAI21X1_612 INVX1_367/Y NOR2X1_122/Y OAI21X1_612/C gnd OAI21X1_612/Y vdd OAI21X1
XOAI21X1_601 INVX1_110/Y NOR2X1_111/Y OAI21X1_601/C gnd OAI21X1_601/Y vdd OAI21X1
XOAI21X1_634 BUFX4_456/Y BUFX4_121/Y INVX1_433/A gnd OAI21X1_634/Y vdd OAI21X1
XOAI21X1_645 BUFX4_299/Y OAI21X1_651/B OAI21X1_645/C gnd OAI21X1_645/Y vdd OAI21X1
XOAI21X1_656 INVX1_242/Y NOR2X1_145/B OAI21X1_656/C gnd OAI21X1_656/Y vdd OAI21X1
XOAI21X1_667 INVX1_499/Y NOR2X1_155/Y OAI21X1_667/C gnd OAI21X1_667/Y vdd OAI21X1
XOAI21X1_678 BUFX4_426/Y NAND2X1_174/Y OAI21X1_677/Y gnd OAI21X1_678/Y vdd OAI21X1
XOAI21X1_689 BUFX4_462/Y BUFX4_66/Y INVX1_501/A gnd OAI21X1_690/C vdd OAI21X1
XAOI21X1_9 AOI21X1_1/A NOR2X1_14/B NOR2X1_13/Y gnd AOI21X1_9/Y vdd AOI21X1
XMUX2X1_101 MUX2X1_101/A MUX2X1_101/B BUFX4_1/Y gnd MUX2X1_101/Y vdd MUX2X1
XMUX2X1_112 MUX2X1_112/A MUX2X1_112/B BUFX4_81/Y gnd MUX2X1_112/Y vdd MUX2X1
XMUX2X1_123 MUX2X1_122/Y MUX2X1_123/B BUFX4_363/Y gnd MUX2X1_123/Y vdd MUX2X1
XMUX2X1_134 MUX2X1_134/A MUX2X1_134/B BUFX4_81/Y gnd MUX2X1_135/A vdd MUX2X1
XMUX2X1_156 MUX2X1_155/Y MUX2X1_154/Y BUFX4_363/Y gnd MUX2X1_156/Y vdd MUX2X1
XMUX2X1_145 MUX2X1_145/A MUX2X1_145/B BUFX4_50/Y gnd MUX2X1_147/B vdd MUX2X1
XDFFPOSX1_570 NAND2X1_309/B CLKBUF1_95/Y OAI21X1_292/Y gnd vdd DFFPOSX1
XDFFPOSX1_592 NOR2X1_70/A CLKBUF1_6/Y AOI21X1_56/Y gnd vdd DFFPOSX1
XMUX2X1_167 MUX2X1_167/A MUX2X1_167/B BUFX4_51/Y gnd MUX2X1_167/Y vdd MUX2X1
XDFFPOSX1_581 INVX1_289/A CLKBUF1_3/Y OAI21X1_309/Y gnd vdd DFFPOSX1
XMUX2X1_189 MUX2X1_189/A MUX2X1_187/Y BUFX4_363/Y gnd MUX2X1_189/Y vdd MUX2X1
XMUX2X1_178 MUX2X1_178/A MUX2X1_178/B BUFX4_80/Y gnd MUX2X1_180/B vdd MUX2X1
XNAND2X1_673 BUFX4_235/Y NOR2X1_153/A gnd NAND2X1_673/Y vdd NAND2X1
XNAND2X1_662 BUFX4_215/Y NAND2X1_662/B gnd NAND2X1_662/Y vdd NAND2X1
XNAND2X1_640 BUFX4_272/Y OAI21X1_29/C gnd NAND2X1_640/Y vdd NAND2X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XNAND2X1_651 BUFX4_193/Y NAND2X1_651/B gnd NAND2X1_651/Y vdd NAND2X1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XNAND2X1_684 AOI22X1_67/Y AOI22X1_68/Y gnd AOI22X1_69/D vdd NAND2X1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XNAND2X1_695 BUFX4_275/Y NOR2X1_330/A gnd NAND2X1_695/Y vdd NAND2X1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XFILL_44_4_1 gnd vdd FILL
XDFFPOSX1_4 INVX1_190/A CLKBUF1_23/Y DFFPOSX1_4/D gnd vdd DFFPOSX1
XNOR2X1_7 NOR2X1_7/A NOR2X1_2/Y gnd NOR2X1_7/Y vdd NOR2X1
XFILL_35_4_1 gnd vdd FILL
XAOI21X1_17 AOI21X1_1/A NOR2X1_27/B NOR2X1_23/Y gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_39 BUFX4_287/Y NOR2X1_43/B NOR2X1_49/Y gnd AOI21X1_39/Y vdd AOI21X1
XAOI21X1_28 BUFX4_304/Y NOR2X1_38/B NOR2X1_36/Y gnd AOI21X1_28/Y vdd AOI21X1
XFILL_1_4_1 gnd vdd FILL
XFILL_26_4_1 gnd vdd FILL
XOAI21X1_431 BUFX4_403/Y BUFX4_337/Y INVX1_486/A gnd OAI21X1_432/C vdd OAI21X1
XOAI21X1_420 BUFX4_419/Y NAND2X1_92/Y OAI21X1_420/C gnd OAI21X1_420/Y vdd OAI21X1
XOAI21X1_442 BUFX4_400/Y NAND2X1_93/Y OAI21X1_442/C gnd OAI21X1_442/Y vdd OAI21X1
XOAI21X1_464 BUFX4_377/Y NAND2X1_94/Y OAI21X1_464/C gnd OAI21X1_464/Y vdd OAI21X1
XOAI21X1_453 BUFX4_310/Y BUFX4_340/Y INVX1_167/A gnd OAI21X1_454/C vdd OAI21X1
XOAI21X1_475 BUFX4_370/Y BUFX4_336/Y NAND2X1_592/B gnd OAI21X1_475/Y vdd OAI21X1
XOAI21X1_486 NAND2X1_96/Y BUFX4_117/Y OAI21X1_486/C gnd OAI21X1_486/Y vdd OAI21X1
XOAI21X1_497 BUFX4_414/Y BUFX4_336/Y OAI21X1_497/C gnd OAI21X1_497/Y vdd OAI21X1
XINVX1_506 INVX1_506/A gnd INVX1_506/Y vdd INVX1
XFILL_9_5_1 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XNAND2X1_470 BUFX4_255/Y NOR2X1_183/A gnd NAND2X1_470/Y vdd NAND2X1
XNAND2X1_481 BUFX4_273/Y NOR2X1_280/A gnd NAND2X1_481/Y vdd NAND2X1
XNAND2X1_492 BUFX4_196/Y NOR2X1_346/A gnd NAND2X1_492/Y vdd NAND2X1
XFILL_17_4_1 gnd vdd FILL
XOAI21X1_1705 BUFX4_377/Y NAND2X1_872/Y OAI21X1_1705/C gnd DFFPOSX1_352/D vdd OAI21X1
XOAI21X1_80 BUFX4_298/Y OAI21X1_82/B OAI21X1_80/C gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 BUFX4_86/Y INVX2_1/A OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XFILL_41_2_1 gnd vdd FILL
XOAI21X1_250 BUFX4_394/Y NAND2X1_49/Y OAI21X1_249/Y gnd OAI21X1_250/Y vdd OAI21X1
XOAI21X1_283 BUFX4_165/Y BUFX4_437/Y INVX1_352/A gnd OAI21X1_283/Y vdd OAI21X1
XOAI21X1_272 INVX1_479/Y NOR2X1_51/Y NAND2X1_65/Y gnd OAI21X1_272/Y vdd OAI21X1
XOAI21X1_261 INVX1_286/Y NOR2X1_41/Y NAND2X1_54/Y gnd OAI21X1_261/Y vdd OAI21X1
XOAI21X1_294 BUFX4_116/Y NAND2X1_67/Y OAI21X1_294/C gnd OAI21X1_294/Y vdd OAI21X1
XINVX1_314 INVX1_314/A gnd INVX1_314/Y vdd INVX1
XINVX1_303 INVX1_303/A gnd INVX1_303/Y vdd INVX1
XINVX1_325 INVX1_325/A gnd INVX1_325/Y vdd INVX1
XINVX1_369 INVX1_369/A gnd INVX1_369/Y vdd INVX1
XINVX1_336 INVX1_336/A gnd INVX1_336/Y vdd INVX1
XINVX1_358 INVX1_358/A gnd INVX1_358/Y vdd INVX1
XINVX1_347 INVX1_347/A gnd INVX1_347/Y vdd INVX1
XAOI21X1_307 BUFX4_103/Y NOR2X1_387/B NOR2X1_385/Y gnd AOI21X1_307/Y vdd AOI21X1
XFILL_32_2_1 gnd vdd FILL
XOAI21X1_1513 BUFX4_147/Y BUFX4_92/Y NAND2X1_491/B gnd OAI21X1_1513/Y vdd OAI21X1
XOAI21X1_1502 BUFX4_282/Y NAND2X1_834/Y OAI21X1_1501/Y gnd OAI21X1_1502/Y vdd OAI21X1
XDFFPOSX1_17 NOR2X1_276/A CLKBUF1_44/Y DFFPOSX1_17/D gnd vdd DFFPOSX1
XOAI21X1_1546 NAND2X1_837/Y BUFX4_398/Y OAI21X1_1546/C gnd DFFPOSX1_229/D vdd OAI21X1
XOAI21X1_1557 NAND2X1_839/Y BUFX4_424/Y OAI21X1_1557/C gnd DFFPOSX1_242/D vdd OAI21X1
XOAI21X1_1524 NAND2X1_836/Y BUFX4_424/Y OAI21X1_1524/C gnd DFFPOSX1_210/D vdd OAI21X1
XOAI21X1_1535 BUFX4_405/Y BUFX4_94/Y INVX1_458/A gnd OAI21X1_1536/C vdd OAI21X1
XDFFPOSX1_28 INVX1_189/A CLKBUF1_23/Y DFFPOSX1_28/D gnd vdd DFFPOSX1
XDFFPOSX1_39 INVX1_383/A CLKBUF1_23/Y DFFPOSX1_39/D gnd vdd DFFPOSX1
XOAI21X1_1579 BUFX4_398/Y NAND2X1_840/Y OAI21X1_1578/Y gnd OAI21X1_1579/Y vdd OAI21X1
XOAI21X1_1568 BUFX4_171/Y BUFX4_93/Y INVX1_460/A gnd OAI21X1_1569/C vdd OAI21X1
XFILL_23_2_1 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XCLKBUF1_81 BUFX4_18/Y gnd CLKBUF1_81/Y vdd CLKBUF1
XCLKBUF1_70 BUFX4_15/Y gnd CLKBUF1_70/Y vdd CLKBUF1
XCLKBUF1_92 BUFX4_9/Y gnd CLKBUF1_92/Y vdd CLKBUF1
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XINVX1_144 INVX1_144/A gnd INVX1_144/Y vdd INVX1
XINVX1_166 INVX1_166/A gnd INVX1_166/Y vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XINVX1_177 INVX1_177/A gnd INVX1_177/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XBUFX4_420 INVX8_3/Y gnd BUFX4_420/Y vdd BUFX4
XBUFX4_431 d[7] gnd BUFX4_431/Y vdd BUFX4
XBUFX4_464 BUFX4_467/A gnd INVX2_7/A vdd BUFX4
XBUFX4_442 BUFX4_439/A gnd BUFX4_442/Y vdd BUFX4
XBUFX4_453 d[1] gnd BUFX4_453/Y vdd BUFX4
XFILL_27_1 gnd vdd FILL
XAOI21X1_104 BUFX4_96/Y NOR2X1_126/B NOR2X1_130/Y gnd AOI21X1_104/Y vdd AOI21X1
XAOI21X1_115 BUFX4_374/Y NOR2X1_139/B NOR2X1_143/Y gnd AOI21X1_115/Y vdd AOI21X1
XAOI21X1_126 BUFX4_126/Y NOR2X1_158/B NOR2X1_158/Y gnd AOI21X1_126/Y vdd AOI21X1
XAOI21X1_137 BUFX4_114/Y NOR2X1_173/B NOR2X1_171/Y gnd AOI21X1_137/Y vdd AOI21X1
XAOI21X1_148 BUFX4_402/Y NOR2X1_186/B NOR2X1_184/Y gnd AOI21X1_148/Y vdd AOI21X1
XAOI21X1_159 BUFX4_285/Y NOR2X1_197/B NOR2X1_197/Y gnd AOI21X1_159/Y vdd AOI21X1
XOAI21X1_1310 INVX1_318/Y NOR2X1_264/Y NAND2X1_771/Y gnd DFFPOSX1_6/D vdd OAI21X1
XOAI21X1_1321 INVX1_36/Y NOR2X1_284/Y NAND2X1_783/Y gnd DFFPOSX1_49/D vdd OAI21X1
XOAI21X1_1332 BUFX4_420/Y NAND2X1_792/Y OAI21X1_1331/Y gnd DFFPOSX1_66/D vdd OAI21X1
XOAI21X1_1354 BUFX4_397/Y NAND2X1_793/Y OAI21X1_1353/Y gnd DFFPOSX1_77/D vdd OAI21X1
XOAI21X1_1365 INVX1_258/Y NOR2X1_297/Y NAND2X1_798/Y gnd DFFPOSX1_85/D vdd OAI21X1
XOAI21X1_1343 BUFX4_460/Y INVX2_7/A INVX1_449/A gnd OAI21X1_1344/C vdd OAI21X1
XDFFPOSX1_933 INVX1_311/A CLKBUF1_86/Y OAI21X1_717/Y gnd vdd DFFPOSX1
XDFFPOSX1_911 NAND2X1_676/B CLKBUF1_9/Y OAI21X1_704/Y gnd vdd DFFPOSX1
XDFFPOSX1_922 NOR2X1_181/A CLKBUF1_21/Y AOI21X1_145/Y gnd vdd DFFPOSX1
XDFFPOSX1_900 INVX1_245/A CLKBUF1_51/Y OAI21X1_682/Y gnd vdd DFFPOSX1
XDFFPOSX1_955 NOR2X1_204/A CLKBUF1_86/Y AOI21X1_164/Y gnd vdd DFFPOSX1
XDFFPOSX1_944 NOR2X1_198/A CLKBUF1_9/Y AOI21X1_160/Y gnd vdd DFFPOSX1
XDFFPOSX1_966 INVX1_377/A CLKBUF1_69/Y OAI21X1_739/Y gnd vdd DFFPOSX1
XOAI21X1_1376 INVX1_451/Y NOR2X1_309/Y NAND2X1_809/Y gnd OAI21X1_1376/Y vdd OAI21X1
XOAI21X1_1387 BUFX4_166/Y BUFX4_466/Y INVX1_324/A gnd OAI21X1_1387/Y vdd OAI21X1
XOAI21X1_1398 BUFX4_112/Y NAND2X1_812/Y OAI21X1_1398/C gnd OAI21X1_1398/Y vdd OAI21X1
XDFFPOSX1_999 INVX1_443/A CLKBUF1_85/Y OAI21X1_789/Y gnd vdd DFFPOSX1
XDFFPOSX1_977 MUX2X1_23/B CLKBUF1_65/Y OAI21X1_761/Y gnd vdd DFFPOSX1
XDFFPOSX1_988 NOR2X1_214/A CLKBUF1_88/Y AOI21X1_173/Y gnd vdd DFFPOSX1
XFILL_46_1_1 gnd vdd FILL
XDFFPOSX1_207 NAND2X1_629/B CLKBUF1_5/Y DFFPOSX1_207/D gnd vdd DFFPOSX1
XDFFPOSX1_218 NOR2X1_343/A CLKBUF1_5/Y AOI21X1_272/Y gnd vdd DFFPOSX1
XDFFPOSX1_229 INVX1_267/A CLKBUF1_66/Y DFFPOSX1_229/D gnd vdd DFFPOSX1
XBUFX4_261 BUFX4_29/Y gnd BUFX4_261/Y vdd BUFX4
XBUFX4_272 BUFX4_29/Y gnd BUFX4_272/Y vdd BUFX4
XNOR2X1_310 INVX4_2/Y NOR2X1_275/B gnd INVX8_15/A vdd NOR2X1
XBUFX4_250 BUFX4_27/Y gnd BUFX4_250/Y vdd BUFX4
XFILL_37_1_1 gnd vdd FILL
XNOR2X1_343 NOR2X1_343/A NOR2X1_342/B gnd NOR2X1_343/Y vdd NOR2X1
XBUFX4_283 INVX8_8/Y gnd BUFX4_283/Y vdd BUFX4
XNOR2X1_332 BUFX4_389/Y BUFX4_371/Y gnd NOR2X1_338/B vdd NOR2X1
XNOR2X1_321 BUFX4_389/Y NOR2X1_41/B gnd NOR2X1_321/Y vdd NOR2X1
XBUFX4_294 BUFX4_294/A gnd INVX1_2/A vdd BUFX4
XNOR2X1_354 NOR2X1_354/A NOR2X1_352/B gnd NOR2X1_354/Y vdd NOR2X1
XNOR2X1_365 NOR2X1_365/A NOR2X1_367/B gnd NOR2X1_365/Y vdd NOR2X1
XNOR2X1_376 NOR2X1_376/A NOR2X1_373/B gnd NOR2X1_376/Y vdd NOR2X1
XNOR2X1_387 NOR2X1_387/A NOR2X1_387/B gnd NOR2X1_387/Y vdd NOR2X1
XOAI21X1_805 INVX1_20/Y BUFX4_206/Y OAI21X1_805/C gnd AOI22X1_1/D vdd OAI21X1
XOAI21X1_838 INVX1_50/Y BUFX4_260/Y NAND2X1_260/Y gnd MUX2X1_34/A vdd OAI21X1
XOAI21X1_849 INVX1_61/Y MUX2X1_5/S NAND2X1_272/Y gnd MUX2X1_43/B vdd OAI21X1
XFILL_20_0_1 gnd vdd FILL
XOAI21X1_816 INVX1_31/Y BUFX4_222/Y OAI21X1_816/C gnd AOI22X1_5/A vdd OAI21X1
XOAI21X1_827 OAI21X1_827/A OAI21X1_827/B BUFX4_155/Y gnd NAND3X1_5/B vdd OAI21X1
XMUX2X1_305 MUX2X1_305/A MUX2X1_305/B BUFX4_33/Y gnd MUX2X1_306/A vdd MUX2X1
XOAI21X1_1140 INVX1_352/Y BUFX4_270/Y NAND2X1_585/Y gnd MUX2X1_260/A vdd OAI21X1
XOAI21X1_1162 INVX1_374/Y BUFX4_215/Y NAND2X1_608/Y gnd MUX2X1_277/A vdd OAI21X1
XMUX2X1_327 MUX2X1_327/A MUX2X1_325/Y MUX2X1_96/S gnd MUX2X1_327/Y vdd MUX2X1
XDFFPOSX1_730 NOR2X1_84/A CLKBUF1_33/Y AOI21X1_66/Y gnd vdd DFFPOSX1
XOAI21X1_1151 INVX1_363/Y BUFX4_193/Y NAND2X1_596/Y gnd MUX2X1_269/B vdd OAI21X1
XMUX2X1_316 MUX2X1_316/A MUX2X1_316/B BUFX4_82/Y gnd MUX2X1_318/B vdd MUX2X1
XDFFPOSX1_741 INVX1_299/A CLKBUF1_77/Y OAI21X1_557/Y gnd vdd DFFPOSX1
XMUX2X1_338 MUX2X1_338/A MUX2X1_338/B BUFX4_82/Y gnd MUX2X1_339/A vdd MUX2X1
XOAI21X1_1173 INVX1_385/Y BUFX4_237/Y NAND2X1_621/Y gnd MUX2X1_286/B vdd OAI21X1
XOAI21X1_1184 INVX1_396/Y BUFX4_259/Y NAND2X1_632/Y gnd MUX2X1_293/A vdd OAI21X1
XMUX2X1_349 MUX2X1_349/A MUX2X1_349/B BUFX4_4/Y gnd MUX2X1_349/Y vdd MUX2X1
XDFFPOSX1_774 INVX1_365/A CLKBUF1_100/Y OAI21X1_580/Y gnd vdd DFFPOSX1
XDFFPOSX1_763 NOR2X1_105/A CLKBUF1_4/Y AOI21X1_83/Y gnd vdd DFFPOSX1
XOAI21X1_1195 INVX1_407/Y MUX2X1_4/S NAND2X1_644/Y gnd MUX2X1_302/B vdd OAI21X1
XDFFPOSX1_752 NOR2X1_100/A CLKBUF1_13/Y AOI21X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_785 MUX2X1_2/B CLKBUF1_74/Y AOI21X1_89/Y gnd vdd DFFPOSX1
XNAND2X1_822 BUFX4_139/Y NOR2X1_321/Y gnd NAND2X1_822/Y vdd NAND2X1
XDFFPOSX1_796 NOR2X1_117/A CLKBUF1_62/Y AOI21X1_93/Y gnd vdd DFFPOSX1
XNAND2X1_800 BUFX4_137/Y NOR2X1_297/Y gnd NAND2X1_800/Y vdd NAND2X1
XNAND2X1_811 INVX2_7/Y INVX4_3/Y gnd NAND2X1_811/Y vdd NAND2X1
XNAND2X1_844 BUFX4_162/Y NOR2X1_358/Y gnd NAND2X1_844/Y vdd NAND2X1
XNAND2X1_855 BUFX4_142/Y NOR2X1_368/Y gnd NAND2X1_855/Y vdd NAND2X1
XNAND2X1_833 INVX8_16/A INVX2_8/Y gnd NAND2X1_833/Y vdd NAND2X1
XNAND2X1_866 INVX8_5/A NOR2X1_378/Y gnd NAND2X1_866/Y vdd NAND2X1
XFILL_3_1_1 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_40_8_0 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XFILL_19_1_1 gnd vdd FILL
XNOR2X1_61 NOR2X1_61/A NOR2X1_61/B gnd NOR2X1_61/Y vdd NOR2X1
XNOR2X1_72 NOR2X1_72/A NOR2X1_72/B gnd NOR2X1_77/B vdd NOR2X1
XNOR2X1_50 NOR2X1_50/A NOR2X1_43/B gnd NOR2X1_50/Y vdd NOR2X1
XNOR2X1_83 NOR2X1_83/A NOR2X1_90/B gnd NOR2X1_83/Y vdd NOR2X1
XNOR2X1_94 NOR2X1_94/A NOR2X1_96/B gnd NOR2X1_94/Y vdd NOR2X1
XFILL_31_8_0 gnd vdd FILL
XNAND2X1_107 BUFX4_139/Y NOR2X1_81/Y gnd OAI21X1_551/C vdd NAND2X1
XNAND2X1_129 BUFX4_332/Y NOR2X1_111/Y gnd OAI21X1_602/C vdd NAND2X1
XNAND2X1_118 BUFX4_449/Y NOR2X1_101/Y gnd OAI21X1_562/C vdd NAND2X1
XNAND2X1_5 BUFX4_320/Y NAND2X1_5/B gnd BUFX4_178/A vdd NAND2X1
XNOR2X1_151 NOR2X1_151/A NOR2X1_153/B gnd NOR2X1_151/Y vdd NOR2X1
XNOR2X1_140 NOR2X1_140/A NOR2X1_139/B gnd NOR2X1_140/Y vdd NOR2X1
XMUX2X1_90 MUX2X1_89/Y MUX2X1_88/Y BUFX4_363/Y gnd MUX2X1_90/Y vdd MUX2X1
XNOR2X1_173 NOR2X1_173/A NOR2X1_173/B gnd NOR2X1_173/Y vdd NOR2X1
XNOR2X1_162 NOR2X1_162/A NOR2X1_158/B gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_184 NOR2X1_184/A NOR2X1_186/B gnd NOR2X1_184/Y vdd NOR2X1
XNOR2X1_195 NOR2X1_195/A NOR2X1_197/B gnd NOR2X1_195/Y vdd NOR2X1
XFILL_22_8_0 gnd vdd FILL
XOAI21X1_624 BUFX4_456/Y BUFX4_120/Y INVX1_113/A gnd OAI21X1_624/Y vdd OAI21X1
XOAI21X1_613 INVX1_431/Y NOR2X1_122/Y OAI21X1_613/C gnd OAI21X1_613/Y vdd OAI21X1
XOAI21X1_602 INVX1_174/Y NOR2X1_111/Y OAI21X1_602/C gnd OAI21X1_602/Y vdd OAI21X1
XOAI21X1_635 BUFX4_287/Y OAI21X1_635/B OAI21X1_634/Y gnd OAI21X1_635/Y vdd OAI21X1
XOAI21X1_646 BUFX4_153/Y BUFX4_120/Y NAND2X1_534/B gnd OAI21X1_647/C vdd OAI21X1
XOAI21X1_657 INVX1_306/Y NOR2X1_145/B NAND2X1_155/Y gnd OAI21X1_657/Y vdd OAI21X1
XOAI21X1_679 BUFX4_462/Y BUFX4_66/Y INVX1_181/A gnd OAI21X1_679/Y vdd OAI21X1
XOAI21X1_668 INVX1_116/Y NOR2X1_166/Y OAI21X1_668/C gnd OAI21X1_668/Y vdd OAI21X1
XMUX2X1_102 MUX2X1_101/Y MUX2X1_100/Y MUX2X1_69/S gnd MUX2X1_102/Y vdd MUX2X1
XMUX2X1_113 MUX2X1_113/A MUX2X1_113/B BUFX4_82/Y gnd MUX2X1_114/A vdd MUX2X1
XMUX2X1_135 MUX2X1_135/A MUX2X1_133/Y MUX2X1_69/S gnd MUX2X1_135/Y vdd MUX2X1
XMUX2X1_124 MUX2X1_124/A MUX2X1_124/B BUFX4_2/Y gnd MUX2X1_124/Y vdd MUX2X1
XMUX2X1_146 MUX2X1_146/A MUX2X1_146/B BUFX4_3/Y gnd MUX2X1_147/A vdd MUX2X1
XDFFPOSX1_571 NAND2X1_378/B CLKBUF1_11/Y OAI21X1_294/Y gnd vdd DFFPOSX1
XMUX2X1_179 MUX2X1_179/A MUX2X1_179/B BUFX4_81/Y gnd MUX2X1_180/A vdd MUX2X1
XMUX2X1_168 MUX2X1_167/Y MUX2X1_166/Y MUX2X1_69/S gnd MUX2X1_168/Y vdd MUX2X1
XDFFPOSX1_582 INVX1_353/A CLKBUF1_83/Y OAI21X1_310/Y gnd vdd DFFPOSX1
XMUX2X1_157 MUX2X1_157/A MUX2X1_157/B BUFX4_81/Y gnd MUX2X1_157/Y vdd MUX2X1
XDFFPOSX1_560 NOR2X1_60/A CLKBUF1_41/Y AOI21X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_593 INVX1_50/A CLKBUF1_28/Y OAI21X1_314/Y gnd vdd DFFPOSX1
XNAND2X1_630 BUFX4_254/Y NOR2X1_348/A gnd NAND2X1_630/Y vdd NAND2X1
XNAND2X1_641 BUFX4_274/Y OAI21X1_61/C gnd NAND2X1_641/Y vdd NAND2X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XNAND2X1_663 BUFX4_217/Y OAI21X1_541/C gnd NAND2X1_663/Y vdd NAND2X1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XNAND2X1_652 BUFX4_195/Y NOR2X1_49/A gnd NAND2X1_652/Y vdd NAND2X1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XNAND2X1_685 AOI22X1_64/Y AOI22X1_69/Y gnd NAND2X1_685/Y vdd NAND2X1
XNAND2X1_696 BUFX4_277/Y NOR2X1_340/A gnd NAND2X1_696/Y vdd NAND2X1
XNAND2X1_674 BUFX4_237/Y NOR2X1_164/A gnd NAND2X1_674/Y vdd NAND2X1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XDFFPOSX1_5 INVX1_254/A CLKBUF1_86/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XFILL_13_8_0 gnd vdd FILL
XNOR2X1_8 NOR2X1_8/A NOR2X1_2/Y gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 BUFX4_423/Y NOR2X1_27/B NOR2X1_24/Y gnd AOI21X1_18/Y vdd AOI21X1
XAOI21X1_29 BUFX4_395/Y NOR2X1_38/B NOR2X1_37/Y gnd AOI21X1_29/Y vdd AOI21X1
XOAI21X1_432 BUFX4_377/Y NAND2X1_92/Y OAI21X1_432/C gnd OAI21X1_432/Y vdd OAI21X1
XOAI21X1_421 BUFX4_403/Y NOR2X1_72/A INVX1_166/A gnd OAI21X1_422/C vdd OAI21X1
XOAI21X1_410 INVX1_101/Y NOR2X1_71/Y NAND2X1_85/Y gnd OAI21X1_410/Y vdd OAI21X1
XOAI21X1_443 BUFX4_83/Y BUFX4_341/Y NAND2X1_591/B gnd OAI21X1_444/C vdd OAI21X1
XOAI21X1_454 BUFX4_109/Y NAND2X1_94/Y OAI21X1_454/C gnd OAI21X1_454/Y vdd OAI21X1
XOAI21X1_465 BUFX4_370/Y BUFX4_336/Y NAND2X1_265/B gnd OAI21X1_465/Y vdd OAI21X1
XOAI21X1_487 BUFX4_169/Y BUFX4_342/Y INVX1_232/A gnd OAI21X1_488/C vdd OAI21X1
XOAI21X1_476 BUFX4_101/Y NAND2X1_95/Y OAI21X1_475/Y gnd OAI21X1_476/Y vdd OAI21X1
XOAI21X1_498 BUFX4_124/Y NAND2X1_97/Y OAI21X1_497/Y gnd OAI21X1_498/Y vdd OAI21X1
XINVX1_507 INVX1_507/A gnd INVX1_507/Y vdd INVX1
XDFFPOSX1_390 INVX1_341/A CLKBUF1_77/Y OAI21X1_70/Y gnd vdd DFFPOSX1
XFILL_8_0_1 gnd vdd FILL
XNAND2X1_471 BUFX4_257/Y NOR2X1_194/A gnd NAND2X1_471/Y vdd NAND2X1
XNAND2X1_460 AOI22X1_35/Y AOI22X1_36/Y gnd AOI22X1_39/A vdd NAND2X1
XNAND2X1_493 INVX8_1/A NOR2X1_354/A gnd NAND2X1_493/Y vdd NAND2X1
XNAND2X1_482 BUFX4_275/Y NOR2X1_290/A gnd NAND2X1_482/Y vdd NAND2X1
XFILL_45_7_0 gnd vdd FILL
XFILL_36_7_0 gnd vdd FILL
XOAI21X1_81 NOR2X1_41/B NOR2X1_2/A INVX1_278/A gnd OAI21X1_82/C vdd OAI21X1
XOAI21X1_70 INVX1_341/Y NOR2X1_1/Y NAND2X1_11/Y gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_92 BUFX4_425/Y OAI21X1_96/B OAI21X1_91/Y gnd OAI21X1_92/Y vdd OAI21X1
XFILL_2_7_0 gnd vdd FILL
XFILL_27_7_0 gnd vdd FILL
XOAI21X1_240 BUFX4_379/Y NAND2X1_48/Y OAI21X1_239/Y gnd OAI21X1_240/Y vdd OAI21X1
XFILL_10_6_0 gnd vdd FILL
XOAI21X1_273 BUFX4_165/Y BUFX4_437/Y INVX1_48/A gnd OAI21X1_274/C vdd OAI21X1
XOAI21X1_262 INVX1_350/Y NOR2X1_41/Y NAND2X1_55/Y gnd OAI21X1_262/Y vdd OAI21X1
XOAI21X1_251 BUFX4_150/Y INVX2_2/A OAI21X1_251/C gnd OAI21X1_252/C vdd OAI21X1
XOAI21X1_284 NAND2X1_66/Y BUFX4_97/Y OAI21X1_283/Y gnd OAI21X1_284/Y vdd OAI21X1
XOAI21X1_295 BUFX4_411/Y BUFX4_433/Y NAND2X1_447/B gnd OAI21X1_295/Y vdd OAI21X1
XINVX1_304 INVX1_304/A gnd INVX1_304/Y vdd INVX1
XINVX1_315 INVX1_315/A gnd INVX1_315/Y vdd INVX1
XINVX1_326 INVX1_326/A gnd INVX1_326/Y vdd INVX1
XINVX1_359 INVX1_359/A gnd INVX1_359/Y vdd INVX1
XINVX1_337 INVX1_337/A gnd INVX1_337/Y vdd INVX1
XINVX1_348 INVX1_348/A gnd INVX1_348/Y vdd INVX1
XNAND2X1_290 BUFX4_216/Y NOR2X1_361/A gnd OAI21X1_866/C vdd NAND2X1
XFILL_18_7_0 gnd vdd FILL
XAOI21X1_308 BUFX4_284/Y NOR2X1_387/B NOR2X1_386/Y gnd AOI21X1_308/Y vdd AOI21X1
XOAI21X1_1514 BUFX4_402/Y NAND2X1_835/Y OAI21X1_1513/Y gnd OAI21X1_1514/Y vdd OAI21X1
XOAI21X1_1503 NOR2X1_61/B BUFX4_94/Y INVX1_457/A gnd OAI21X1_1503/Y vdd OAI21X1
XDFFPOSX1_18 NOR2X1_277/A CLKBUF1_2/Y DFFPOSX1_18/D gnd vdd DFFPOSX1
XOAI21X1_1525 BUFX4_405/Y BUFX4_91/Y INVX1_138/A gnd OAI21X1_1525/Y vdd OAI21X1
XOAI21X1_1547 BUFX4_312/Y BUFX4_95/Y INVX1_331/A gnd OAI21X1_1547/Y vdd OAI21X1
XOAI21X1_1536 NAND2X1_836/Y BUFX4_375/Y OAI21X1_1536/C gnd DFFPOSX1_216/D vdd OAI21X1
XDFFPOSX1_29 INVX1_253/A CLKBUF1_18/Y DFFPOSX1_29/D gnd vdd DFFPOSX1
XOAI21X1_1558 BUFX4_166/Y BUFX4_92/Y INVX1_140/A gnd OAI21X1_1559/C vdd OAI21X1
XOAI21X1_1569 NAND2X1_839/Y BUFX4_380/Y OAI21X1_1569/C gnd DFFPOSX1_248/D vdd OAI21X1
XCLKBUF1_60 BUFX4_10/Y gnd CLKBUF1_60/Y vdd CLKBUF1
XCLKBUF1_82 BUFX4_18/Y gnd CLKBUF1_82/Y vdd CLKBUF1
XCLKBUF1_71 BUFX4_11/Y gnd CLKBUF1_71/Y vdd CLKBUF1
XCLKBUF1_93 BUFX4_11/Y gnd CLKBUF1_93/Y vdd CLKBUF1
XFILL_42_5_0 gnd vdd FILL
XINVX1_101 INVX1_101/A gnd INVX1_101/Y vdd INVX1
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XINVX1_123 INVX1_123/A gnd INVX1_123/Y vdd INVX1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_167 INVX1_167/A gnd INVX1_167/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XINVX1_189 INVX1_189/A gnd INVX1_189/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XBUFX4_421 INVX8_3/Y gnd BUFX4_421/Y vdd BUFX4
XBUFX4_410 INVX8_16/Y gnd BUFX4_410/Y vdd BUFX4
XBUFX4_465 BUFX4_467/A gnd BUFX4_465/Y vdd BUFX4
XBUFX4_443 BUFX4_439/A gnd BUFX4_443/Y vdd BUFX4
XBUFX4_454 INVX8_10/Y gnd BUFX4_454/Y vdd BUFX4
XBUFX4_432 BUFX4_436/A gnd BUFX4_432/Y vdd BUFX4
XFILL_33_5_0 gnd vdd FILL
XAOI21X1_105 BUFX4_279/Y NOR2X1_126/B NOR2X1_131/Y gnd AOI21X1_105/Y vdd AOI21X1
XAOI21X1_138 BUFX4_299/Y NOR2X1_173/B NOR2X1_172/Y gnd AOI21X1_138/Y vdd AOI21X1
XAOI21X1_149 BUFX4_98/Y NOR2X1_186/B NOR2X1_185/Y gnd AOI21X1_149/Y vdd AOI21X1
XAOI21X1_116 BUFX4_126/Y NOR2X1_145/B NOR2X1_145/Y gnd AOI21X1_116/Y vdd AOI21X1
XAOI21X1_127 BUFX4_418/Y NOR2X1_158/B NOR2X1_159/Y gnd AOI21X1_127/Y vdd AOI21X1
XOAI21X1_1311 INVX1_382/Y NOR2X1_264/Y NAND2X1_772/Y gnd DFFPOSX1_7/D vdd OAI21X1
XOAI21X1_1300 INVX1_189/Y NOR2X1_254/Y NAND2X1_759/Y gnd DFFPOSX1_28/D vdd OAI21X1
XOAI21X1_1322 INVX1_64/Y NOR2X1_284/Y NAND2X1_784/Y gnd DFFPOSX1_50/D vdd OAI21X1
XOAI21X1_1333 BUFX4_460/Y BUFX4_465/Y INVX1_129/A gnd OAI21X1_1333/Y vdd OAI21X1
XOAI21X1_1344 BUFX4_373/Y NAND2X1_792/Y OAI21X1_1344/C gnd DFFPOSX1_72/D vdd OAI21X1
XDFFPOSX1_923 NOR2X1_182/A CLKBUF1_86/Y AOI21X1_146/Y gnd vdd DFFPOSX1
XDFFPOSX1_912 NAND2X1_745/B CLKBUF1_9/Y OAI21X1_706/Y gnd vdd DFFPOSX1
XDFFPOSX1_901 INVX1_309/A CLKBUF1_9/Y OAI21X1_684/Y gnd vdd DFFPOSX1
XOAI21X1_1355 BUFX4_154/Y INVX2_7/A NAND2X1_552/B gnd OAI21X1_1355/Y vdd OAI21X1
XOAI21X1_1377 BUFX4_168/Y BUFX4_468/Y INVX1_40/A gnd OAI21X1_1377/Y vdd OAI21X1
XDFFPOSX1_945 MUX2X1_19/B CLKBUF1_86/Y AOI21X1_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_956 NOR2X1_205/A CLKBUF1_101/Y AOI21X1_165/Y gnd vdd DFFPOSX1
XDFFPOSX1_934 INVX1_375/A CLKBUF1_14/Y OAI21X1_718/Y gnd vdd DFFPOSX1
XOAI21X1_1388 NAND2X1_811/Y BUFX4_99/Y OAI21X1_1387/Y gnd OAI21X1_1388/Y vdd OAI21X1
XOAI21X1_1366 INVX1_322/Y NOR2X1_297/Y NAND2X1_799/Y gnd DFFPOSX1_86/D vdd OAI21X1
XOAI21X1_1399 BUFX4_416/Y INVX2_7/A NAND2X1_417/B gnd OAI21X1_1400/C vdd OAI21X1
XDFFPOSX1_978 INVX1_122/A CLKBUF1_65/Y OAI21X1_763/Y gnd vdd DFFPOSX1
XDFFPOSX1_989 NOR2X1_215/A CLKBUF1_65/Y AOI21X1_174/Y gnd vdd DFFPOSX1
XDFFPOSX1_967 INVX1_441/A CLKBUF1_59/Y OAI21X1_741/Y gnd vdd DFFPOSX1
XFILL_24_5_0 gnd vdd FILL
XFILL_7_6_0 gnd vdd FILL
XFILL_15_5_0 gnd vdd FILL
XDFFPOSX1_219 NOR2X1_344/A CLKBUF1_76/Y AOI21X1_273/Y gnd vdd DFFPOSX1
XDFFPOSX1_208 NAND2X1_698/B CLKBUF1_35/Y DFFPOSX1_208/D gnd vdd DFFPOSX1
XBUFX4_240 BUFX4_27/Y gnd BUFX4_240/Y vdd BUFX4
XNOR2X1_300 NOR2X1_300/A NOR2X1_303/B gnd NOR2X1_300/Y vdd NOR2X1
XBUFX4_273 BUFX4_30/Y gnd BUFX4_273/Y vdd BUFX4
XBUFX4_251 BUFX4_30/Y gnd BUFX4_251/Y vdd BUFX4
XBUFX4_262 BUFX4_23/Y gnd BUFX4_262/Y vdd BUFX4
XBUFX4_284 INVX8_8/Y gnd BUFX4_284/Y vdd BUFX4
XNOR2X1_333 NOR2X1_333/A NOR2X1_338/B gnd NOR2X1_333/Y vdd NOR2X1
XNOR2X1_322 BUFX4_389/Y BUFX4_84/Y gnd NOR2X1_325/B vdd NOR2X1
XBUFX4_295 BUFX4_294/A gnd BUFX4_295/Y vdd BUFX4
XNOR2X1_311 BUFX4_466/Y BUFX4_371/Y gnd NOR2X1_315/B vdd NOR2X1
XNOR2X1_344 NOR2X1_344/A NOR2X1_342/B gnd NOR2X1_344/Y vdd NOR2X1
XNOR2X1_355 NOR2X1_355/A NOR2X1_352/B gnd NOR2X1_355/Y vdd NOR2X1
XNOR2X1_366 NOR2X1_366/A NOR2X1_367/B gnd NOR2X1_366/Y vdd NOR2X1
XNOR2X1_377 NOR2X1_377/A NOR2X1_373/B gnd NOR2X1_377/Y vdd NOR2X1
XOAI21X1_806 INVX8_1/Y OAI21X1_49/C OAI21X1_806/C gnd NAND3X1_2/A vdd OAI21X1
XOAI21X1_839 INVX1_51/Y BUFX4_262/Y NAND2X1_261/Y gnd MUX2X1_35/B vdd OAI21X1
XOAI21X1_817 INVX1_32/Y BUFX4_224/Y NAND2X1_229/Y gnd AOI22X1_5/D vdd OAI21X1
XOAI21X1_828 INVX1_41/Y BUFX4_242/Y OAI21X1_828/C gnd NAND2X1_248/B vdd OAI21X1
XOAI21X1_1130 INVX1_342/Y BUFX4_250/Y NAND2X1_574/Y gnd MUX2X1_253/A vdd OAI21X1
XDFFPOSX1_720 OAI21X1_543/C CLKBUF1_46/Y OAI21X1_544/Y gnd vdd DFFPOSX1
XOAI21X1_1163 INVX1_375/Y BUFX4_217/Y NAND2X1_609/Y gnd MUX2X1_278/B vdd OAI21X1
XOAI21X1_1141 INVX1_353/Y BUFX4_272/Y NAND2X1_586/Y gnd MUX2X1_262/B vdd OAI21X1
XMUX2X1_306 MUX2X1_306/A MUX2X1_304/Y MUX2X1_42/S gnd MUX2X1_306/Y vdd MUX2X1
XMUX2X1_328 MUX2X1_328/A MUX2X1_328/B BUFX4_34/Y gnd MUX2X1_330/B vdd MUX2X1
XDFFPOSX1_731 NOR2X1_85/A CLKBUF1_72/Y AOI21X1_67/Y gnd vdd DFFPOSX1
XOAI21X1_1152 INVX1_364/Y BUFX4_195/Y NAND2X1_597/Y gnd MUX2X1_269/A vdd OAI21X1
XMUX2X1_317 MUX2X1_317/A MUX2X1_317/B BUFX4_42/Y gnd MUX2X1_318/A vdd MUX2X1
XMUX2X1_339 MUX2X1_339/A MUX2X1_339/B MUX2X1_42/S gnd AOI22X1_71/A vdd MUX2X1
XOAI21X1_1174 INVX1_386/Y BUFX4_239/Y NAND2X1_622/Y gnd MUX2X1_286/A vdd OAI21X1
XDFFPOSX1_775 INVX1_429/A CLKBUF1_100/Y OAI21X1_582/Y gnd vdd DFFPOSX1
XDFFPOSX1_742 INVX1_363/A CLKBUF1_100/Y OAI21X1_558/Y gnd vdd DFFPOSX1
XOAI21X1_1196 INVX1_408/Y MUX2X1_8/S NAND2X1_645/Y gnd MUX2X1_302/A vdd OAI21X1
XOAI21X1_1185 INVX1_397/Y BUFX4_261/Y NAND2X1_634/Y gnd MUX2X1_295/B vdd OAI21X1
XDFFPOSX1_764 NOR2X1_106/A CLKBUF1_26/Y AOI21X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_753 INVX1_60/A CLKBUF1_48/Y OAI21X1_561/Y gnd vdd DFFPOSX1
XDFFPOSX1_786 INVX1_110/A CLKBUF1_74/Y OAI21X1_601/Y gnd vdd DFFPOSX1
XDFFPOSX1_797 NOR2X1_118/A CLKBUF1_13/Y AOI21X1_94/Y gnd vdd DFFPOSX1
XNAND2X1_801 BUFX4_428/Y NOR2X1_297/Y gnd NAND2X1_801/Y vdd NAND2X1
XNAND2X1_812 INVX8_16/A INVX2_7/Y gnd NAND2X1_812/Y vdd NAND2X1
XNAND2X1_834 INVX8_10/A INVX2_9/Y gnd NAND2X1_834/Y vdd NAND2X1
XNAND2X1_845 BUFX4_449/Y NOR2X1_358/Y gnd NAND2X1_845/Y vdd NAND2X1
XNAND2X1_823 BUFX4_430/Y NOR2X1_321/Y gnd NAND2X1_823/Y vdd NAND2X1
XNAND2X1_867 INVX8_6/A NOR2X1_378/Y gnd NAND2X1_867/Y vdd NAND2X1
XNAND2X1_856 BUFX4_445/Y NOR2X1_368/Y gnd NAND2X1_856/Y vdd NAND2X1
XFILL_40_8_1 gnd vdd FILL
XFILL_47_4_0 gnd vdd FILL
XNOR2X1_62 BUFX4_385/Y NOR2X1_2/B gnd NOR2X1_67/B vdd NOR2X1
XNOR2X1_73 NOR2X1_73/A NOR2X1_77/B gnd NOR2X1_73/Y vdd NOR2X1
XNOR2X1_40 NOR2X1_40/A NOR2X1_38/B gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_51 BUFX4_432/Y NOR2X1_51/B gnd NOR2X1_51/Y vdd NOR2X1
XNOR2X1_84 NOR2X1_84/A NOR2X1_90/B gnd NOR2X1_84/Y vdd NOR2X1
XNOR2X1_95 NOR2X1_95/A NOR2X1_96/B gnd NOR2X1_95/Y vdd NOR2X1
XFILL_31_8_1 gnd vdd FILL
XFILL_30_3_0 gnd vdd FILL
XNAND2X1_108 BUFX4_430/Y NOR2X1_81/Y gnd NAND2X1_108/Y vdd NAND2X1
XNAND2X1_119 NAND2X1_8/A NOR2X1_101/Y gnd OAI21X1_563/C vdd NAND2X1
XNAND2X1_6 INVX8_2/A NOR2X1_1/Y gnd NAND2X1_6/Y vdd NAND2X1
XFILL_38_4_0 gnd vdd FILL
XNOR2X1_141 NOR2X1_141/A NOR2X1_139/B gnd NOR2X1_141/Y vdd NOR2X1
XNOR2X1_130 NOR2X1_130/A NOR2X1_126/B gnd NOR2X1_130/Y vdd NOR2X1
XMUX2X1_80 MUX2X1_80/A MUX2X1_80/B BUFX4_35/Y gnd MUX2X1_80/Y vdd MUX2X1
XNOR2X1_152 NOR2X1_152/A NOR2X1_153/B gnd NOR2X1_152/Y vdd NOR2X1
XNOR2X1_163 NOR2X1_163/A NOR2X1_158/B gnd NOR2X1_163/Y vdd NOR2X1
XNOR2X1_185 NOR2X1_185/A NOR2X1_186/B gnd NOR2X1_185/Y vdd NOR2X1
XMUX2X1_91 MUX2X1_91/A MUX2X1_91/B BUFX4_82/Y gnd MUX2X1_91/Y vdd MUX2X1
XNOR2X1_174 NOR2X1_174/A NOR2X1_173/B gnd NOR2X1_174/Y vdd NOR2X1
XNOR2X1_196 NOR2X1_196/A NOR2X1_197/B gnd NOR2X1_196/Y vdd NOR2X1
XFILL_22_8_1 gnd vdd FILL
XFILL_21_3_0 gnd vdd FILL
XOAI21X1_614 INVX1_495/Y NOR2X1_122/Y OAI21X1_614/C gnd OAI21X1_614/Y vdd OAI21X1
XOAI21X1_603 INVX1_238/Y NOR2X1_111/Y OAI21X1_603/C gnd OAI21X1_603/Y vdd OAI21X1
XOAI21X1_647 BUFX4_396/Y OAI21X1_651/B OAI21X1_647/C gnd OAI21X1_647/Y vdd OAI21X1
XOAI21X1_636 BUFX4_456/Y BUFX4_120/Y INVX1_497/A gnd OAI21X1_637/C vdd OAI21X1
XOAI21X1_625 BUFX4_418/Y OAI21X1_635/B OAI21X1_624/Y gnd OAI21X1_625/Y vdd OAI21X1
XOAI21X1_669 INVX1_180/Y NOR2X1_166/Y NAND2X1_167/Y gnd OAI21X1_669/Y vdd OAI21X1
XOAI21X1_658 INVX1_370/Y NOR2X1_145/B NAND2X1_156/Y gnd OAI21X1_658/Y vdd OAI21X1
XMUX2X1_114 MUX2X1_114/A MUX2X1_112/Y MUX2X1_48/S gnd MUX2X1_114/Y vdd MUX2X1
XMUX2X1_103 MUX2X1_103/A MUX2X1_103/B BUFX4_32/Y gnd MUX2X1_103/Y vdd MUX2X1
XMUX2X1_136 MUX2X1_136/A MUX2X1_136/B BUFX4_82/Y gnd MUX2X1_136/Y vdd MUX2X1
XMUX2X1_125 MUX2X1_125/A MUX2X1_125/B BUFX4_33/Y gnd MUX2X1_126/A vdd MUX2X1
XMUX2X1_147 MUX2X1_147/A MUX2X1_147/B MUX2X1_48/S gnd AOI22X1_31/A vdd MUX2X1
XDFFPOSX1_550 INVX1_351/A CLKBUF1_46/Y OAI21X1_270/Y gnd vdd DFFPOSX1
XDFFPOSX1_561 INVX1_48/A CLKBUF1_80/Y OAI21X1_274/Y gnd vdd DFFPOSX1
XDFFPOSX1_572 NAND2X1_447/B CLKBUF1_95/Y OAI21X1_296/Y gnd vdd DFFPOSX1
XDFFPOSX1_583 INVX1_417/A CLKBUF1_6/Y OAI21X1_311/Y gnd vdd DFFPOSX1
XMUX2X1_169 MUX2X1_169/A MUX2X1_169/B BUFX4_4/Y gnd MUX2X1_171/B vdd MUX2X1
XMUX2X1_158 MUX2X1_158/A MUX2X1_158/B BUFX4_82/Y gnd MUX2X1_159/A vdd MUX2X1
XDFFPOSX1_594 INVX1_98/A CLKBUF1_70/Y OAI21X1_316/Y gnd vdd DFFPOSX1
XNAND2X1_620 BUFX4_234/Y NOR2X1_292/A gnd NAND2X1_620/Y vdd NAND2X1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XNAND2X1_631 BUFX4_256/Y NOR2X1_356/A gnd NAND2X1_631/Y vdd NAND2X1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XNAND2X1_642 BUFX4_276/Y NOR2X1_9/A gnd NAND2X1_642/Y vdd NAND2X1
XNAND2X1_664 BUFX4_219/Y NOR2X1_89/A gnd NAND2X1_664/Y vdd NAND2X1
XNAND2X1_653 BUFX4_197/Y NOR2X1_59/A gnd NAND2X1_653/Y vdd NAND2X1
XNAND2X1_697 MUX2X1_1/S NAND2X1_697/B gnd NAND2X1_697/Y vdd NAND2X1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XNAND2X1_686 BUFX4_257/Y NOR2X1_263/A gnd NAND2X1_686/Y vdd NAND2X1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XNAND2X1_675 BUFX4_239/Y NOR2X1_175/A gnd NAND2X1_675/Y vdd NAND2X1
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XFILL_4_4_0 gnd vdd FILL
XFILL_29_4_0 gnd vdd FILL
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XDFFPOSX1_6 INVX1_318/A CLKBUF1_90/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XFILL_13_8_1 gnd vdd FILL
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_2/Y gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 AOI21X1_3/A NOR2X1_27/B NOR2X1_25/Y gnd AOI21X1_19/Y vdd AOI21X1
XOAI21X1_400 BUFX4_303/Y NAND2X1_82/Y OAI21X1_399/Y gnd OAI21X1_400/Y vdd OAI21X1
XOAI21X1_422 BUFX4_117/Y NAND2X1_92/Y OAI21X1_422/C gnd OAI21X1_422/Y vdd OAI21X1
XOAI21X1_411 INVX1_165/Y NOR2X1_71/Y NAND2X1_86/Y gnd OAI21X1_411/Y vdd OAI21X1
XOAI21X1_433 BUFX4_83/Y BUFX4_342/Y NAND2X1_264/B gnd OAI21X1_434/C vdd OAI21X1
XOAI21X1_444 BUFX4_101/Y NAND2X1_93/Y OAI21X1_444/C gnd OAI21X1_444/Y vdd OAI21X1
XOAI21X1_455 BUFX4_310/Y BUFX4_341/Y INVX1_231/A gnd OAI21X1_456/C vdd OAI21X1
XOAI21X1_466 BUFX4_124/Y NAND2X1_95/Y OAI21X1_465/Y gnd OAI21X1_466/Y vdd OAI21X1
XOAI21X1_488 NAND2X1_96/Y BUFX4_302/Y OAI21X1_488/C gnd OAI21X1_488/Y vdd OAI21X1
XOAI21X1_477 BUFX4_368/Y BUFX4_340/Y NAND2X1_661/B gnd OAI21X1_478/C vdd OAI21X1
XOAI21X1_499 BUFX4_414/Y NOR2X1_72/A OAI21X1_499/C gnd OAI21X1_500/C vdd OAI21X1
XINVX1_508 INVX1_508/A gnd INVX1_508/Y vdd INVX1
XDFFPOSX1_380 OAI21X1_55/C CLKBUF1_8/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XDFFPOSX1_391 INVX1_405/A CLKBUF1_75/Y OAI21X1_71/Y gnd vdd DFFPOSX1
XNAND2X1_472 BUFX4_259/Y NOR2X1_205/A gnd NAND2X1_472/Y vdd NAND2X1
XNAND2X1_450 BUFX4_217/Y NAND2X1_450/B gnd NAND2X1_450/Y vdd NAND2X1
XNAND2X1_461 BUFX4_237/Y NAND2X1_461/B gnd NAND2X1_461/Y vdd NAND2X1
XNAND2X1_483 BUFX4_277/Y NAND2X1_483/B gnd NAND2X1_483/Y vdd NAND2X1
XNAND2X1_494 BUFX4_200/Y NAND2X1_494/B gnd NAND2X1_494/Y vdd NAND2X1
XFILL_45_7_1 gnd vdd FILL
XFILL_44_2_0 gnd vdd FILL
XFILL_36_7_1 gnd vdd FILL
XFILL_35_2_0 gnd vdd FILL
XOAI21X1_60 BUFX4_102/Y NAND2X1_4/Y OAI21X1_59/Y gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_71 INVX1_405/Y NOR2X1_1/Y OAI21X1_71/C gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_93 BUFX4_86/Y INVX2_1/A OAI21X1_93/C gnd OAI21X1_94/C vdd OAI21X1
XOAI21X1_82 BUFX4_399/Y OAI21X1_82/B OAI21X1_82/C gnd OAI21X1_82/Y vdd OAI21X1
XFILL_2_7_1 gnd vdd FILL
XFILL_27_7_1 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XFILL_26_2_0 gnd vdd FILL
XOAI21X1_230 BUFX4_114/Y NAND2X1_48/Y OAI21X1_229/Y gnd OAI21X1_230/Y vdd OAI21X1
XOAI21X1_241 BUFX4_154/Y BUFX4_436/Y OAI21X1_241/C gnd OAI21X1_241/Y vdd OAI21X1
XFILL_10_6_1 gnd vdd FILL
XOAI21X1_274 NAND2X1_66/Y BUFX4_126/Y OAI21X1_274/C gnd OAI21X1_274/Y vdd OAI21X1
XOAI21X1_263 INVX1_414/Y NOR2X1_41/Y NAND2X1_56/Y gnd OAI21X1_263/Y vdd OAI21X1
XOAI21X1_252 AOI21X1_6/A NAND2X1_49/Y OAI21X1_252/C gnd OAI21X1_252/Y vdd OAI21X1
XOAI21X1_285 BUFX4_165/Y BUFX4_434/Y INVX1_416/A gnd OAI21X1_285/Y vdd OAI21X1
XOAI21X1_296 BUFX4_299/Y NAND2X1_67/Y OAI21X1_295/Y gnd OAI21X1_296/Y vdd OAI21X1
XINVX1_305 INVX1_305/A gnd INVX1_305/Y vdd INVX1
XINVX1_316 INVX1_316/A gnd INVX1_316/Y vdd INVX1
XINVX1_349 INVX1_349/A gnd INVX1_349/Y vdd INVX1
XINVX1_338 INVX1_338/A gnd INVX1_338/Y vdd INVX1
XINVX1_327 INVX1_327/A gnd INVX1_327/Y vdd INVX1
XFILL_9_3_0 gnd vdd FILL
XNAND2X1_280 INVX8_1/A NAND2X1_280/B gnd NAND2X1_280/Y vdd NAND2X1
XNAND2X1_291 BUFX4_218/Y NOR2X1_371/A gnd OAI21X1_867/C vdd NAND2X1
XFILL_18_7_1 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XAOI21X1_309 BUFX4_378/Y NOR2X1_387/B NOR2X1_387/Y gnd AOI21X1_309/Y vdd AOI21X1
XOAI21X1_1504 BUFX4_375/Y NAND2X1_834/Y OAI21X1_1503/Y gnd OAI21X1_1504/Y vdd OAI21X1
XOAI21X1_1526 NAND2X1_836/Y BUFX4_115/Y OAI21X1_1525/Y gnd DFFPOSX1_211/D vdd OAI21X1
XOAI21X1_1515 BUFX4_146/Y BUFX4_94/Y NAND2X1_560/B gnd OAI21X1_1515/Y vdd OAI21X1
XOAI21X1_1548 NAND2X1_837/Y BUFX4_96/Y OAI21X1_1547/Y gnd DFFPOSX1_230/D vdd OAI21X1
XOAI21X1_1537 BUFX4_312/Y BUFX4_89/Y INVX1_15/A gnd OAI21X1_1537/Y vdd OAI21X1
XDFFPOSX1_19 NOR2X1_278/A CLKBUF1_71/Y DFFPOSX1_19/D gnd vdd DFFPOSX1
XOAI21X1_1559 NAND2X1_839/Y BUFX4_113/Y OAI21X1_1559/C gnd OAI21X1_1559/Y vdd OAI21X1
XCLKBUF1_50 BUFX4_13/Y gnd CLKBUF1_50/Y vdd CLKBUF1
XCLKBUF1_83 BUFX4_15/Y gnd CLKBUF1_83/Y vdd CLKBUF1
XCLKBUF1_72 BUFX4_9/Y gnd CLKBUF1_72/Y vdd CLKBUF1
XCLKBUF1_61 BUFX4_11/Y gnd CLKBUF1_61/Y vdd CLKBUF1
XCLKBUF1_94 BUFX4_13/Y gnd CLKBUF1_94/Y vdd CLKBUF1
XFILL_41_0_0 gnd vdd FILL
XFILL_42_5_1 gnd vdd FILL
XINVX1_102 INVX1_102/A gnd INVX1_102/Y vdd INVX1
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XINVX1_135 INVX1_135/A gnd INVX1_135/Y vdd INVX1
XINVX1_179 INVX1_179/A gnd INVX1_179/Y vdd INVX1
XBUFX4_400 INVX8_6/Y gnd BUFX4_400/Y vdd BUFX4
XBUFX4_422 INVX8_3/Y gnd BUFX4_422/Y vdd BUFX4
XBUFX4_411 INVX8_16/Y gnd BUFX4_411/Y vdd BUFX4
XBUFX4_444 d[4] gnd BUFX4_444/Y vdd BUFX4
XBUFX4_455 INVX8_10/Y gnd BUFX4_455/Y vdd BUFX4
XBUFX4_433 BUFX4_436/A gnd BUFX4_433/Y vdd BUFX4
XBUFX4_466 BUFX4_467/A gnd BUFX4_466/Y vdd BUFX4
XFILL_33_5_1 gnd vdd FILL
XAOI21X1_106 BUFX4_374/Y NOR2X1_126/B NOR2X1_132/Y gnd AOI21X1_106/Y vdd AOI21X1
XFILL_32_0_0 gnd vdd FILL
XAOI21X1_117 BUFX4_126/Y NOR2X1_153/B NOR2X1_147/Y gnd AOI21X1_117/Y vdd AOI21X1
XAOI21X1_139 BUFX4_394/Y NOR2X1_173/B NOR2X1_173/Y gnd AOI21X1_139/Y vdd AOI21X1
XAOI21X1_128 BUFX4_116/Y NOR2X1_158/B NOR2X1_160/Y gnd AOI21X1_128/Y vdd AOI21X1
XOAI21X1_1312 INVX1_446/Y NOR2X1_264/Y NAND2X1_773/Y gnd DFFPOSX1_8/D vdd OAI21X1
XOAI21X1_1301 INVX1_253/Y NOR2X1_254/Y NAND2X1_760/Y gnd DFFPOSX1_29/D vdd OAI21X1
XOAI21X1_1323 INVX1_128/Y NOR2X1_284/Y NAND2X1_785/Y gnd DFFPOSX1_51/D vdd OAI21X1
XOAI21X1_1345 BUFX4_154/Y BUFX4_467/Y DFFPOSX1_73/Q gnd OAI21X1_1345/Y vdd OAI21X1
XOAI21X1_1334 BUFX4_112/Y NAND2X1_792/Y OAI21X1_1333/Y gnd DFFPOSX1_67/D vdd OAI21X1
XDFFPOSX1_924 NOR2X1_183/A CLKBUF1_101/Y AOI21X1_147/Y gnd vdd DFFPOSX1
XDFFPOSX1_913 MUX2X1_16/B CLKBUF1_101/Y AOI21X1_143/Y gnd vdd DFFPOSX1
XDFFPOSX1_902 INVX1_373/A CLKBUF1_21/Y OAI21X1_686/Y gnd vdd DFFPOSX1
XOAI21X1_1356 BUFX4_99/Y NAND2X1_793/Y OAI21X1_1355/Y gnd DFFPOSX1_78/D vdd OAI21X1
XOAI21X1_1389 BUFX4_168/Y BUFX4_467/Y INVX1_388/A gnd OAI21X1_1389/Y vdd OAI21X1
XOAI21X1_1378 NAND2X1_811/Y BUFX4_125/Y OAI21X1_1377/Y gnd OAI21X1_1378/Y vdd OAI21X1
XDFFPOSX1_946 INVX1_120/A CLKBUF1_90/Y OAI21X1_721/Y gnd vdd DFFPOSX1
XDFFPOSX1_957 NOR2X1_206/A CLKBUF1_18/Y AOI21X1_166/Y gnd vdd DFFPOSX1
XDFFPOSX1_935 INVX1_439/A CLKBUF1_23/Y OAI21X1_719/Y gnd vdd DFFPOSX1
XOAI21X1_1367 INVX1_386/Y NOR2X1_297/Y NAND2X1_800/Y gnd DFFPOSX1_87/D vdd OAI21X1
XDFFPOSX1_979 INVX1_186/A CLKBUF1_73/Y OAI21X1_765/Y gnd vdd DFFPOSX1
XDFFPOSX1_968 INVX1_505/A CLKBUF1_67/Y OAI21X1_743/Y gnd vdd DFFPOSX1
XFILL_24_5_1 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XFILL_7_6_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_15_5_1 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XDFFPOSX1_209 MUX2X1_30/B CLKBUF1_76/Y DFFPOSX1_209/D gnd vdd DFFPOSX1
XBUFX4_230 BUFX4_28/Y gnd BUFX4_230/Y vdd BUFX4
XBUFX4_241 BUFX4_30/Y gnd BUFX4_241/Y vdd BUFX4
XBUFX4_263 BUFX4_28/Y gnd BUFX4_263/Y vdd BUFX4
XBUFX4_252 BUFX4_25/Y gnd BUFX4_252/Y vdd BUFX4
XNOR2X1_301 NOR2X1_301/A NOR2X1_303/B gnd NOR2X1_301/Y vdd NOR2X1
XBUFX4_274 BUFX4_24/Y gnd BUFX4_274/Y vdd BUFX4
XBUFX4_285 INVX8_8/Y gnd BUFX4_285/Y vdd BUFX4
XNOR2X1_334 NOR2X1_334/A NOR2X1_338/B gnd NOR2X1_334/Y vdd NOR2X1
XNOR2X1_323 NOR2X1_323/A NOR2X1_325/B gnd NOR2X1_323/Y vdd NOR2X1
XBUFX4_296 BUFX4_294/A gnd NOR2X1_91/A vdd BUFX4
XNOR2X1_312 NOR2X1_312/A NOR2X1_315/B gnd NOR2X1_312/Y vdd NOR2X1
XNOR2X1_345 NOR2X1_345/A NOR2X1_342/B gnd NOR2X1_345/Y vdd NOR2X1
XNOR2X1_356 NOR2X1_356/A NOR2X1_352/B gnd NOR2X1_356/Y vdd NOR2X1
XFILL_32_1 gnd vdd FILL
XNOR2X1_367 NOR2X1_367/A NOR2X1_367/B gnd NOR2X1_367/Y vdd NOR2X1
XNOR2X1_378 OAI21X1_1/B NOR2X1_61/B gnd NOR2X1_378/Y vdd NOR2X1
XOAI21X1_807 INVX1_22/Y BUFX4_208/Y NAND2X1_218/Y gnd OAI21X1_807/Y vdd OAI21X1
XOAI21X1_818 INVX1_33/Y BUFX4_226/Y OAI21X1_818/C gnd NAND2X1_232/B vdd OAI21X1
XOAI21X1_829 INVX1_42/Y BUFX4_244/Y OAI21X1_829/C gnd NAND2X1_250/B vdd OAI21X1
XOAI21X1_1120 INVX1_332/Y BUFX4_230/Y NAND2X1_563/Y gnd MUX2X1_245/A vdd OAI21X1
XOAI21X1_1131 INVX1_343/Y BUFX4_252/Y NAND2X1_575/Y gnd MUX2X1_254/B vdd OAI21X1
XOAI21X1_1142 INVX1_354/Y BUFX4_274/Y NAND2X1_587/Y gnd MUX2X1_262/A vdd OAI21X1
XOAI21X1_1164 INVX1_376/Y BUFX4_219/Y NAND2X1_610/Y gnd MUX2X1_278/A vdd OAI21X1
XMUX2X1_329 MUX2X1_329/A MUX2X1_329/B BUFX4_54/Y gnd MUX2X1_329/Y vdd MUX2X1
XMUX2X1_318 MUX2X1_318/A MUX2X1_318/B BUFX4_362/Y gnd AOI22X1_66/D vdd MUX2X1
XOAI21X1_1153 INVX1_365/Y BUFX4_197/Y NAND2X1_599/Y gnd MUX2X1_271/B vdd OAI21X1
XDFFPOSX1_732 NOR2X1_86/A CLKBUF1_29/Y AOI21X1_68/Y gnd vdd DFFPOSX1
XMUX2X1_307 MUX2X1_307/A MUX2X1_307/B BUFX4_53/Y gnd MUX2X1_309/B vdd MUX2X1
XDFFPOSX1_721 INVX1_58/A CLKBUF1_49/Y OAI21X1_545/Y gnd vdd DFFPOSX1
XDFFPOSX1_710 INVX1_361/A CLKBUF1_54/Y OAI21X1_524/Y gnd vdd DFFPOSX1
XOAI21X1_1197 INVX1_409/Y MUX2X1_11/S NAND2X1_646/Y gnd MUX2X1_304/B vdd OAI21X1
XDFFPOSX1_765 NOR2X1_107/A CLKBUF1_94/Y AOI21X1_85/Y gnd vdd DFFPOSX1
XDFFPOSX1_743 INVX1_427/A CLKBUF1_4/Y OAI21X1_559/Y gnd vdd DFFPOSX1
XOAI21X1_1175 INVX1_387/Y BUFX4_241/Y NAND2X1_623/Y gnd MUX2X1_287/B vdd OAI21X1
XOAI21X1_1186 INVX1_398/Y BUFX4_263/Y NAND2X1_635/Y gnd MUX2X1_295/A vdd OAI21X1
XDFFPOSX1_754 INVX1_108/A CLKBUF1_57/Y OAI21X1_562/Y gnd vdd DFFPOSX1
XNAND2X1_813 AOI22X1_9/A BUFX4_321/Y gnd BUFX4_392/A vdd NAND2X1
XDFFPOSX1_798 NOR2X1_119/A CLKBUF1_62/Y AOI21X1_95/Y gnd vdd DFFPOSX1
XDFFPOSX1_787 INVX1_174/A CLKBUF1_62/Y OAI21X1_602/Y gnd vdd DFFPOSX1
XNAND2X1_802 BUFX4_162/Y NOR2X1_309/Y gnd NAND2X1_802/Y vdd NAND2X1
XDFFPOSX1_776 INVX1_493/A CLKBUF1_92/Y OAI21X1_584/Y gnd vdd DFFPOSX1
XNAND2X1_835 INVX8_11/A INVX2_9/Y gnd NAND2X1_835/Y vdd NAND2X1
XNAND2X1_824 BUFX4_164/Y NOR2X1_331/Y gnd NAND2X1_824/Y vdd NAND2X1
XNAND2X1_846 NAND2X1_8/A NOR2X1_358/Y gnd NAND2X1_846/Y vdd NAND2X1
XNAND2X1_868 INVX8_7/A NOR2X1_378/Y gnd NAND2X1_868/Y vdd NAND2X1
XNAND2X1_857 BUFX4_327/Y NOR2X1_368/Y gnd NAND2X1_857/Y vdd NAND2X1
XFILL_47_4_1 gnd vdd FILL
XNOR2X1_30 NOR2X1_30/A NOR2X1_27/B gnd NOR2X1_30/Y vdd NOR2X1
XNOR2X1_63 NOR2X1_63/A NOR2X1_67/B gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_52 BUFX4_432/Y NOR2X1_52/B gnd NOR2X1_55/B vdd NOR2X1
XNOR2X1_41 BUFX4_432/Y NOR2X1_41/B gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_74 NOR2X1_74/A NOR2X1_77/B gnd NOR2X1_74/Y vdd NOR2X1
XNOR2X1_85 NOR2X1_85/A NOR2X1_90/B gnd NOR2X1_85/Y vdd NOR2X1
XNOR2X1_96 NOR2X1_96/A NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XFILL_30_3_1 gnd vdd FILL
XNAND2X1_109 BUFX4_162/Y NOR2X1_91/Y gnd OAI21X1_553/C vdd NAND2X1
XNAND2X1_7 BUFX4_449/Y NOR2X1_1/Y gnd NAND2X1_7/Y vdd NAND2X1
XFILL_38_4_1 gnd vdd FILL
XMUX2X1_70 MUX2X1_70/A MUX2X1_70/B BUFX4_43/Y gnd MUX2X1_70/Y vdd MUX2X1
XNOR2X1_142 NOR2X1_142/A NOR2X1_139/B gnd NOR2X1_142/Y vdd NOR2X1
XNOR2X1_131 NOR2X1_131/A NOR2X1_126/B gnd NOR2X1_131/Y vdd NOR2X1
XMUX2X1_81 MUX2X1_80/Y MUX2X1_81/B MUX2X1_48/S gnd MUX2X1_81/Y vdd MUX2X1
XNOR2X1_120 NOR2X1_120/A NOR2X1_118/B gnd AOI21X1_96/C vdd NOR2X1
XNOR2X1_153 NOR2X1_153/A NOR2X1_153/B gnd NOR2X1_153/Y vdd NOR2X1
XNOR2X1_164 NOR2X1_164/A NOR2X1_158/B gnd NOR2X1_164/Y vdd NOR2X1
XMUX2X1_92 MUX2X1_92/A MUX2X1_92/B MUX2X1_3/S gnd MUX2X1_93/A vdd MUX2X1
XNOR2X1_175 NOR2X1_175/A NOR2X1_173/B gnd NOR2X1_175/Y vdd NOR2X1
XNOR2X1_186 NOR2X1_186/A NOR2X1_186/B gnd NOR2X1_186/Y vdd NOR2X1
XNOR2X1_197 NOR2X1_197/A NOR2X1_197/B gnd NOR2X1_197/Y vdd NOR2X1
XOAI21X1_615 INVX1_112/Y NOR2X1_133/Y OAI21X1_615/C gnd OAI21X1_615/Y vdd OAI21X1
XFILL_21_3_1 gnd vdd FILL
XOAI21X1_604 INVX1_302/Y NOR2X1_111/Y OAI21X1_604/C gnd OAI21X1_604/Y vdd OAI21X1
XOAI21X1_637 BUFX4_372/Y OAI21X1_635/B OAI21X1_637/C gnd OAI21X1_637/Y vdd OAI21X1
XOAI21X1_626 BUFX4_456/Y INVX1_4/A INVX1_177/A gnd OAI21X1_626/Y vdd OAI21X1
XOAI21X1_648 BUFX4_153/Y INVX1_4/A NAND2X1_603/B gnd OAI21X1_648/Y vdd OAI21X1
XOAI21X1_659 INVX1_434/Y NOR2X1_145/B NAND2X1_157/Y gnd OAI21X1_659/Y vdd OAI21X1
XMUX2X1_104 MUX2X1_104/A MUX2X1_104/B BUFX4_52/Y gnd MUX2X1_105/A vdd MUX2X1
XDFFPOSX1_540 NOR2X1_46/A CLKBUF1_95/Y AOI21X1_36/Y gnd vdd DFFPOSX1
XMUX2X1_137 MUX2X1_137/A MUX2X1_137/B BUFX4_42/Y gnd MUX2X1_137/Y vdd MUX2X1
XMUX2X1_126 MUX2X1_126/A MUX2X1_124/Y BUFX4_364/Y gnd AOI22X1_26/D vdd MUX2X1
XMUX2X1_115 MUX2X1_115/A MUX2X1_115/B BUFX4_41/Y gnd MUX2X1_117/B vdd MUX2X1
XDFFPOSX1_562 INVX1_96/A CLKBUF1_80/Y OAI21X1_276/Y gnd vdd DFFPOSX1
XDFFPOSX1_573 NAND2X1_516/B CLKBUF1_19/Y OAI21X1_298/Y gnd vdd DFFPOSX1
XMUX2X1_148 MUX2X1_148/A MUX2X1_148/B BUFX4_34/Y gnd MUX2X1_150/B vdd MUX2X1
XMUX2X1_159 MUX2X1_159/A MUX2X1_157/Y BUFX4_364/Y gnd AOI22X1_33/A vdd MUX2X1
XDFFPOSX1_551 INVX1_415/A CLKBUF1_27/Y OAI21X1_271/Y gnd vdd DFFPOSX1
XNAND2X1_610 BUFX4_218/Y NOR2X1_207/A gnd NAND2X1_610/Y vdd NAND2X1
XDFFPOSX1_595 INVX1_162/A CLKBUF1_28/Y OAI21X1_318/Y gnd vdd DFFPOSX1
XDFFPOSX1_584 INVX1_481/A CLKBUF1_83/Y OAI21X1_312/Y gnd vdd DFFPOSX1
XNAND2X1_621 BUFX4_236/Y NAND2X1_621/B gnd NAND2X1_621/Y vdd NAND2X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XNAND2X1_632 BUFX4_258/Y NAND2X1_632/B gnd NAND2X1_632/Y vdd NAND2X1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XNAND2X1_643 BUFX4_278/Y NAND2X1_643/B gnd NAND2X1_643/Y vdd NAND2X1
XNAND2X1_654 BUFX4_199/Y NAND2X1_654/B gnd NAND2X1_654/Y vdd NAND2X1
XNAND2X1_687 BUFX4_259/Y NOR2X1_273/A gnd NAND2X1_687/Y vdd NAND2X1
XNAND2X1_676 BUFX4_241/Y NAND2X1_676/B gnd NAND2X1_676/Y vdd NAND2X1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XNAND2X1_665 BUFX4_221/Y NOR2X1_99/A gnd NAND2X1_665/Y vdd NAND2X1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XFILL_4_4_1 gnd vdd FILL
XNAND2X1_698 MUX2X1_4/S NAND2X1_698/B gnd NAND2X1_698/Y vdd NAND2X1
XFILL_29_4_1 gnd vdd FILL
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XDFFPOSX1_7 INVX1_382/A CLKBUF1_14/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XFILL_12_3_1 gnd vdd FILL
XOAI21X1_423 BUFX4_403/Y BUFX4_342/Y INVX1_230/A gnd OAI21X1_424/C vdd OAI21X1
XOAI21X1_401 NOR2X1_32/B NOR2X1_61/A NAND2X1_520/B gnd OAI21X1_402/C vdd OAI21X1
XOAI21X1_412 INVX1_229/Y NOR2X1_71/Y NAND2X1_87/Y gnd OAI21X1_412/Y vdd OAI21X1
XOAI21X1_434 BUFX4_124/Y NAND2X1_93/Y OAI21X1_434/C gnd OAI21X1_434/Y vdd OAI21X1
XOAI21X1_456 BUFX4_302/Y NAND2X1_94/Y OAI21X1_456/C gnd OAI21X1_456/Y vdd OAI21X1
XOAI21X1_445 BUFX4_88/Y NOR2X1_72/A OAI21X1_445/C gnd OAI21X1_446/C vdd OAI21X1
XOAI21X1_489 BUFX4_169/Y INVX2_4/A INVX1_296/A gnd OAI21X1_489/Y vdd OAI21X1
XOAI21X1_467 BUFX4_370/Y BUFX4_336/Y NAND2X1_316/B gnd OAI21X1_468/C vdd OAI21X1
XOAI21X1_478 BUFX4_284/Y NAND2X1_95/Y OAI21X1_478/C gnd OAI21X1_478/Y vdd OAI21X1
XINVX1_509 INVX1_509/A gnd INVX1_509/Y vdd INVX1
XDFFPOSX1_381 OAI21X1_57/C CLKBUF1_28/Y OAI21X1_58/Y gnd vdd DFFPOSX1
XDFFPOSX1_370 INVX1_84/A CLKBUF1_64/Y OAI21X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_392 INVX1_469/A CLKBUF1_69/Y OAI21X1_72/Y gnd vdd DFFPOSX1
XNAND2X1_451 BUFX4_219/Y NAND2X1_451/B gnd NAND2X1_451/Y vdd NAND2X1
XNAND2X1_440 BUFX4_199/Y NOR2X1_16/A gnd NAND2X1_440/Y vdd NAND2X1
XNAND2X1_462 BUFX4_239/Y NOR2X1_117/A gnd NAND2X1_462/Y vdd NAND2X1
XNAND2X1_484 MUX2X1_1/S NOR2X1_304/A gnd NAND2X1_484/Y vdd NAND2X1
XNAND2X1_473 BUFX4_261/Y NAND2X1_473/B gnd NAND2X1_473/Y vdd NAND2X1
XNAND2X1_495 AOI22X1_40/Y AOI22X1_41/Y gnd AOI22X1_44/A vdd NAND2X1
XFILL_44_2_1 gnd vdd FILL
XOAI21X1_990 INVX1_202/Y BUFX4_267/Y OAI21X1_990/C gnd MUX2X1_148/A vdd OAI21X1
XFILL_35_2_1 gnd vdd FILL
XOAI21X1_50 BUFX4_123/Y NAND2X1_4/Y OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_61 BUFX4_415/Y BUFX4_317/Y OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_72 INVX1_469/Y NOR2X1_1/Y NAND2X1_13/Y gnd OAI21X1_72/Y vdd OAI21X1
XOAI21X1_94 BUFX4_110/Y OAI21X1_96/B OAI21X1_94/C gnd OAI21X1_94/Y vdd OAI21X1
XOAI21X1_83 NOR2X1_81/B INVX2_1/A INVX1_342/A gnd OAI21X1_84/C vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XFILL_26_2_1 gnd vdd FILL
XOAI21X1_231 BUFX4_461/Y BUFX4_434/Y INVX1_221/A gnd OAI21X1_231/Y vdd OAI21X1
XOAI21X1_220 INVX1_220/Y NOR2X1_31/Y NAND2X1_42/Y gnd OAI21X1_220/Y vdd OAI21X1
XOAI21X1_242 BUFX4_129/Y NAND2X1_49/Y OAI21X1_241/Y gnd OAI21X1_242/Y vdd OAI21X1
XOAI21X1_264 INVX1_478/Y NOR2X1_41/Y NAND2X1_57/Y gnd OAI21X1_264/Y vdd OAI21X1
XOAI21X1_253 BUFX4_150/Y BUFX4_432/Y NAND2X1_651/B gnd OAI21X1_253/Y vdd OAI21X1
XOAI21X1_286 NAND2X1_66/Y BUFX4_287/Y OAI21X1_285/Y gnd OAI21X1_286/Y vdd OAI21X1
XOAI21X1_275 BUFX4_165/Y BUFX4_434/Y INVX1_96/A gnd OAI21X1_275/Y vdd OAI21X1
XINVX1_306 INVX1_306/A gnd INVX1_306/Y vdd INVX1
XOAI21X1_297 BUFX4_412/Y INVX2_2/A NAND2X1_516/B gnd OAI21X1_297/Y vdd OAI21X1
XINVX1_317 INVX1_317/A gnd INVX1_317/Y vdd INVX1
XINVX1_328 INVX1_328/A gnd INVX1_328/Y vdd INVX1
XINVX1_339 INVX1_339/A gnd INVX1_339/Y vdd INVX1
XFILL_9_3_1 gnd vdd FILL
XNAND2X1_270 MUX2X1_1/S NOR2X1_103/A gnd OAI21X1_848/C vdd NAND2X1
XNAND2X1_281 BUFX4_200/Y NOR2X1_324/A gnd OAI21X1_858/C vdd NAND2X1
XNAND2X1_292 BUFX4_220/Y NAND2X1_292/B gnd OAI21X1_868/C vdd NAND2X1
XFILL_17_2_1 gnd vdd FILL
XOAI21X1_1505 BUFX4_146/Y BUFX4_89/Y MUX2X1_29/A gnd OAI21X1_1506/C vdd OAI21X1
XOAI21X1_1527 BUFX4_405/Y BUFX4_91/Y INVX1_202/A gnd OAI21X1_1528/C vdd OAI21X1
XOAI21X1_1516 BUFX4_98/Y NAND2X1_835/Y OAI21X1_1515/Y gnd DFFPOSX1_206/D vdd OAI21X1
XOAI21X1_1538 NAND2X1_837/Y BUFX4_128/Y OAI21X1_1537/Y gnd DFFPOSX1_225/D vdd OAI21X1
XOAI21X1_1549 BUFX4_312/Y BUFX4_93/Y INVX1_395/A gnd OAI21X1_1550/C vdd OAI21X1
XCLKBUF1_51 BUFX4_16/Y gnd CLKBUF1_51/Y vdd CLKBUF1
XCLKBUF1_40 BUFX4_13/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XCLKBUF1_84 BUFX4_12/Y gnd CLKBUF1_84/Y vdd CLKBUF1
XCLKBUF1_73 BUFX4_15/Y gnd CLKBUF1_73/Y vdd CLKBUF1
XCLKBUF1_62 BUFX4_9/Y gnd CLKBUF1_62/Y vdd CLKBUF1
XCLKBUF1_95 BUFX4_18/Y gnd CLKBUF1_95/Y vdd CLKBUF1
XFILL_41_0_1 gnd vdd FILL
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_136 INVX1_136/A gnd INVX1_136/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XINVX1_169 INVX1_169/A gnd INVX1_169/Y vdd INVX1
XBUFX4_401 INVX8_6/Y gnd BUFX4_401/Y vdd BUFX4
XBUFX4_412 INVX8_16/Y gnd BUFX4_412/Y vdd BUFX4
XBUFX4_434 BUFX4_436/A gnd BUFX4_434/Y vdd BUFX4
XBUFX4_456 INVX8_10/Y gnd BUFX4_456/Y vdd BUFX4
XBUFX4_423 INVX8_3/Y gnd BUFX4_423/Y vdd BUFX4
XBUFX4_445 d[4] gnd BUFX4_445/Y vdd BUFX4
XBUFX4_467 BUFX4_467/A gnd BUFX4_467/Y vdd BUFX4
XFILL_32_0_1 gnd vdd FILL
XAOI21X1_129 BUFX4_299/Y NOR2X1_158/B NOR2X1_161/Y gnd AOI21X1_129/Y vdd AOI21X1
XAOI21X1_107 BUFX4_124/Y NOR2X1_133/Y NOR2X1_134/Y gnd AOI21X1_107/Y vdd AOI21X1
XAOI21X1_118 BUFX4_418/Y NOR2X1_153/B NOR2X1_148/Y gnd AOI21X1_118/Y vdd AOI21X1
XOAI21X1_1313 INVX1_35/Y NOR2X1_274/Y NAND2X1_775/Y gnd DFFPOSX1_33/D vdd OAI21X1
XOAI21X1_1302 INVX1_317/Y NOR2X1_254/Y NAND2X1_761/Y gnd DFFPOSX1_30/D vdd OAI21X1
XOAI21X1_1346 BUFX4_125/Y NAND2X1_793/Y OAI21X1_1345/Y gnd DFFPOSX1_73/D vdd OAI21X1
XOAI21X1_1335 BUFX4_454/Y BUFX4_468/Y INVX1_193/A gnd OAI21X1_1335/Y vdd OAI21X1
XDFFPOSX1_914 INVX1_118/A CLKBUF1_76/Y OAI21X1_707/Y gnd vdd DFFPOSX1
XDFFPOSX1_903 INVX1_437/A CLKBUF1_101/Y OAI21X1_688/Y gnd vdd DFFPOSX1
XOAI21X1_1324 INVX1_192/Y NOR2X1_284/Y NAND2X1_786/Y gnd DFFPOSX1_52/D vdd OAI21X1
XOAI21X1_1379 BUFX4_168/Y BUFX4_468/Y INVX1_68/A gnd OAI21X1_1380/C vdd OAI21X1
XDFFPOSX1_936 INVX1_503/A CLKBUF1_90/Y OAI21X1_720/Y gnd vdd DFFPOSX1
XDFFPOSX1_925 NOR2X1_184/A CLKBUF1_9/Y AOI21X1_148/Y gnd vdd DFFPOSX1
XDFFPOSX1_947 INVX1_184/A CLKBUF1_14/Y OAI21X1_722/Y gnd vdd DFFPOSX1
XOAI21X1_1357 BUFX4_154/Y BUFX4_463/Y NAND2X1_621/B gnd OAI21X1_1357/Y vdd OAI21X1
XOAI21X1_1368 INVX1_450/Y NOR2X1_297/Y NAND2X1_801/Y gnd DFFPOSX1_88/D vdd OAI21X1
XDFFPOSX1_958 NOR2X1_207/A CLKBUF1_90/Y AOI21X1_167/Y gnd vdd DFFPOSX1
XDFFPOSX1_969 MUX2X1_22/A CLKBUF1_67/Y OAI21X1_745/Y gnd vdd DFFPOSX1
XFILL_23_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XFILL_43_8_0 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XBUFX4_220 BUFX4_31/Y gnd BUFX4_220/Y vdd BUFX4
XBUFX4_264 BUFX4_31/Y gnd BUFX4_264/Y vdd BUFX4
XBUFX4_231 BUFX4_31/Y gnd BUFX4_231/Y vdd BUFX4
XBUFX4_253 BUFX4_23/Y gnd BUFX4_253/Y vdd BUFX4
XBUFX4_242 BUFX4_27/Y gnd BUFX4_242/Y vdd BUFX4
XNOR2X1_302 NOR2X1_302/A NOR2X1_303/B gnd NOR2X1_302/Y vdd NOR2X1
XBUFX4_275 BUFX4_30/Y gnd BUFX4_275/Y vdd BUFX4
XNOR2X1_324 NOR2X1_324/A NOR2X1_325/B gnd NOR2X1_324/Y vdd NOR2X1
XBUFX4_297 INVX8_5/Y gnd BUFX4_297/Y vdd BUFX4
XNOR2X1_313 NOR2X1_313/A NOR2X1_315/B gnd NOR2X1_313/Y vdd NOR2X1
XBUFX4_286 INVX8_8/Y gnd BUFX4_286/Y vdd BUFX4
XNOR2X1_346 NOR2X1_346/A NOR2X1_342/B gnd NOR2X1_346/Y vdd NOR2X1
XNOR2X1_357 NOR2X1_357/A NOR2X1_352/B gnd NOR2X1_357/Y vdd NOR2X1
XNOR2X1_335 NOR2X1_335/A NOR2X1_338/B gnd NOR2X1_335/Y vdd NOR2X1
XFILL_34_8_0 gnd vdd FILL
XNOR2X1_368 INVX2_10/A NOR2X1_51/B gnd NOR2X1_368/Y vdd NOR2X1
XNOR2X1_379 INVX2_11/A NOR2X1_72/B gnd NOR2X1_387/B vdd NOR2X1
XFILL_25_1 gnd vdd FILL
XOAI21X1_808 INVX1_23/Y BUFX4_210/Y NAND2X1_220/Y gnd AOI22X1_2/A vdd OAI21X1
XOAI21X1_819 INVX1_34/Y BUFX4_228/Y NAND2X1_233/Y gnd OAI21X1_819/Y vdd OAI21X1
XOAI21X1_1121 INVX1_333/Y BUFX4_232/Y NAND2X1_565/Y gnd MUX2X1_247/B vdd OAI21X1
XOAI21X1_1110 INVX1_322/Y BUFX4_210/Y NAND2X1_553/Y gnd MUX2X1_238/A vdd OAI21X1
XDFFPOSX1_700 NAND2X1_455/B CLKBUF1_38/Y OAI21X1_504/Y gnd vdd DFFPOSX1
XOAI21X1_1143 INVX1_355/Y BUFX4_276/Y NAND2X1_588/Y gnd MUX2X1_263/B vdd OAI21X1
XOAI21X1_1165 INVX1_377/Y BUFX4_221/Y NAND2X1_611/Y gnd MUX2X1_280/B vdd OAI21X1
XDFFPOSX1_722 INVX1_106/A CLKBUF1_72/Y OAI21X1_546/Y gnd vdd DFFPOSX1
XMUX2X1_319 MUX2X1_319/A MUX2X1_319/B BUFX4_58/Y gnd MUX2X1_321/B vdd MUX2X1
XOAI21X1_1154 INVX1_366/Y BUFX4_199/Y NAND2X1_600/Y gnd MUX2X1_271/A vdd OAI21X1
XMUX2X1_308 MUX2X1_308/A MUX2X1_308/B BUFX4_6/Y gnd MUX2X1_309/A vdd MUX2X1
XOAI21X1_1132 INVX1_344/Y BUFX4_254/Y NAND2X1_576/Y gnd MUX2X1_254/A vdd OAI21X1
XDFFPOSX1_711 INVX1_425/A CLKBUF1_54/Y OAI21X1_526/Y gnd vdd DFFPOSX1
XOAI21X1_1198 INVX1_410/Y BUFX4_188/Y NAND2X1_647/Y gnd MUX2X1_304/A vdd OAI21X1
XDFFPOSX1_766 NOR2X1_108/A CLKBUF1_72/Y AOI21X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_755 INVX1_172/A CLKBUF1_4/Y OAI21X1_563/Y gnd vdd DFFPOSX1
XDFFPOSX1_733 NOR2X1_87/A CLKBUF1_94/Y AOI21X1_69/Y gnd vdd DFFPOSX1
XOAI21X1_1176 INVX1_388/Y BUFX4_243/Y NAND2X1_624/Y gnd MUX2X1_287/A vdd OAI21X1
XOAI21X1_1187 INVX1_399/Y BUFX4_265/Y NAND2X1_636/Y gnd MUX2X1_296/B vdd OAI21X1
XDFFPOSX1_744 INVX1_491/A CLKBUF1_92/Y OAI21X1_560/Y gnd vdd DFFPOSX1
XDFFPOSX1_777 MUX2X1_1/A CLKBUF1_74/Y OAI21X1_586/Y gnd vdd DFFPOSX1
XNAND2X1_803 INVX8_3/A NOR2X1_309/Y gnd NAND2X1_803/Y vdd NAND2X1
XDFFPOSX1_788 INVX1_238/A CLKBUF1_62/Y OAI21X1_603/Y gnd vdd DFFPOSX1
XDFFPOSX1_799 NOR2X1_120/A CLKBUF1_92/Y AOI21X1_96/Y gnd vdd DFFPOSX1
XNAND2X1_836 INVX2_9/Y INVX8_12/A gnd NAND2X1_836/Y vdd NAND2X1
XNAND2X1_825 BUFX4_453/Y NOR2X1_331/Y gnd NAND2X1_825/Y vdd NAND2X1
XNAND2X1_814 INVX8_10/A INVX2_8/Y gnd NAND2X1_814/Y vdd NAND2X1
XNAND2X1_869 INVX8_8/A NOR2X1_378/Y gnd NAND2X1_869/Y vdd NAND2X1
XNAND2X1_847 NAND2X1_9/A NOR2X1_358/Y gnd NAND2X1_847/Y vdd NAND2X1
XNAND2X1_858 BUFX4_137/Y NOR2X1_368/Y gnd NAND2X1_858/Y vdd NAND2X1
XFILL_0_8_0 gnd vdd FILL
XFILL_25_8_0 gnd vdd FILL
XNOR2X1_20 NOR2X1_20/A NOR2X1_14/B gnd NOR2X1_20/Y vdd NOR2X1
XNOR2X1_53 NOR2X1_53/A NOR2X1_55/B gnd NOR2X1_53/Y vdd NOR2X1
XNOR2X1_64 NOR2X1_64/A NOR2X1_67/B gnd NOR2X1_64/Y vdd NOR2X1
XNOR2X1_31 BUFX4_135/Y BUFX4_166/Y gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_42 BUFX4_432/Y BUFX4_84/Y gnd NOR2X1_43/B vdd NOR2X1
XFILL_16_8_0 gnd vdd FILL
XNOR2X1_75 NOR2X1_75/A NOR2X1_77/B gnd NOR2X1_75/Y vdd NOR2X1
XNOR2X1_86 NOR2X1_86/A NOR2X1_90/B gnd NOR2X1_86/Y vdd NOR2X1
XNOR2X1_97 NOR2X1_97/A NOR2X1_96/B gnd NOR2X1_97/Y vdd NOR2X1
XNAND2X1_8 NAND2X1_8/A NOR2X1_1/Y gnd NAND2X1_8/Y vdd NAND2X1
XMUX2X1_71 MUX2X1_71/A MUX2X1_71/B BUFX4_59/Y gnd MUX2X1_71/Y vdd MUX2X1
XMUX2X1_60 MUX2X1_59/Y MUX2X1_58/Y BUFX4_364/Y gnd MUX2X1_60/Y vdd MUX2X1
XNOR2X1_132 NOR2X1_132/A NOR2X1_126/B gnd NOR2X1_132/Y vdd NOR2X1
XNOR2X1_121 NOR2X1_121/A NOR2X1_118/B gnd NOR2X1_121/Y vdd NOR2X1
XNOR2X1_110 NOR2X1_110/A NOR2X1_103/B gnd NOR2X1_110/Y vdd NOR2X1
XNOR2X1_176 NOR2X1_176/A NOR2X1_173/B gnd NOR2X1_176/Y vdd NOR2X1
XNOR2X1_154 NOR2X1_154/A NOR2X1_153/B gnd NOR2X1_154/Y vdd NOR2X1
XNOR2X1_165 NOR2X1_165/A NOR2X1_158/B gnd NOR2X1_165/Y vdd NOR2X1
XMUX2X1_93 MUX2X1_93/A MUX2X1_91/Y BUFX4_364/Y gnd MUX2X1_93/Y vdd MUX2X1
XNOR2X1_143 NOR2X1_143/A NOR2X1_139/B gnd NOR2X1_143/Y vdd NOR2X1
XMUX2X1_82 MUX2X1_82/A MUX2X1_82/B BUFX4_55/Y gnd MUX2X1_84/B vdd MUX2X1
XNOR2X1_198 NOR2X1_198/A NOR2X1_197/B gnd NOR2X1_198/Y vdd NOR2X1
XNOR2X1_187 NOR2X1_187/A NOR2X1_186/B gnd NOR2X1_187/Y vdd NOR2X1
XOAI21X1_605 INVX1_366/Y NOR2X1_111/Y NAND2X1_132/Y gnd OAI21X1_605/Y vdd OAI21X1
XOAI21X1_638 BUFX4_153/Y BUFX4_121/Y MUX2X1_8/A gnd OAI21X1_639/C vdd OAI21X1
XOAI21X1_627 BUFX4_116/Y OAI21X1_635/B OAI21X1_626/Y gnd OAI21X1_627/Y vdd OAI21X1
XOAI21X1_616 INVX1_176/Y NOR2X1_133/Y OAI21X1_616/C gnd OAI21X1_616/Y vdd OAI21X1
XOAI21X1_649 BUFX4_104/Y OAI21X1_651/B OAI21X1_648/Y gnd OAI21X1_649/Y vdd OAI21X1
XMUX2X1_105 MUX2X1_105/A MUX2X1_103/Y BUFX4_357/Y gnd AOI22X1_22/A vdd MUX2X1
XDFFPOSX1_541 NOR2X1_47/A CLKBUF1_91/Y AOI21X1_37/Y gnd vdd DFFPOSX1
XMUX2X1_138 MUX2X1_137/Y MUX2X1_136/Y BUFX4_357/Y gnd MUX2X1_138/Y vdd MUX2X1
XMUX2X1_127 MUX2X1_127/A MUX2X1_127/B BUFX4_53/Y gnd MUX2X1_129/B vdd MUX2X1
XMUX2X1_116 MUX2X1_116/A MUX2X1_116/B BUFX4_57/Y gnd MUX2X1_117/A vdd MUX2X1
XDFFPOSX1_530 INVX1_94/A CLKBUF1_57/Y OAI21X1_258/Y gnd vdd DFFPOSX1
XDFFPOSX1_552 INVX1_479/A CLKBUF1_95/Y OAI21X1_272/Y gnd vdd DFFPOSX1
XMUX2X1_149 MUX2X1_149/A MUX2X1_149/B BUFX4_54/Y gnd MUX2X1_149/Y vdd MUX2X1
XDFFPOSX1_574 NAND2X1_585/B CLKBUF1_41/Y OAI21X1_300/Y gnd vdd DFFPOSX1
XDFFPOSX1_563 INVX1_160/A CLKBUF1_19/Y OAI21X1_278/Y gnd vdd DFFPOSX1
XDFFPOSX1_585 NOR2X1_63/A CLKBUF1_22/Y AOI21X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_596 INVX1_226/A CLKBUF1_79/Y OAI21X1_320/Y gnd vdd DFFPOSX1
XNAND2X1_611 BUFX4_220/Y NAND2X1_611/B gnd NAND2X1_611/Y vdd NAND2X1
XNAND2X1_600 INVX8_1/A NOR2X1_119/A gnd NAND2X1_600/Y vdd NAND2X1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XNAND2X1_655 BUFX4_201/Y NOR2X1_69/A gnd NAND2X1_655/Y vdd NAND2X1
XINVX1_12 a[6] gnd INVX1_12/Y vdd INVX1
XNAND2X1_633 AOI22X1_60/Y AOI22X1_61/Y gnd AOI22X1_64/A vdd NAND2X1
XNAND2X1_644 MUX2X1_2/S OAI21X1_133/C gnd NAND2X1_644/Y vdd NAND2X1
XNAND2X1_622 BUFX4_238/Y NOR2X1_306/A gnd NAND2X1_622/Y vdd NAND2X1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XNAND2X1_677 BUFX4_243/Y NOR2X1_186/A gnd NAND2X1_677/Y vdd NAND2X1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XNAND2X1_688 BUFX4_261/Y NOR2X1_283/A gnd NAND2X1_688/Y vdd NAND2X1
XNAND2X1_666 BUFX4_223/Y NOR2X1_109/A gnd NAND2X1_666/Y vdd NAND2X1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XNAND2X1_699 MUX2X1_8/S NOR2X1_349/A gnd NAND2X1_699/Y vdd NAND2X1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XDFFPOSX1_8 INVX1_446/A CLKBUF1_90/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XFILL_40_6_0 gnd vdd FILL
XAOI21X1_290 BUFX4_399/Y NOR2X1_367/B NOR2X1_364/Y gnd AOI21X1_290/Y vdd AOI21X1
XFILL_48_7_0 gnd vdd FILL
XFILL_31_6_0 gnd vdd FILL
XFILL_39_7_0 gnd vdd FILL
XFILL_22_6_0 gnd vdd FILL
XOAI21X1_402 BUFX4_398/Y NAND2X1_82/Y OAI21X1_402/C gnd OAI21X1_402/Y vdd OAI21X1
XOAI21X1_413 INVX1_293/Y NOR2X1_71/Y NAND2X1_88/Y gnd OAI21X1_413/Y vdd OAI21X1
XOAI21X1_424 BUFX4_302/Y NAND2X1_92/Y OAI21X1_424/C gnd OAI21X1_424/Y vdd OAI21X1
XOAI21X1_457 BUFX4_310/Y BUFX4_336/Y INVX1_295/A gnd OAI21X1_458/C vdd OAI21X1
XOAI21X1_435 BUFX4_88/Y BUFX4_337/Y NAND2X1_315/B gnd OAI21X1_436/C vdd OAI21X1
XOAI21X1_446 BUFX4_284/Y NAND2X1_93/Y OAI21X1_446/C gnd OAI21X1_446/Y vdd OAI21X1
XOAI21X1_479 BUFX4_370/Y INVX2_4/A NAND2X1_730/B gnd OAI21X1_479/Y vdd OAI21X1
XOAI21X1_468 BUFX4_421/Y NAND2X1_95/Y OAI21X1_468/C gnd OAI21X1_468/Y vdd OAI21X1
XDFFPOSX1_382 OAI21X1_59/C CLKBUF1_28/Y OAI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_360 INVX1_467/A CLKBUF1_8/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_371 INVX1_148/A CLKBUF1_16/Y OAI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_393 NOR2X1_3/A CLKBUF1_93/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XNAND2X1_452 BUFX4_221/Y NOR2X1_76/A gnd NAND2X1_452/Y vdd NAND2X1
XNAND2X1_441 BUFX4_201/Y NOR2X1_26/A gnd NAND2X1_441/Y vdd NAND2X1
XNAND2X1_463 BUFX4_241/Y NOR2X1_128/A gnd NAND2X1_463/Y vdd NAND2X1
XNAND2X1_430 BUFX4_278/Y NAND2X1_430/B gnd OAI21X1_996/C vdd NAND2X1
XFILL_5_7_0 gnd vdd FILL
XNAND2X1_474 BUFX4_263/Y NOR2X1_214/A gnd NAND2X1_474/Y vdd NAND2X1
XNAND2X1_496 BUFX4_202/Y NAND2X1_496/B gnd NAND2X1_496/Y vdd NAND2X1
XNAND2X1_485 MUX2X1_4/S NOR2X1_316/A gnd NAND2X1_485/Y vdd NAND2X1
XFILL_13_6_0 gnd vdd FILL
XOAI21X1_991 INVX1_203/Y BUFX4_269/Y OAI21X1_991/C gnd MUX2X1_149/B vdd OAI21X1
XOAI21X1_980 INVX1_192/Y BUFX4_247/Y OAI21X1_980/C gnd MUX2X1_140/A vdd OAI21X1
XOAI21X1_51 BUFX4_415/Y BUFX4_317/Y OAI21X1_51/C gnd OAI21X1_52/C vdd OAI21X1
XOAI21X1_62 BUFX4_283/Y NAND2X1_4/Y OAI21X1_61/Y gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_40 NAND2X1_3/Y BUFX4_300/Y OAI21X1_40/C gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_73 NOR2X1_41/B NOR2X1_2/A INVX1_27/A gnd OAI21X1_74/C vdd OAI21X1
XOAI21X1_84 BUFX4_103/Y OAI21X1_82/B OAI21X1_84/C gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_95 BUFX4_86/Y NOR2X1_1/A OAI21X1_95/C gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_210 INVX1_91/Y NOR2X1_21/Y NAND2X1_32/Y gnd OAI21X1_210/Y vdd OAI21X1
XOAI21X1_221 INVX1_284/Y NOR2X1_31/Y NAND2X1_43/Y gnd OAI21X1_221/Y vdd OAI21X1
XOAI21X1_232 BUFX4_299/Y NAND2X1_48/Y OAI21X1_231/Y gnd OAI21X1_232/Y vdd OAI21X1
XOAI21X1_243 BUFX4_150/Y INVX2_2/A NAND2X1_306/B gnd OAI21X1_243/Y vdd OAI21X1
XOAI21X1_254 BUFX4_287/Y NAND2X1_49/Y OAI21X1_253/Y gnd OAI21X1_254/Y vdd OAI21X1
XOAI21X1_265 INVX1_47/Y NOR2X1_51/Y NAND2X1_58/Y gnd OAI21X1_265/Y vdd OAI21X1
XOAI21X1_276 NAND2X1_66/Y BUFX4_422/Y OAI21X1_275/Y gnd OAI21X1_276/Y vdd OAI21X1
XINVX1_307 INVX1_307/A gnd INVX1_307/Y vdd INVX1
XOAI21X1_298 BUFX4_394/Y NAND2X1_67/Y OAI21X1_297/Y gnd OAI21X1_298/Y vdd OAI21X1
XOAI21X1_287 BUFX4_165/Y BUFX4_434/Y INVX1_480/A gnd OAI21X1_288/C vdd OAI21X1
XINVX1_318 INVX1_318/A gnd INVX1_318/Y vdd INVX1
XINVX1_329 INVX1_329/A gnd INVX1_329/Y vdd INVX1
XDFFPOSX1_190 NAND2X1_559/B CLKBUF1_78/Y OAI21X1_1484/Y gnd vdd DFFPOSX1
XNAND2X1_260 BUFX4_259/Y NAND2X1_260/B gnd NAND2X1_260/Y vdd NAND2X1
XNAND2X1_271 AOI22X1_7/Y AOI22X1_8/Y gnd AOI22X1_9/C vdd NAND2X1
XNAND2X1_293 BUFX4_222/Y NOR2X1_381/A gnd OAI21X1_869/C vdd NAND2X1
XNAND2X1_282 BUFX4_202/Y NOR2X1_334/A gnd OAI21X1_859/C vdd NAND2X1
XFILL_45_5_0 gnd vdd FILL
XOAI21X1_1517 BUFX4_147/Y BUFX4_92/Y NAND2X1_629/B gnd OAI21X1_1518/C vdd OAI21X1
XOAI21X1_1539 NOR2X1_21/B INVX2_9/A INVX1_75/A gnd OAI21X1_1540/C vdd OAI21X1
XOAI21X1_1528 NAND2X1_836/Y BUFX4_303/Y OAI21X1_1528/C gnd OAI21X1_1528/Y vdd OAI21X1
XOAI21X1_1506 BUFX4_128/Y NAND2X1_835/Y OAI21X1_1506/C gnd OAI21X1_1506/Y vdd OAI21X1
XFILL_36_5_0 gnd vdd FILL
XCLKBUF1_41 BUFX4_18/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XCLKBUF1_30 BUFX4_13/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XCLKBUF1_52 BUFX4_17/Y gnd CLKBUF1_52/Y vdd CLKBUF1
XCLKBUF1_63 BUFX4_11/Y gnd CLKBUF1_63/Y vdd CLKBUF1
XCLKBUF1_74 BUFX4_9/Y gnd CLKBUF1_74/Y vdd CLKBUF1
XCLKBUF1_96 BUFX4_10/Y gnd CLKBUF1_96/Y vdd CLKBUF1
XCLKBUF1_85 BUFX4_15/Y gnd CLKBUF1_85/Y vdd CLKBUF1
XFILL_2_5_0 gnd vdd FILL
XFILL_27_5_0 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XINVX1_115 INVX1_115/A gnd INVX1_115/Y vdd INVX1
XINVX1_159 INVX1_159/A gnd INVX1_159/Y vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd INVX1_137/Y vdd INVX1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XBUFX4_402 INVX8_6/Y gnd BUFX4_402/Y vdd BUFX4
XBUFX4_413 INVX8_16/Y gnd NOR2X1_32/B vdd BUFX4
XBUFX4_435 BUFX4_436/A gnd INVX2_2/A vdd BUFX4
XBUFX4_424 INVX8_3/Y gnd BUFX4_424/Y vdd BUFX4
XBUFX4_446 d[4] gnd INVX8_6/A vdd BUFX4
XBUFX4_468 BUFX4_467/A gnd BUFX4_468/Y vdd BUFX4
XFILL_18_5_0 gnd vdd FILL
XBUFX4_457 INVX8_10/Y gnd BUFX4_457/Y vdd BUFX4
XAOI21X1_119 BUFX4_116/Y NOR2X1_153/B NOR2X1_149/Y gnd AOI21X1_119/Y vdd AOI21X1
XAOI21X1_108 BUFX4_124/Y NOR2X1_139/B NOR2X1_136/Y gnd AOI21X1_108/Y vdd AOI21X1
XOAI21X1_1303 INVX1_381/Y NOR2X1_254/Y NAND2X1_762/Y gnd DFFPOSX1_31/D vdd OAI21X1
XOAI21X1_1314 INVX1_63/Y NOR2X1_274/Y NAND2X1_776/Y gnd DFFPOSX1_34/D vdd OAI21X1
XOAI21X1_1336 BUFX4_305/Y NAND2X1_792/Y OAI21X1_1335/Y gnd DFFPOSX1_68/D vdd OAI21X1
XDFFPOSX1_915 INVX1_182/A CLKBUF1_21/Y OAI21X1_708/Y gnd vdd DFFPOSX1
XDFFPOSX1_904 INVX1_501/A CLKBUF1_101/Y OAI21X1_690/Y gnd vdd DFFPOSX1
XOAI21X1_1325 INVX1_256/Y NOR2X1_284/Y NAND2X1_787/Y gnd DFFPOSX1_53/D vdd OAI21X1
XOAI21X1_1347 BUFX4_151/Y BUFX4_463/Y NAND2X1_276/B gnd OAI21X1_1347/Y vdd OAI21X1
XDFFPOSX1_926 NOR2X1_185/A CLKBUF1_51/Y AOI21X1_149/Y gnd vdd DFFPOSX1
XDFFPOSX1_937 MUX2X1_18/A CLKBUF1_101/Y AOI21X1_153/Y gnd vdd DFFPOSX1
XDFFPOSX1_948 INVX1_248/A CLKBUF1_87/Y OAI21X1_723/Y gnd vdd DFFPOSX1
XOAI21X1_1369 INVX1_39/Y NOR2X1_309/Y NAND2X1_802/Y gnd DFFPOSX1_97/D vdd OAI21X1
XOAI21X1_1358 BUFX4_286/Y NAND2X1_793/Y OAI21X1_1357/Y gnd DFFPOSX1_79/D vdd OAI21X1
XDFFPOSX1_959 NOR2X1_208/A CLKBUF1_9/Y AOI21X1_168/Y gnd vdd DFFPOSX1
XFILL_43_8_1 gnd vdd FILL
XFILL_42_3_0 gnd vdd FILL
XBUFX4_210 BUFX4_26/Y gnd BUFX4_210/Y vdd BUFX4
XBUFX4_221 BUFX4_27/Y gnd BUFX4_221/Y vdd BUFX4
XBUFX4_254 BUFX4_24/Y gnd BUFX4_254/Y vdd BUFX4
XBUFX4_232 BUFX4_28/Y gnd BUFX4_232/Y vdd BUFX4
XBUFX4_243 BUFX4_27/Y gnd BUFX4_243/Y vdd BUFX4
XNOR2X1_303 NOR2X1_303/A NOR2X1_303/B gnd NOR2X1_303/Y vdd NOR2X1
XBUFX4_265 BUFX4_31/Y gnd BUFX4_265/Y vdd BUFX4
XBUFX4_276 BUFX4_28/Y gnd BUFX4_276/Y vdd BUFX4
XBUFX4_298 INVX8_5/Y gnd BUFX4_298/Y vdd BUFX4
XNOR2X1_325 NOR2X1_325/A NOR2X1_325/B gnd NOR2X1_325/Y vdd NOR2X1
XNOR2X1_314 NOR2X1_314/A NOR2X1_315/B gnd NOR2X1_314/Y vdd NOR2X1
XBUFX4_287 INVX8_8/Y gnd BUFX4_287/Y vdd BUFX4
XNOR2X1_347 NOR2X1_347/A NOR2X1_342/B gnd NOR2X1_347/Y vdd NOR2X1
XNOR2X1_336 NOR2X1_336/A NOR2X1_338/B gnd NOR2X1_336/Y vdd NOR2X1
XNOR2X1_358 BUFX4_348/Y NOR2X1_41/B gnd NOR2X1_358/Y vdd NOR2X1
XFILL_34_8_1 gnd vdd FILL
XFILL_33_3_0 gnd vdd FILL
XNOR2X1_369 INVX2_10/A BUFX4_371/Y gnd NOR2X1_373/B vdd NOR2X1
XOAI21X1_809 INVX1_24/Y BUFX4_212/Y NAND2X1_221/Y gnd AOI22X1_2/D vdd OAI21X1
XOAI21X1_1100 INVX1_312/Y BUFX4_190/Y NAND2X1_541/Y gnd MUX2X1_230/A vdd OAI21X1
XOAI21X1_1111 INVX1_323/Y BUFX4_212/Y NAND2X1_554/Y gnd MUX2X1_239/B vdd OAI21X1
XOAI21X1_1122 INVX1_334/Y BUFX4_234/Y NAND2X1_566/Y gnd MUX2X1_247/A vdd OAI21X1
XDFFPOSX1_712 INVX1_489/A CLKBUF1_7/Y OAI21X1_528/Y gnd vdd DFFPOSX1
XDFFPOSX1_701 NAND2X1_524/B CLKBUF1_70/Y OAI21X1_506/Y gnd vdd DFFPOSX1
XOAI21X1_1133 INVX1_345/Y BUFX4_256/Y NAND2X1_577/Y gnd MUX2X1_256/B vdd OAI21X1
XOAI21X1_1144 INVX1_356/Y BUFX4_278/Y NAND2X1_589/Y gnd MUX2X1_263/A vdd OAI21X1
XOAI21X1_1155 INVX1_367/Y BUFX4_201/Y NAND2X1_601/Y gnd MUX2X1_272/B vdd OAI21X1
XDFFPOSX1_723 INVX1_170/A CLKBUF1_30/Y OAI21X1_547/Y gnd vdd DFFPOSX1
XMUX2X1_309 MUX2X1_309/A MUX2X1_309/B INVX2_6/A gnd AOI22X1_65/A vdd MUX2X1
XOAI21X1_1166 INVX1_378/Y BUFX4_223/Y NAND2X1_612/Y gnd MUX2X1_280/A vdd OAI21X1
XDFFPOSX1_734 NOR2X1_88/A CLKBUF1_29/Y AOI21X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_756 INVX1_236/A CLKBUF1_29/Y OAI21X1_564/Y gnd vdd DFFPOSX1
XDFFPOSX1_745 NOR2X1_93/A CLKBUF1_39/Y AOI21X1_73/Y gnd vdd DFFPOSX1
XOAI21X1_1177 INVX1_389/Y BUFX4_245/Y NAND2X1_625/Y gnd MUX2X1_289/B vdd OAI21X1
XOAI21X1_1188 INVX1_400/Y BUFX4_267/Y NAND2X1_637/Y gnd MUX2X1_296/A vdd OAI21X1
XOAI21X1_1199 INVX1_411/Y BUFX4_190/Y NAND2X1_648/Y gnd MUX2X1_305/B vdd OAI21X1
XDFFPOSX1_767 NOR2X1_109/A CLKBUF1_49/Y AOI21X1_87/Y gnd vdd DFFPOSX1
XNAND2X1_804 INVX8_4/A NOR2X1_309/Y gnd NAND2X1_804/Y vdd NAND2X1
XDFFPOSX1_778 OAI21X1_587/C CLKBUF1_74/Y OAI21X1_588/Y gnd vdd DFFPOSX1
XDFFPOSX1_789 INVX1_302/A CLKBUF1_92/Y OAI21X1_604/Y gnd vdd DFFPOSX1
XNAND2X1_837 INVX2_9/Y INVX8_14/A gnd NAND2X1_837/Y vdd NAND2X1
XNAND2X1_826 BUFX4_335/Y NOR2X1_331/Y gnd NAND2X1_826/Y vdd NAND2X1
XINVX1_490 INVX1_490/A gnd INVX1_490/Y vdd INVX1
XNAND2X1_815 INVX8_11/A INVX2_8/Y gnd NAND2X1_815/Y vdd NAND2X1
XNAND2X1_848 BUFX4_444/Y NOR2X1_358/Y gnd NAND2X1_848/Y vdd NAND2X1
XNAND2X1_859 BUFX4_428/Y NOR2X1_368/Y gnd NAND2X1_859/Y vdd NAND2X1
XFILL_0_8_1 gnd vdd FILL
XFILL_25_8_1 gnd vdd FILL
XFILL_24_3_0 gnd vdd FILL
XFILL_7_4_0 gnd vdd FILL
XNOR2X1_21 BUFX4_135/Y NOR2X1_21/B gnd NOR2X1_21/Y vdd NOR2X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_2/Y gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_43 NOR2X1_43/A NOR2X1_43/B gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_54 NOR2X1_54/A NOR2X1_55/B gnd NOR2X1_54/Y vdd NOR2X1
XNOR2X1_32 BUFX4_135/Y NOR2X1_32/B gnd NOR2X1_38/B vdd NOR2X1
XNOR2X1_65 NOR2X1_65/A NOR2X1_67/B gnd NOR2X1_65/Y vdd NOR2X1
XFILL_16_8_1 gnd vdd FILL
XNOR2X1_76 NOR2X1_76/A NOR2X1_77/B gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_87 NOR2X1_87/A NOR2X1_90/B gnd NOR2X1_87/Y vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNOR2X1_98 NOR2X1_98/A NOR2X1_96/B gnd NOR2X1_98/Y vdd NOR2X1
XNAND2X1_9 NAND2X1_9/A NOR2X1_1/Y gnd NAND2X1_9/Y vdd NAND2X1
XNOR2X1_100 NOR2X1_100/A NOR2X1_96/B gnd AOI21X1_80/C vdd NOR2X1
XMUX2X1_72 MUX2X1_71/Y MUX2X1_70/Y BUFX4_357/Y gnd MUX2X1_72/Y vdd MUX2X1
XNOR2X1_133 BUFX4_105/Y BUFX4_166/Y gnd NOR2X1_133/Y vdd NOR2X1
XNOR2X1_122 BUFX4_105/Y NOR2X1_91/B gnd NOR2X1_122/Y vdd NOR2X1
XMUX2X1_50 MUX2X1_50/A MUX2X1_50/B BUFX4_21/Y gnd MUX2X1_51/A vdd MUX2X1
XMUX2X1_61 MUX2X1_61/A MUX2X1_61/B BUFX4_7/Y gnd MUX2X1_61/Y vdd MUX2X1
XNOR2X1_111 BUFX4_105/Y NOR2X1_81/B gnd NOR2X1_111/Y vdd NOR2X1
XMUX2X1_83 MUX2X1_83/A MUX2X1_83/B BUFX4_8/Y gnd MUX2X1_84/A vdd MUX2X1
XNOR2X1_155 BUFX4_118/Y NOR2X1_91/B gnd NOR2X1_155/Y vdd NOR2X1
XNOR2X1_144 BUFX4_118/Y NOR2X1_81/B gnd NOR2X1_145/B vdd NOR2X1
XNOR2X1_166 BUFX4_118/Y BUFX4_165/Y gnd NOR2X1_166/Y vdd NOR2X1
XMUX2X1_94 MUX2X1_94/A MUX2X1_94/B BUFX4_56/Y gnd MUX2X1_96/B vdd MUX2X1
XNOR2X1_188 INVX1_5/A NOR2X1_21/B gnd NOR2X1_189/B vdd NOR2X1
XNOR2X1_199 BUFX4_64/Y BUFX4_166/Y gnd NOR2X1_199/Y vdd NOR2X1
XNOR2X1_177 BUFX4_64/Y BUFX4_405/Y gnd NOR2X1_177/Y vdd NOR2X1
XOAI21X1_606 INVX1_430/Y NOR2X1_111/Y OAI21X1_606/C gnd OAI21X1_606/Y vdd OAI21X1
XOAI21X1_628 BUFX4_456/Y BUFX4_120/Y INVX1_241/A gnd OAI21X1_628/Y vdd OAI21X1
XOAI21X1_639 BUFX4_126/Y OAI21X1_651/B OAI21X1_639/C gnd OAI21X1_639/Y vdd OAI21X1
XOAI21X1_617 INVX1_240/Y NOR2X1_133/Y NAND2X1_144/Y gnd OAI21X1_617/Y vdd OAI21X1
XDFFPOSX1_520 INVX1_477/A CLKBUF1_80/Y OAI21X1_240/Y gnd vdd DFFPOSX1
XMUX2X1_106 MUX2X1_106/A MUX2X1_106/B BUFX4_5/Y gnd MUX2X1_106/Y vdd MUX2X1
XMUX2X1_128 MUX2X1_128/A MUX2X1_128/B BUFX4_6/Y gnd MUX2X1_128/Y vdd MUX2X1
XMUX2X1_117 MUX2X1_117/A MUX2X1_117/B MUX2X1_84/S gnd AOI22X1_25/A vdd MUX2X1
XDFFPOSX1_531 INVX1_158/A CLKBUF1_1/Y OAI21X1_259/Y gnd vdd DFFPOSX1
XDFFPOSX1_553 NOR2X1_53/A CLKBUF1_1/Y AOI21X1_41/Y gnd vdd DFFPOSX1
XMUX2X1_139 MUX2X1_139/A MUX2X1_139/B BUFX4_58/Y gnd MUX2X1_139/Y vdd MUX2X1
XDFFPOSX1_564 INVX1_224/A CLKBUF1_46/Y OAI21X1_280/Y gnd vdd DFFPOSX1
XDFFPOSX1_542 NOR2X1_48/A CLKBUF1_57/Y AOI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_586 NOR2X1_64/A CLKBUF1_22/Y AOI21X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_597 INVX1_290/A CLKBUF1_79/Y OAI21X1_322/Y gnd vdd DFFPOSX1
XNAND2X1_601 BUFX4_200/Y NOR2X1_130/A gnd NAND2X1_601/Y vdd NAND2X1
XNAND2X1_612 BUFX4_222/Y NOR2X1_216/A gnd NAND2X1_612/Y vdd NAND2X1
XDFFPOSX1_575 NAND2X1_654/B CLKBUF1_57/Y OAI21X1_302/Y gnd vdd DFFPOSX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_13 a[5] gnd INVX1_13/Y vdd INVX1
XNAND2X1_634 BUFX4_260/Y NAND2X1_634/B gnd NAND2X1_634/Y vdd NAND2X1
XNAND2X1_645 MUX2X1_5/S NAND2X1_645/B gnd NAND2X1_645/Y vdd NAND2X1
XNAND2X1_623 BUFX4_240/Y NOR2X1_318/A gnd NAND2X1_623/Y vdd NAND2X1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XNAND2X1_656 BUFX4_203/Y NAND2X1_656/B gnd NAND2X1_656/Y vdd NAND2X1
XNAND2X1_678 BUFX4_245/Y NOR2X1_197/A gnd NAND2X1_678/Y vdd NAND2X1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XNAND2X1_667 AOI22X1_65/Y AOI22X1_66/Y gnd AOI22X1_69/A vdd NAND2X1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XNAND2X1_689 BUFX4_263/Y NOR2X1_293/A gnd NAND2X1_689/Y vdd NAND2X1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XDFFPOSX1_9 DFFPOSX1_9/Q CLKBUF1_23/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XFILL_40_6_1 gnd vdd FILL
XAOI21X1_280 BUFX4_113/Y NOR2X1_352/B NOR2X1_352/Y gnd AOI21X1_280/Y vdd AOI21X1
XAOI21X1_291 BUFX4_97/Y NOR2X1_367/B NOR2X1_365/Y gnd AOI21X1_291/Y vdd AOI21X1
XFILL_48_7_1 gnd vdd FILL
XFILL_47_2_0 gnd vdd FILL
XFILL_31_6_1 gnd vdd FILL
XFILL_30_1_0 gnd vdd FILL
XFILL_39_7_1 gnd vdd FILL
XFILL_38_2_0 gnd vdd FILL
XFILL_22_6_1 gnd vdd FILL
XOAI21X1_403 BUFX4_415/Y NOR2X1_61/A NAND2X1_589/B gnd OAI21X1_404/C vdd OAI21X1
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_414 INVX1_357/Y NOR2X1_71/Y NAND2X1_89/Y gnd OAI21X1_414/Y vdd OAI21X1
XOAI21X1_425 BUFX4_406/Y BUFX4_341/Y INVX1_294/A gnd OAI21X1_425/Y vdd OAI21X1
XOAI21X1_447 BUFX4_88/Y BUFX4_337/Y NAND2X1_729/B gnd OAI21X1_448/C vdd OAI21X1
XOAI21X1_436 BUFX4_419/Y NAND2X1_93/Y OAI21X1_436/C gnd OAI21X1_436/Y vdd OAI21X1
XOAI21X1_469 BUFX4_368/Y BUFX4_340/Y NAND2X1_385/B gnd OAI21X1_470/C vdd OAI21X1
XOAI21X1_458 BUFX4_401/Y NAND2X1_94/Y OAI21X1_458/C gnd OAI21X1_458/Y vdd OAI21X1
XDFFPOSX1_383 OAI21X1_61/C CLKBUF1_8/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_361 OAI21X1_17/C CLKBUF1_34/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_372 INVX1_212/A CLKBUF1_34/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_350 NAND2X1_570/B CLKBUF1_45/Y DFFPOSX1_350/D gnd vdd DFFPOSX1
XDFFPOSX1_394 NOR2X1_4/A CLKBUF1_94/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XNAND2X1_420 BUFX4_260/Y NOR2X1_336/A gnd OAI21X1_987/C vdd NAND2X1
XNAND2X1_453 BUFX4_223/Y OAI21X1_439/C gnd NAND2X1_453/Y vdd NAND2X1
XNAND2X1_431 MUX2X1_2/S NOR2X1_383/A gnd OAI21X1_997/C vdd NAND2X1
XNAND2X1_442 BUFX4_203/Y NOR2X1_36/A gnd NAND2X1_442/Y vdd NAND2X1
XFILL_5_7_1 gnd vdd FILL
XNAND2X1_475 BUFX4_265/Y NOR2X1_223/A gnd NAND2X1_475/Y vdd NAND2X1
XNAND2X1_464 BUFX4_243/Y NOR2X1_139/A gnd NAND2X1_464/Y vdd NAND2X1
XNAND2X1_497 BUFX4_204/Y NOR2X1_364/A gnd NAND2X1_497/Y vdd NAND2X1
XNAND2X1_486 MUX2X1_8/S NAND2X1_486/B gnd NAND2X1_486/Y vdd NAND2X1
XFILL_4_2_0 gnd vdd FILL
XFILL_29_2_0 gnd vdd FILL
XFILL_13_6_1 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_970 INVX1_182/Y BUFX4_227/Y NAND2X1_401/Y gnd MUX2X1_133/A vdd OAI21X1
XOAI21X1_981 INVX1_193/Y BUFX4_249/Y OAI21X1_981/C gnd MUX2X1_142/B vdd OAI21X1
XOAI21X1_992 INVX1_204/Y BUFX4_271/Y OAI21X1_992/C gnd MUX2X1_149/A vdd OAI21X1
XOAI21X1_63 BUFX4_415/Y BUFX4_314/Y OAI21X1_63/C gnd OAI21X1_64/C vdd OAI21X1
XOAI21X1_52 BUFX4_424/Y NAND2X1_4/Y OAI21X1_52/C gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_41 BUFX4_169/Y BUFX4_314/Y INVX1_276/A gnd OAI21X1_42/C vdd OAI21X1
XOAI21X1_30 BUFX4_283/Y NAND2X1_2/Y OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_74 BUFX4_127/Y OAI21X1_82/B OAI21X1_74/C gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_85 NOR2X1_41/B NOR2X1_2/A INVX1_406/A gnd OAI21X1_86/C vdd OAI21X1
XOAI21X1_96 BUFX4_297/Y OAI21X1_96/B OAI21X1_95/Y gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_200 BUFX4_375/Y NAND2X1_22/Y OAI21X1_200/C gnd OAI21X1_200/Y vdd OAI21X1
XOAI21X1_211 INVX1_155/Y NOR2X1_21/Y NAND2X1_33/Y gnd OAI21X1_211/Y vdd OAI21X1
XOAI21X1_222 INVX1_348/Y NOR2X1_31/Y NAND2X1_44/Y gnd OAI21X1_222/Y vdd OAI21X1
XOAI21X1_233 BUFX4_461/Y BUFX4_436/Y INVX1_285/A gnd OAI21X1_233/Y vdd OAI21X1
XOAI21X1_244 BUFX4_422/Y NAND2X1_49/Y OAI21X1_243/Y gnd OAI21X1_244/Y vdd OAI21X1
XOAI21X1_255 BUFX4_150/Y INVX2_2/A NAND2X1_720/B gnd OAI21X1_255/Y vdd OAI21X1
XOAI21X1_288 NAND2X1_66/Y BUFX4_379/Y OAI21X1_288/C gnd OAI21X1_288/Y vdd OAI21X1
XOAI21X1_266 INVX1_95/Y NOR2X1_51/Y NAND2X1_59/Y gnd OAI21X1_266/Y vdd OAI21X1
XOAI21X1_299 BUFX4_411/Y BUFX4_432/Y NAND2X1_585/B gnd OAI21X1_299/Y vdd OAI21X1
XOAI21X1_277 BUFX4_165/Y BUFX4_432/Y INVX1_160/A gnd OAI21X1_277/Y vdd OAI21X1
XINVX1_308 INVX1_308/A gnd INVX1_308/Y vdd INVX1
XINVX1_319 INVX1_319/A gnd INVX1_319/Y vdd INVX1
XDFFPOSX1_191 NAND2X1_628/B CLKBUF1_84/Y OAI21X1_1486/Y gnd vdd DFFPOSX1
XDFFPOSX1_180 INVX1_200/A CLKBUF1_84/Y DFFPOSX1_180/D gnd vdd DFFPOSX1
XNAND2X1_261 BUFX4_261/Y NAND2X1_261/B gnd NAND2X1_261/Y vdd NAND2X1
XNAND2X1_250 BUFX4_20/Y NAND2X1_250/B gnd AOI21X1_205/B vdd NAND2X1
XNAND2X1_283 BUFX4_204/Y NAND2X1_283/B gnd OAI21X1_860/C vdd NAND2X1
XNAND2X1_294 BUFX4_224/Y NAND2X1_294/B gnd NAND2X1_294/Y vdd NAND2X1
XNAND2X1_272 MUX2X1_4/S NOR2X1_257/A gnd NAND2X1_272/Y vdd NAND2X1
XFILL_45_5_1 gnd vdd FILL
XFILL_44_0_0 gnd vdd FILL
XOAI21X1_1518 BUFX4_282/Y NAND2X1_835/Y OAI21X1_1518/C gnd DFFPOSX1_207/D vdd OAI21X1
XOAI21X1_1529 BUFX4_405/Y BUFX4_91/Y INVX1_266/A gnd OAI21X1_1530/C vdd OAI21X1
XOAI21X1_1507 BUFX4_147/Y BUFX4_91/Y NAND2X1_284/B gnd OAI21X1_1508/C vdd OAI21X1
XFILL_6_1 gnd vdd FILL
XFILL_48_1 gnd vdd FILL
XFILL_36_5_1 gnd vdd FILL
XFILL_35_0_0 gnd vdd FILL
XCLKBUF1_42 BUFX4_12/Y gnd CLKBUF1_42/Y vdd CLKBUF1
XCLKBUF1_31 BUFX4_13/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XCLKBUF1_20 BUFX4_12/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XCLKBUF1_53 BUFX4_14/Y gnd CLKBUF1_53/Y vdd CLKBUF1
XCLKBUF1_64 BUFX4_17/Y gnd CLKBUF1_64/Y vdd CLKBUF1
XCLKBUF1_75 BUFX4_13/Y gnd CLKBUF1_75/Y vdd CLKBUF1
XCLKBUF1_86 BUFX4_16/Y gnd CLKBUF1_86/Y vdd CLKBUF1
XCLKBUF1_97 BUFX4_15/Y gnd CLKBUF1_97/Y vdd CLKBUF1
XFILL_2_5_1 gnd vdd FILL
XFILL_27_5_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_10_4_1 gnd vdd FILL
XINVX1_116 INVX1_116/A gnd INVX1_116/Y vdd INVX1
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XINVX1_138 INVX1_138/A gnd INVX1_138/Y vdd INVX1
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XBUFX4_403 INVX8_12/Y gnd BUFX4_403/Y vdd BUFX4
XBUFX4_436 BUFX4_436/A gnd BUFX4_436/Y vdd BUFX4
XBUFX4_414 INVX8_16/Y gnd BUFX4_414/Y vdd BUFX4
XBUFX4_447 d[4] gnd BUFX4_447/Y vdd BUFX4
XBUFX4_425 INVX8_3/Y gnd BUFX4_425/Y vdd BUFX4
XFILL_18_5_1 gnd vdd FILL
XBUFX4_458 INVX8_10/Y gnd NOR2X1_1/B vdd BUFX4
XFILL_17_0_0 gnd vdd FILL
XAOI21X1_109 BUFX4_421/Y NOR2X1_139/B NOR2X1_137/Y gnd AOI21X1_109/Y vdd AOI21X1
XOAI21X1_1304 INVX1_445/Y NOR2X1_254/Y NAND2X1_763/Y gnd DFFPOSX1_32/D vdd OAI21X1
XOAI21X1_1337 BUFX4_460/Y BUFX4_465/Y INVX1_257/A gnd OAI21X1_1338/C vdd OAI21X1
XDFFPOSX1_905 MUX2X1_15/A CLKBUF1_9/Y OAI21X1_692/Y gnd vdd DFFPOSX1
XOAI21X1_1326 INVX1_320/Y NOR2X1_284/Y NAND2X1_788/Y gnd DFFPOSX1_54/D vdd OAI21X1
XOAI21X1_1315 INVX1_127/Y NOR2X1_274/Y NAND2X1_777/Y gnd DFFPOSX1_35/D vdd OAI21X1
XOAI21X1_1359 BUFX4_154/Y BUFX4_468/Y NAND2X1_690/B gnd OAI21X1_1359/Y vdd OAI21X1
XDFFPOSX1_916 INVX1_246/A CLKBUF1_90/Y OAI21X1_709/Y gnd vdd DFFPOSX1
XDFFPOSX1_938 NOR2X1_192/A CLKBUF1_86/Y AOI21X1_154/Y gnd vdd DFFPOSX1
XDFFPOSX1_927 NOR2X1_186/A CLKBUF1_86/Y AOI21X1_150/Y gnd vdd DFFPOSX1
XOAI21X1_1348 BUFX4_420/Y NAND2X1_793/Y OAI21X1_1347/Y gnd DFFPOSX1_74/D vdd OAI21X1
XDFFPOSX1_949 INVX1_312/A CLKBUF1_44/Y OAI21X1_724/Y gnd vdd DFFPOSX1
XFILL_42_3_1 gnd vdd FILL
XBUFX4_211 BUFX4_26/Y gnd BUFX4_211/Y vdd BUFX4
XBUFX4_200 BUFX4_23/Y gnd BUFX4_200/Y vdd BUFX4
XBUFX4_255 BUFX4_24/Y gnd BUFX4_255/Y vdd BUFX4
XBUFX4_233 BUFX4_30/Y gnd BUFX4_233/Y vdd BUFX4
XBUFX4_222 BUFX4_23/Y gnd BUFX4_222/Y vdd BUFX4
XBUFX4_244 BUFX4_27/Y gnd BUFX4_244/Y vdd BUFX4
XNOR2X1_304 NOR2X1_304/A NOR2X1_303/B gnd NOR2X1_304/Y vdd NOR2X1
XBUFX4_266 BUFX4_31/Y gnd BUFX4_266/Y vdd BUFX4
XBUFX4_288 BUFX4_288/A gnd BUFX4_288/Y vdd BUFX4
XBUFX4_277 BUFX4_28/Y gnd BUFX4_277/Y vdd BUFX4
XNOR2X1_315 NOR2X1_315/A NOR2X1_315/B gnd NOR2X1_315/Y vdd NOR2X1
XNOR2X1_348 NOR2X1_348/A NOR2X1_342/B gnd NOR2X1_348/Y vdd NOR2X1
XNOR2X1_326 NOR2X1_326/A NOR2X1_325/B gnd NOR2X1_326/Y vdd NOR2X1
XNOR2X1_359 BUFX4_348/Y BUFX4_84/Y gnd NOR2X1_367/B vdd NOR2X1
XNOR2X1_337 NOR2X1_337/A NOR2X1_338/B gnd NOR2X1_337/Y vdd NOR2X1
XBUFX4_299 INVX8_5/Y gnd BUFX4_299/Y vdd BUFX4
XFILL_33_3_1 gnd vdd FILL
XOAI21X1_1101 INVX1_313/Y BUFX4_192/Y NAND2X1_542/Y gnd MUX2X1_232/B vdd OAI21X1
XOAI21X1_1112 INVX1_324/Y BUFX4_214/Y NAND2X1_555/Y gnd MUX2X1_239/A vdd OAI21X1
XDFFPOSX1_702 NAND2X1_593/B CLKBUF1_45/Y OAI21X1_508/Y gnd vdd DFFPOSX1
XOAI21X1_1134 INVX1_346/Y BUFX4_258/Y NAND2X1_578/Y gnd MUX2X1_256/A vdd OAI21X1
XOAI21X1_1156 INVX1_368/Y BUFX4_203/Y NAND2X1_602/Y gnd MUX2X1_272/A vdd OAI21X1
XOAI21X1_1145 INVX1_357/Y MUX2X1_2/S NAND2X1_590/Y gnd MUX2X1_265/B vdd OAI21X1
XDFFPOSX1_713 NAND2X1_267/B CLKBUF1_46/Y OAI21X1_530/Y gnd vdd DFFPOSX1
XOAI21X1_1123 INVX1_335/Y BUFX4_236/Y NAND2X1_567/Y gnd MUX2X1_248/B vdd OAI21X1
XOAI21X1_1189 INVX1_401/Y BUFX4_269/Y NAND2X1_638/Y gnd MUX2X1_298/B vdd OAI21X1
XOAI21X1_1167 INVX1_379/Y BUFX4_225/Y NAND2X1_613/Y gnd MUX2X1_281/B vdd OAI21X1
XDFFPOSX1_724 INVX1_234/A CLKBUF1_72/Y OAI21X1_548/Y gnd vdd DFFPOSX1
XDFFPOSX1_757 INVX1_300/A CLKBUF1_94/Y OAI21X1_565/Y gnd vdd DFFPOSX1
XDFFPOSX1_735 NOR2X1_89/A CLKBUF1_29/Y AOI21X1_71/Y gnd vdd DFFPOSX1
XOAI21X1_1178 INVX1_390/Y BUFX4_247/Y NAND2X1_626/Y gnd MUX2X1_289/A vdd OAI21X1
XDFFPOSX1_746 NOR2X1_94/A CLKBUF1_13/Y AOI21X1_74/Y gnd vdd DFFPOSX1
XINVX1_480 INVX1_480/A gnd INVX1_480/Y vdd INVX1
XDFFPOSX1_779 NAND2X1_392/B CLKBUF1_62/Y OAI21X1_590/Y gnd vdd DFFPOSX1
XDFFPOSX1_768 NOR2X1_110/A CLKBUF1_54/Y AOI21X1_88/Y gnd vdd DFFPOSX1
XNAND2X1_805 INVX8_5/A NOR2X1_309/Y gnd NAND2X1_805/Y vdd NAND2X1
XNAND2X1_816 BUFX4_163/Y NOR2X1_321/Y gnd NAND2X1_816/Y vdd NAND2X1
XNAND2X1_827 BUFX4_145/Y NOR2X1_331/Y gnd NAND2X1_827/Y vdd NAND2X1
XINVX1_491 INVX1_491/A gnd INVX1_491/Y vdd INVX1
XNAND2X1_838 INVX8_2/A NOR2X1_352/B gnd NAND2X1_838/Y vdd NAND2X1
XNAND2X1_849 BUFX4_326/Y NOR2X1_358/Y gnd NAND2X1_849/Y vdd NAND2X1
XFILL_24_3_1 gnd vdd FILL
XOAI21X1_1690 BUFX4_83/Y INVX2_11/A NAND2X1_220/B gnd OAI21X1_1691/C vdd OAI21X1
XFILL_7_4_1 gnd vdd FILL
XNOR2X1_11 BUFX4_135/Y NOR2X1_41/B gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_55 NOR2X1_55/A NOR2X1_55/B gnd NOR2X1_55/Y vdd NOR2X1
XNOR2X1_44 NOR2X1_44/A NOR2X1_43/B gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_33 NOR2X1_33/A NOR2X1_38/B gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_22 BUFX4_135/Y NOR2X1_22/B gnd NOR2X1_27/B vdd NOR2X1
XNOR2X1_66 NOR2X1_66/A NOR2X1_67/B gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_77 NOR2X1_77/A NOR2X1_77/B gnd NOR2X1_77/Y vdd NOR2X1
XNOR2X1_88 NOR2X1_88/A NOR2X1_90/B gnd NOR2X1_88/Y vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_99 NOR2X1_99/A NOR2X1_96/B gnd NOR2X1_99/Y vdd NOR2X1
XNOR2X1_123 MUX2X1_4/B NOR2X1_122/Y gnd NOR2X1_123/Y vdd NOR2X1
XMUX2X1_51 MUX2X1_51/A MUX2X1_51/B MUX2X1_84/S gnd MUX2X1_51/Y vdd MUX2X1
XNOR2X1_112 MUX2X1_2/B NOR2X1_111/Y gnd NOR2X1_112/Y vdd NOR2X1
XMUX2X1_62 MUX2X1_62/A MUX2X1_62/B BUFX4_38/Y gnd MUX2X1_63/A vdd MUX2X1
XMUX2X1_40 MUX2X1_40/A MUX2X1_40/B BUFX4_37/Y gnd MUX2X1_40/Y vdd MUX2X1
XNOR2X1_101 INVX1_2/A BUFX4_165/Y gnd NOR2X1_101/Y vdd NOR2X1
XNOR2X1_134 MUX2X1_5/B NOR2X1_133/Y gnd NOR2X1_134/Y vdd NOR2X1
XMUX2X1_73 MUX2X1_73/A MUX2X1_73/B BUFX4_22/Y gnd MUX2X1_75/B vdd MUX2X1
XMUX2X1_84 MUX2X1_84/A MUX2X1_84/B MUX2X1_84/S gnd MUX2X1_84/Y vdd MUX2X1
XNOR2X1_156 MUX2X1_11/B NOR2X1_155/Y gnd NOR2X1_156/Y vdd NOR2X1
XMUX2X1_95 MUX2X1_95/A MUX2X1_95/B BUFX4_19/Y gnd MUX2X1_96/A vdd MUX2X1
XNOR2X1_167 MUX2X1_12/B NOR2X1_166/Y gnd NOR2X1_167/Y vdd NOR2X1
XNOR2X1_145 MUX2X1_9/B NOR2X1_145/B gnd NOR2X1_145/Y vdd NOR2X1
XNOR2X1_189 MUX2X1_18/B NOR2X1_189/B gnd NOR2X1_189/Y vdd NOR2X1
XNOR2X1_178 MUX2X1_16/B NOR2X1_177/Y gnd NOR2X1_178/Y vdd NOR2X1
XOAI21X1_629 BUFX4_299/Y OAI21X1_635/B OAI21X1_628/Y gnd OAI21X1_629/Y vdd OAI21X1
XOAI21X1_618 INVX1_304/Y NOR2X1_133/Y OAI21X1_618/C gnd OAI21X1_618/Y vdd OAI21X1
XOAI21X1_607 INVX1_494/Y NOR2X1_111/Y OAI21X1_607/C gnd OAI21X1_607/Y vdd OAI21X1
XDFFPOSX1_521 OAI21X1_241/C CLKBUF1_1/Y OAI21X1_242/Y gnd vdd DFFPOSX1
XMUX2X1_118 MUX2X1_118/A MUX2X1_118/B BUFX4_20/Y gnd MUX2X1_120/B vdd MUX2X1
XMUX2X1_107 MUX2X1_107/A MUX2X1_107/B BUFX4_36/Y gnd MUX2X1_107/Y vdd MUX2X1
XDFFPOSX1_510 NOR2X1_38/A CLKBUF1_30/Y AOI21X1_30/Y gnd vdd DFFPOSX1
XMUX2X1_129 MUX2X1_128/Y MUX2X1_129/B MUX2X1_96/S gnd AOI22X1_27/A vdd MUX2X1
XDFFPOSX1_532 INVX1_222/A CLKBUF1_46/Y OAI21X1_260/Y gnd vdd DFFPOSX1
XDFFPOSX1_565 INVX1_288/A CLKBUF1_91/Y OAI21X1_282/Y gnd vdd DFFPOSX1
XDFFPOSX1_554 NOR2X1_54/A CLKBUF1_15/Y AOI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_543 NOR2X1_49/A CLKBUF1_57/Y AOI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_587 NOR2X1_65/A CLKBUF1_22/Y AOI21X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_598 INVX1_354/A CLKBUF1_79/Y OAI21X1_324/Y gnd vdd DFFPOSX1
XNAND2X1_602 BUFX4_202/Y NOR2X1_141/A gnd NAND2X1_602/Y vdd NAND2X1
XDFFPOSX1_576 OAI21X1_303/C CLKBUF1_82/Y OAI21X1_304/Y gnd vdd DFFPOSX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XNAND2X1_613 BUFX4_224/Y NOR2X1_225/A gnd NAND2X1_613/Y vdd NAND2X1
XNAND2X1_646 MUX2X1_9/S NAND2X1_646/B gnd NAND2X1_646/Y vdd NAND2X1
XNAND2X1_635 BUFX4_262/Y NOR2X1_366/A gnd NAND2X1_635/Y vdd NAND2X1
XNAND2X1_624 BUFX4_242/Y NAND2X1_624/B gnd NAND2X1_624/Y vdd NAND2X1
XNAND2X1_657 BUFX4_205/Y NAND2X1_657/B gnd NAND2X1_657/Y vdd NAND2X1
XNAND2X1_679 BUFX4_247/Y NOR2X1_208/A gnd NAND2X1_679/Y vdd NAND2X1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XNAND2X1_668 BUFX4_225/Y OAI21X1_597/C gnd NAND2X1_668/Y vdd NAND2X1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XAOI21X1_270 BUFX4_373/Y NOR2X1_338/B NOR2X1_340/Y gnd AOI21X1_270/Y vdd AOI21X1
XAOI21X1_281 BUFX4_303/Y NOR2X1_352/B NOR2X1_353/Y gnd AOI21X1_281/Y vdd AOI21X1
XAOI21X1_292 BUFX4_280/Y NOR2X1_367/B NOR2X1_366/Y gnd AOI21X1_292/Y vdd AOI21X1
XFILL_47_2_1 gnd vdd FILL
XFILL_30_1_1 gnd vdd FILL
XFILL_38_2_1 gnd vdd FILL
XOAI21X1_404 BUFX4_102/Y NAND2X1_82/Y OAI21X1_404/C gnd OAI21X1_404/Y vdd OAI21X1
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_426 BUFX4_401/Y NAND2X1_92/Y OAI21X1_425/Y gnd OAI21X1_426/Y vdd OAI21X1
XOAI21X1_448 BUFX4_378/Y NAND2X1_93/Y OAI21X1_448/C gnd OAI21X1_448/Y vdd OAI21X1
XOAI21X1_437 BUFX4_88/Y NOR2X1_72/A NAND2X1_384/B gnd OAI21X1_438/C vdd OAI21X1
XOAI21X1_415 INVX1_421/Y NOR2X1_71/Y NAND2X1_90/Y gnd OAI21X1_415/Y vdd OAI21X1
XOAI21X1_459 BUFX4_310/Y BUFX4_336/Y INVX1_359/A gnd OAI21X1_460/C vdd OAI21X1
XDFFPOSX1_340 INVX1_210/A CLKBUF1_28/Y DFFPOSX1_340/D gnd vdd DFFPOSX1
XDFFPOSX1_351 NAND2X1_639/B CLKBUF1_8/Y OAI21X1_1703/Y gnd vdd DFFPOSX1
XDFFPOSX1_373 INVX1_276/A CLKBUF1_34/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_362 OAI21X1_19/C CLKBUF1_8/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_384 OAI21X1_63/C CLKBUF1_28/Y OAI21X1_64/Y gnd vdd DFFPOSX1
XNAND2X1_410 BUFX4_240/Y NOR2X1_259/A gnd NAND2X1_410/Y vdd NAND2X1
XDFFPOSX1_395 NOR2X1_5/A CLKBUF1_75/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XNAND2X1_421 BUFX4_262/Y NAND2X1_421/B gnd OAI21X1_988/C vdd NAND2X1
XNAND2X1_432 MUX2X1_5/S NAND2X1_432/B gnd NAND2X1_432/Y vdd NAND2X1
XNAND2X1_454 BUFX4_225/Y NAND2X1_454/B gnd NAND2X1_454/Y vdd NAND2X1
XNAND2X1_443 AOI22X1_32/Y AOI22X1_33/Y gnd AOI22X1_34/D vdd NAND2X1
XNAND2X1_465 BUFX4_245/Y NAND2X1_465/B gnd NAND2X1_465/Y vdd NAND2X1
XNAND2X1_476 BUFX4_267/Y NOR2X1_234/A gnd NAND2X1_476/Y vdd NAND2X1
XNAND2X1_487 MUX2X1_11/S NAND2X1_487/B gnd NAND2X1_487/Y vdd NAND2X1
XFILL_4_2_1 gnd vdd FILL
XFILL_29_2_1 gnd vdd FILL
XNAND2X1_498 BUFX4_206/Y NOR2X1_374/A gnd NAND2X1_498/Y vdd NAND2X1
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_960 INVX1_172/Y BUFX4_207/Y OAI21X1_960/C gnd MUX2X1_125/A vdd OAI21X1
XOAI21X1_982 INVX1_194/Y BUFX4_251/Y OAI21X1_982/C gnd MUX2X1_142/A vdd OAI21X1
XOAI21X1_971 INVX1_183/Y BUFX4_229/Y NAND2X1_402/Y gnd MUX2X1_134/B vdd OAI21X1
XOAI21X1_993 INVX1_205/Y BUFX4_273/Y NAND2X1_427/Y gnd MUX2X1_151/B vdd OAI21X1
XOAI21X1_20 BUFX4_424/Y NAND2X1_2/Y OAI21X1_20/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_42 NAND2X1_3/Y BUFX4_401/Y OAI21X1_42/C gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_31 BUFX4_367/Y OAI21X1_7/B OAI21X1_31/C gnd OAI21X1_32/C vdd OAI21X1
XOAI21X1_53 BUFX4_414/Y BUFX4_319/Y OAI21X1_53/C gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_64 BUFX4_380/Y NAND2X1_4/Y OAI21X1_64/C gnd OAI21X1_64/Y vdd OAI21X1
XOAI21X1_75 NOR2X1_81/B NOR2X1_1/A INVX1_86/A gnd OAI21X1_76/C vdd OAI21X1
XOAI21X1_86 BUFX4_280/Y OAI21X1_82/B OAI21X1_86/C gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_97 BUFX4_84/Y NOR2X1_2/A OAI21X1_97/C gnd OAI21X1_98/C vdd OAI21X1
XOAI21X1_201 INVX1_31/Y NOR2X1_11/Y NAND2X1_23/Y gnd OAI21X1_201/Y vdd OAI21X1
XOAI21X1_212 INVX1_219/Y NOR2X1_21/Y NAND2X1_34/Y gnd OAI21X1_212/Y vdd OAI21X1
XOAI21X1_234 BUFX4_394/Y NAND2X1_48/Y OAI21X1_233/Y gnd OAI21X1_234/Y vdd OAI21X1
XOAI21X1_245 BUFX4_154/Y BUFX4_436/Y OAI21X1_245/C gnd OAI21X1_246/C vdd OAI21X1
XOAI21X1_256 BUFX4_379/Y NAND2X1_49/Y OAI21X1_255/Y gnd OAI21X1_256/Y vdd OAI21X1
XOAI21X1_223 INVX1_412/Y NOR2X1_31/Y NAND2X1_45/Y gnd OAI21X1_223/Y vdd OAI21X1
XOAI21X1_267 INVX1_159/Y NOR2X1_51/Y NAND2X1_60/Y gnd OAI21X1_267/Y vdd OAI21X1
XOAI21X1_278 NAND2X1_66/Y BUFX4_116/Y OAI21X1_277/Y gnd OAI21X1_278/Y vdd OAI21X1
XOAI21X1_289 BUFX4_411/Y BUFX4_433/Y NAND2X1_258/B gnd OAI21X1_290/C vdd OAI21X1
XINVX1_309 INVX1_309/A gnd INVX1_309/Y vdd INVX1
XDFFPOSX1_181 INVX1_264/A CLKBUF1_84/Y OAI21X1_1466/Y gnd vdd DFFPOSX1
XDFFPOSX1_170 NOR2X1_334/A CLKBUF1_93/Y AOI21X1_264/Y gnd vdd DFFPOSX1
XDFFPOSX1_192 NAND2X1_697/B CLKBUF1_78/Y OAI21X1_1488/Y gnd vdd DFFPOSX1
XNAND2X1_262 BUFX4_263/Y OAI21X1_393/C gnd OAI21X1_840/C vdd NAND2X1
XNAND2X1_251 BUFX4_245/Y NOR2X1_333/A gnd OAI21X1_830/C vdd NAND2X1
XNAND2X1_240 INVX4_1/Y NAND2X1_240/B gnd AOI21X1_203/A vdd NAND2X1
XNAND2X1_284 BUFX4_206/Y NAND2X1_284/B gnd OAI21X1_861/C vdd NAND2X1
XNAND2X1_273 MUX2X1_8/S NOR2X1_267/A gnd OAI21X1_850/C vdd NAND2X1
XNAND2X1_295 BUFX4_226/Y OAI21X1_19/C gnd NAND2X1_295/Y vdd NAND2X1
XFILL_44_0_1 gnd vdd FILL
XOAI21X1_1508 BUFX4_426/Y NAND2X1_835/Y OAI21X1_1508/C gnd DFFPOSX1_202/D vdd OAI21X1
XOAI21X1_1519 BUFX4_146/Y BUFX4_94/Y NAND2X1_698/B gnd OAI21X1_1519/Y vdd OAI21X1
XOAI21X1_790 BUFX4_308/Y BUFX4_438/Y INVX1_507/A gnd OAI21X1_791/C vdd OAI21X1
XFILL_6_2 gnd vdd FILL
XMUX2X1_290 MUX2X1_290/A MUX2X1_290/B BUFX4_80/Y gnd MUX2X1_291/A vdd MUX2X1
XFILL_35_0_1 gnd vdd FILL
XCLKBUF1_32 BUFX4_14/Y gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_10 BUFX4_17/Y gnd CLKBUF1_10/Y vdd CLKBUF1
XCLKBUF1_21 BUFX4_16/Y gnd CLKBUF1_21/Y vdd CLKBUF1
XCLKBUF1_43 BUFX4_12/Y gnd CLKBUF1_43/Y vdd CLKBUF1
XCLKBUF1_65 BUFX4_15/Y gnd CLKBUF1_65/Y vdd CLKBUF1
XCLKBUF1_54 BUFX4_9/Y gnd CLKBUF1_54/Y vdd CLKBUF1
XCLKBUF1_87 BUFX4_16/Y gnd CLKBUF1_87/Y vdd CLKBUF1
XCLKBUF1_76 BUFX4_17/Y gnd CLKBUF1_76/Y vdd CLKBUF1
XCLKBUF1_98 BUFX4_11/Y gnd CLKBUF1_98/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_26_0_1 gnd vdd FILL
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XINVX1_117 INVX1_117/A gnd INVX1_117/Y vdd INVX1
XINVX1_128 INVX1_128/A gnd INVX1_128/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XBUFX4_404 INVX8_12/Y gnd BUFX4_404/Y vdd BUFX4
XBUFX4_437 BUFX4_436/A gnd BUFX4_437/Y vdd BUFX4
XBUFX4_415 INVX8_16/Y gnd BUFX4_415/Y vdd BUFX4
XBUFX4_426 INVX8_3/Y gnd BUFX4_426/Y vdd BUFX4
XFILL_46_8_0 gnd vdd FILL
XBUFX4_459 INVX8_10/Y gnd NOR2X1_61/B vdd BUFX4
XBUFX4_448 d[4] gnd BUFX4_448/Y vdd BUFX4
XFILL_17_0_1 gnd vdd FILL
XOAI21X1_1305 INVX1_34/Y NOR2X1_264/Y NAND2X1_766/Y gnd DFFPOSX1_1/D vdd OAI21X1
XOAI21X1_1338 BUFX4_397/Y NAND2X1_792/Y OAI21X1_1338/C gnd DFFPOSX1_69/D vdd OAI21X1
XDFFPOSX1_906 OAI21X1_693/C CLKBUF1_21/Y OAI21X1_694/Y gnd vdd DFFPOSX1
XOAI21X1_1327 INVX1_384/Y NOR2X1_284/Y NAND2X1_789/Y gnd DFFPOSX1_55/D vdd OAI21X1
XOAI21X1_1316 INVX1_191/Y NOR2X1_274/Y NAND2X1_778/Y gnd DFFPOSX1_36/D vdd OAI21X1
XOAI21X1_1349 BUFX4_154/Y BUFX4_467/Y DFFPOSX1_75/Q gnd OAI21X1_1349/Y vdd OAI21X1
XDFFPOSX1_928 NOR2X1_187/A CLKBUF1_51/Y AOI21X1_151/Y gnd vdd DFFPOSX1
XDFFPOSX1_939 NOR2X1_193/A CLKBUF1_101/Y AOI21X1_155/Y gnd vdd DFFPOSX1
XDFFPOSX1_917 INVX1_310/A CLKBUF1_18/Y OAI21X1_710/Y gnd vdd DFFPOSX1
XFILL_37_8_0 gnd vdd FILL
XFILL_20_7_0 gnd vdd FILL
XFILL_3_8_0 gnd vdd FILL
XFILL_28_8_0 gnd vdd FILL
XFILL_11_7_0 gnd vdd FILL
XBUFX4_212 BUFX4_29/Y gnd BUFX4_212/Y vdd BUFX4
XBUFX4_201 BUFX4_30/Y gnd BUFX4_201/Y vdd BUFX4
XBUFX4_234 BUFX4_29/Y gnd BUFX4_234/Y vdd BUFX4
XFILL_19_8_0 gnd vdd FILL
XBUFX4_223 BUFX4_28/Y gnd BUFX4_223/Y vdd BUFX4
XBUFX4_245 BUFX4_27/Y gnd BUFX4_245/Y vdd BUFX4
XBUFX4_256 BUFX4_26/Y gnd BUFX4_256/Y vdd BUFX4
XBUFX4_289 BUFX4_288/A gnd INVX1_11/A vdd BUFX4
XBUFX4_278 BUFX4_23/Y gnd BUFX4_278/Y vdd BUFX4
XBUFX4_267 BUFX4_25/Y gnd BUFX4_267/Y vdd BUFX4
XNOR2X1_316 NOR2X1_316/A NOR2X1_315/B gnd NOR2X1_316/Y vdd NOR2X1
XNOR2X1_305 NOR2X1_305/A NOR2X1_303/B gnd NOR2X1_305/Y vdd NOR2X1
XNOR2X1_349 NOR2X1_349/A NOR2X1_342/B gnd NOR2X1_349/Y vdd NOR2X1
XNOR2X1_327 NOR2X1_327/A NOR2X1_325/B gnd NOR2X1_327/Y vdd NOR2X1
XNOR2X1_338 NOR2X1_338/A NOR2X1_338/B gnd NOR2X1_338/Y vdd NOR2X1
XOAI21X1_1102 INVX1_314/Y BUFX4_194/Y NAND2X1_543/Y gnd MUX2X1_232/A vdd OAI21X1
XOAI21X1_1113 INVX1_325/Y BUFX4_216/Y NAND2X1_556/Y gnd MUX2X1_241/B vdd OAI21X1
XOAI21X1_1146 INVX1_358/Y MUX2X1_5/S NAND2X1_591/Y gnd MUX2X1_265/A vdd OAI21X1
XDFFPOSX1_703 NAND2X1_662/B CLKBUF1_38/Y OAI21X1_510/Y gnd vdd DFFPOSX1
XOAI21X1_1135 INVX1_347/Y BUFX4_260/Y NAND2X1_579/Y gnd MUX2X1_257/B vdd OAI21X1
XDFFPOSX1_714 NAND2X1_318/B CLKBUF1_29/Y OAI21X1_532/Y gnd vdd DFFPOSX1
XOAI21X1_1124 INVX1_336/Y BUFX4_238/Y NAND2X1_568/Y gnd MUX2X1_248/A vdd OAI21X1
XOAI21X1_1168 INVX1_380/Y BUFX4_227/Y NAND2X1_614/Y gnd MUX2X1_281/A vdd OAI21X1
XDFFPOSX1_725 INVX1_298/A CLKBUF1_94/Y OAI21X1_549/Y gnd vdd DFFPOSX1
XDFFPOSX1_747 NOR2X1_95/A CLKBUF1_4/Y AOI21X1_75/Y gnd vdd DFFPOSX1
XOAI21X1_1179 INVX1_391/Y BUFX4_249/Y NAND2X1_627/Y gnd MUX2X1_290/B vdd OAI21X1
XDFFPOSX1_736 NOR2X1_90/A CLKBUF1_54/Y AOI21X1_72/Y gnd vdd DFFPOSX1
XOAI21X1_1157 INVX1_369/Y BUFX4_205/Y NAND2X1_603/Y gnd MUX2X1_274/B vdd OAI21X1
XINVX1_470 INVX1_470/A gnd INVX1_470/Y vdd INVX1
XDFFPOSX1_769 MUX2X1_1/B CLKBUF1_74/Y OAI21X1_570/Y gnd vdd DFFPOSX1
XDFFPOSX1_758 INVX1_364/A CLKBUF1_100/Y OAI21X1_566/Y gnd vdd DFFPOSX1
XINVX1_481 INVX1_481/A gnd INVX1_481/Y vdd INVX1
XNAND2X1_806 INVX8_6/A NOR2X1_309/Y gnd NAND2X1_806/Y vdd NAND2X1
XNAND2X1_817 BUFX4_452/Y NOR2X1_321/Y gnd NAND2X1_817/Y vdd NAND2X1
XNAND2X1_828 BUFX4_448/Y NOR2X1_331/Y gnd NAND2X1_828/Y vdd NAND2X1
XINVX1_492 INVX1_492/A gnd INVX1_492/Y vdd INVX1
XNAND2X1_839 INVX2_9/Y INVX4_3/Y gnd NAND2X1_839/Y vdd NAND2X1
XOAI21X1_1691 BUFX4_124/Y NAND2X1_872/Y OAI21X1_1691/C gnd DFFPOSX1_345/D vdd OAI21X1
XOAI21X1_1680 BUFX4_404/Y BUFX4_314/Y INVX1_210/A gnd OAI21X1_1680/Y vdd OAI21X1
XNOR2X1_12 BUFX4_133/Y BUFX4_87/Y gnd NOR2X1_14/B vdd NOR2X1
XNOR2X1_45 NOR2X1_45/A NOR2X1_43/B gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_38/B gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A NOR2X1_27/B gnd NOR2X1_23/Y vdd NOR2X1
XNOR2X1_56 NOR2X1_56/A NOR2X1_55/B gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_67 NOR2X1_67/A NOR2X1_67/B gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_78 NOR2X1_78/A NOR2X1_77/B gnd NOR2X1_78/Y vdd NOR2X1
XNOR2X1_89 NOR2X1_89/A NOR2X1_90/B gnd NOR2X1_89/Y vdd NOR2X1
XFILL_43_6_0 gnd vdd FILL
XMUX2X1_30 MUX2X1_30/A MUX2X1_30/B BUFX4_200/Y gnd MUX2X1_30/Y vdd MUX2X1
XMUX2X1_52 MUX2X1_52/A MUX2X1_52/B BUFX4_46/Y gnd MUX2X1_54/B vdd MUX2X1
XNOR2X1_124 BUFX4_105/Y NOR2X1_22/B gnd NOR2X1_126/B vdd NOR2X1
XNOR2X1_113 BUFX4_108/Y BUFX4_88/Y gnd NOR2X1_118/B vdd NOR2X1
XMUX2X1_63 MUX2X1_63/A MUX2X1_61/Y MUX2X1_96/S gnd MUX2X1_63/Y vdd MUX2X1
XMUX2X1_41 MUX2X1_41/A MUX2X1_41/B INVX4_1/A gnd MUX2X1_42/A vdd MUX2X1
XNOR2X1_102 INVX1_2/A BUFX4_411/Y gnd NOR2X1_103/B vdd NOR2X1
XMUX2X1_85 MUX2X1_85/A MUX2X1_85/B BUFX4_39/Y gnd MUX2X1_87/B vdd MUX2X1
XMUX2X1_74 MUX2X1_74/A MUX2X1_74/B BUFX4_47/Y gnd MUX2X1_74/Y vdd MUX2X1
XNOR2X1_135 BUFX4_105/Y NOR2X1_32/B gnd NOR2X1_139/B vdd NOR2X1
XFILL_34_6_0 gnd vdd FILL
XNOR2X1_146 BUFX4_118/Y BUFX4_86/Y gnd NOR2X1_153/B vdd NOR2X1
XMUX2X1_96 MUX2X1_96/A MUX2X1_96/B MUX2X1_96/S gnd MUX2X1_96/Y vdd MUX2X1
XNOR2X1_157 BUFX4_118/Y NOR2X1_52/B gnd NOR2X1_158/B vdd NOR2X1
XNOR2X1_179 BUFX4_64/Y BUFX4_87/Y gnd NOR2X1_186/B vdd NOR2X1
XNOR2X1_168 BUFX4_118/Y BUFX4_411/Y gnd NOR2X1_173/B vdd NOR2X1
XOAI21X1_619 INVX1_368/Y NOR2X1_133/Y OAI21X1_619/C gnd OAI21X1_619/Y vdd OAI21X1
XOAI21X1_608 INVX1_111/Y NOR2X1_122/Y OAI21X1_608/C gnd OAI21X1_608/Y vdd OAI21X1
XDFFPOSX1_522 NAND2X1_306/B CLKBUF1_19/Y OAI21X1_244/Y gnd vdd DFFPOSX1
XMUX2X1_119 MUX2X1_119/A MUX2X1_119/B BUFX4_45/Y gnd MUX2X1_119/Y vdd MUX2X1
XMUX2X1_108 MUX2X1_107/Y MUX2X1_106/Y MUX2X1_42/S gnd MUX2X1_108/Y vdd MUX2X1
XDFFPOSX1_500 INVX1_220/A CLKBUF1_31/Y OAI21X1_220/Y gnd vdd DFFPOSX1
XDFFPOSX1_511 NOR2X1_39/A CLKBUF1_37/Y AOI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_555 NOR2X1_55/A CLKBUF1_1/Y AOI21X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_533 INVX1_286/A CLKBUF1_11/Y OAI21X1_261/Y gnd vdd DFFPOSX1
XDFFPOSX1_544 NOR2X1_50/A CLKBUF1_57/Y AOI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_566 INVX1_352/A CLKBUF1_19/Y OAI21X1_284/Y gnd vdd DFFPOSX1
XDFFPOSX1_599 INVX1_418/A CLKBUF1_79/Y OAI21X1_326/Y gnd vdd DFFPOSX1
XDFFPOSX1_588 NOR2X1_66/A CLKBUF1_34/Y AOI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_577 INVX1_49/A CLKBUF1_3/Y OAI21X1_305/Y gnd vdd DFFPOSX1
XNAND2X1_603 BUFX4_204/Y NAND2X1_603/B gnd NAND2X1_603/Y vdd NAND2X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XNAND2X1_614 BUFX4_226/Y NOR2X1_236/A gnd NAND2X1_614/Y vdd NAND2X1
XNAND2X1_625 BUFX4_244/Y NAND2X1_625/B gnd NAND2X1_625/Y vdd NAND2X1
XNAND2X1_636 BUFX4_264/Y NOR2X1_376/A gnd NAND2X1_636/Y vdd NAND2X1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XNAND2X1_658 BUFX4_207/Y NAND2X1_658/B gnd NAND2X1_658/Y vdd NAND2X1
XNAND2X1_647 MUX2X1_12/S NOR2X1_19/A gnd NAND2X1_647/Y vdd NAND2X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XNAND2X1_669 BUFX4_227/Y NOR2X1_120/A gnd NAND2X1_669/Y vdd NAND2X1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XFILL_0_6_0 gnd vdd FILL
XFILL_25_6_0 gnd vdd FILL
XAOI21X1_260 BUFX4_99/Y NOR2X1_325/B NOR2X1_328/Y gnd AOI21X1_260/Y vdd AOI21X1
XAOI21X1_282 BUFX4_398/Y NOR2X1_352/B NOR2X1_354/Y gnd AOI21X1_282/Y vdd AOI21X1
XAOI21X1_271 BUFX4_128/Y NOR2X1_342/B NOR2X1_342/Y gnd AOI21X1_271/Y vdd AOI21X1
XAOI21X1_293 BUFX4_379/Y NOR2X1_367/B NOR2X1_367/Y gnd AOI21X1_293/Y vdd AOI21X1
XFILL_8_7_0 gnd vdd FILL
XFILL_16_6_0 gnd vdd FILL
XOAI21X1_405 BUFX4_414/Y BUFX4_381/Y NAND2X1_658/B gnd OAI21X1_405/Y vdd OAI21X1
XOAI21X1_427 BUFX4_403/Y BUFX4_341/Y INVX1_358/A gnd OAI21X1_428/C vdd OAI21X1
XOAI21X1_438 BUFX4_117/Y NAND2X1_93/Y OAI21X1_438/C gnd OAI21X1_438/Y vdd OAI21X1
XOAI21X1_416 INVX1_485/Y NOR2X1_71/Y NAND2X1_91/Y gnd OAI21X1_416/Y vdd OAI21X1
XOAI21X1_449 BUFX4_310/Y BUFX4_341/Y INVX1_55/A gnd OAI21X1_450/C vdd OAI21X1
XDFFPOSX1_330 NOR2X1_381/A CLKBUF1_69/Y AOI21X1_303/Y gnd vdd DFFPOSX1
XDFFPOSX1_363 OAI21X1_21/C CLKBUF1_16/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_341 INVX1_274/A CLKBUF1_99/Y DFFPOSX1_341/D gnd vdd DFFPOSX1
XDFFPOSX1_352 NAND2X1_708/B CLKBUF1_16/Y DFFPOSX1_352/D gnd vdd DFFPOSX1
XDFFPOSX1_374 INVX1_340/A CLKBUF1_34/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XNAND2X1_400 BUFX4_224/Y NAND2X1_400/B gnd NAND2X1_400/Y vdd NAND2X1
XNAND2X1_411 BUFX4_242/Y NOR2X1_269/A gnd NAND2X1_411/Y vdd NAND2X1
XDFFPOSX1_385 INVX1_28/A CLKBUF1_93/Y OAI21X1_65/Y gnd vdd DFFPOSX1
XDFFPOSX1_396 NOR2X1_6/A CLKBUF1_72/Y AOI21X1_4/Y gnd vdd DFFPOSX1
XNAND2X1_433 MUX2X1_9/S OAI21X1_23/C gnd NAND2X1_433/Y vdd NAND2X1
XNAND2X1_422 BUFX4_264/Y NAND2X1_422/B gnd NAND2X1_422/Y vdd NAND2X1
XNAND2X1_444 BUFX4_205/Y NAND2X1_444/B gnd NAND2X1_444/Y vdd NAND2X1
XNAND2X1_455 BUFX4_227/Y NAND2X1_455/B gnd NAND2X1_455/Y vdd NAND2X1
XNAND2X1_477 AOI22X1_37/Y AOI22X1_38/Y gnd AOI22X1_39/D vdd NAND2X1
XNAND2X1_488 BUFX4_188/Y NOR2X1_327/A gnd NAND2X1_488/Y vdd NAND2X1
XNAND2X1_466 BUFX4_247/Y NOR2X1_150/A gnd NAND2X1_466/Y vdd NAND2X1
XNAND2X1_499 BUFX4_208/Y NAND2X1_499/B gnd NAND2X1_499/Y vdd NAND2X1
XFILL_40_4_0 gnd vdd FILL
XOAI21X1_950 INVX1_162/Y MUX2X1_12/S NAND2X1_380/Y gnd MUX2X1_118/A vdd OAI21X1
XOAI21X1_961 INVX1_173/Y BUFX4_209/Y NAND2X1_392/Y gnd MUX2X1_127/B vdd OAI21X1
XOAI21X1_972 INVX1_184/Y BUFX4_231/Y NAND2X1_403/Y gnd MUX2X1_134/A vdd OAI21X1
XOAI21X1_994 INVX1_206/Y BUFX4_275/Y OAI21X1_994/C gnd MUX2X1_151/A vdd OAI21X1
XOAI21X1_983 INVX1_195/Y BUFX4_253/Y OAI21X1_983/C gnd MUX2X1_143/B vdd OAI21X1
XFILL_48_5_0 gnd vdd FILL
XOAI21X1_10 BUFX4_401/Y NAND2X1_1/Y OAI21X1_9/Y gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_21 BUFX4_368/Y BUFX4_319/Y OAI21X1_21/C gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_32 BUFX4_380/Y NAND2X1_2/Y OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_54 BUFX4_109/Y NAND2X1_4/Y OAI21X1_53/Y gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_43 BUFX4_169/Y OAI21X1_7/B INVX1_340/A gnd OAI21X1_44/C vdd OAI21X1
XFILL_31_4_0 gnd vdd FILL
XOAI21X1_65 INVX1_28/Y NOR2X1_1/Y NAND2X1_6/Y gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_87 NOR2X1_81/B INVX2_1/A INVX1_470/A gnd OAI21X1_88/C vdd OAI21X1
XOAI21X1_76 BUFX4_425/Y OAI21X1_82/B OAI21X1_76/C gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_98 BUFX4_399/Y OAI21X1_96/B OAI21X1_98/C gnd OAI21X1_98/Y vdd OAI21X1
XFILL_39_5_0 gnd vdd FILL
XFILL_22_4_0 gnd vdd FILL
XOAI21X1_202 INVX1_90/Y NOR2X1_11/Y NAND2X1_24/Y gnd OAI21X1_202/Y vdd OAI21X1
XOAI21X1_213 INVX1_283/Y NOR2X1_21/Y NAND2X1_35/Y gnd OAI21X1_213/Y vdd OAI21X1
XOAI21X1_246 BUFX4_114/Y NAND2X1_49/Y OAI21X1_246/C gnd OAI21X1_246/Y vdd OAI21X1
XOAI21X1_235 BUFX4_461/Y BUFX4_437/Y INVX1_349/A gnd OAI21X1_235/Y vdd OAI21X1
XOAI21X1_224 INVX1_476/Y NOR2X1_31/Y NAND2X1_46/Y gnd OAI21X1_224/Y vdd OAI21X1
XOAI21X1_257 INVX1_46/Y NOR2X1_41/Y NAND2X1_50/Y gnd OAI21X1_257/Y vdd OAI21X1
XOAI21X1_268 INVX1_223/Y NOR2X1_51/Y NAND2X1_61/Y gnd OAI21X1_268/Y vdd OAI21X1
XOAI21X1_279 BUFX4_165/Y BUFX4_433/Y INVX1_224/A gnd OAI21X1_279/Y vdd OAI21X1
XDFFPOSX1_182 INVX1_328/A CLKBUF1_42/Y OAI21X1_1468/Y gnd vdd DFFPOSX1
XDFFPOSX1_171 NOR2X1_335/A CLKBUF1_63/Y AOI21X1_265/Y gnd vdd DFFPOSX1
XDFFPOSX1_160 NOR2X1_330/A CLKBUF1_68/Y AOI21X1_262/Y gnd vdd DFFPOSX1
XDFFPOSX1_193 MUX2X1_29/B CLKBUF1_36/Y OAI21X1_1490/Y gnd vdd DFFPOSX1
XNAND2X1_241 BUFX4_235/Y NOR2X1_300/A gnd OAI21X1_824/C vdd NAND2X1
XNAND2X1_230 AOI22X1_3/Y AOI22X1_6/Y gnd AOI21X1_200/B vdd NAND2X1
XNAND2X1_252 INVX4_1/Y NAND2X1_252/B gnd NAND2X1_252/Y vdd NAND2X1
XNAND2X1_285 BUFX4_208/Y NOR2X1_343/A gnd OAI21X1_862/C vdd NAND2X1
XFILL_5_5_0 gnd vdd FILL
XNAND2X1_296 BUFX4_228/Y OAI21X1_51/C gnd NAND2X1_296/Y vdd NAND2X1
XNAND2X1_274 MUX2X1_11/S NOR2X1_277/A gnd OAI21X1_851/C vdd NAND2X1
XNAND2X1_263 BUFX4_265/Y NOR2X1_73/A gnd OAI21X1_841/C vdd NAND2X1
XFILL_13_4_0 gnd vdd FILL
XOAI21X1_1509 BUFX4_146/Y BUFX4_89/Y NAND2X1_353/B gnd OAI21X1_1510/C vdd OAI21X1
XOAI21X1_791 BUFX4_378/Y NAND2X1_201/Y OAI21X1_791/C gnd OAI21X1_791/Y vdd OAI21X1
XOAI21X1_780 NOR2X1_91/B BUFX4_441/Y INVX1_187/A gnd OAI21X1_780/Y vdd OAI21X1
XMUX2X1_280 MUX2X1_280/A MUX2X1_280/B BUFX4_48/Y gnd MUX2X1_282/B vdd MUX2X1
XMUX2X1_291 MUX2X1_291/A MUX2X1_291/B BUFX4_364/Y gnd AOI22X1_61/A vdd MUX2X1
XCLKBUF1_11 BUFX4_14/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XCLKBUF1_22 BUFX4_17/Y gnd CLKBUF1_22/Y vdd CLKBUF1
XCLKBUF1_33 BUFX4_9/Y gnd CLKBUF1_33/Y vdd CLKBUF1
XCLKBUF1_66 BUFX4_17/Y gnd CLKBUF1_66/Y vdd CLKBUF1
XCLKBUF1_44 BUFX4_11/Y gnd CLKBUF1_44/Y vdd CLKBUF1
XCLKBUF1_55 BUFX4_12/Y gnd CLKBUF1_55/Y vdd CLKBUF1
XCLKBUF1_99 BUFX4_10/Y gnd CLKBUF1_99/Y vdd CLKBUF1
XCLKBUF1_88 BUFX4_9/Y gnd CLKBUF1_88/Y vdd CLKBUF1
XCLKBUF1_77 BUFX4_14/Y gnd CLKBUF1_77/Y vdd CLKBUF1
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XBUFX4_405 INVX8_12/Y gnd BUFX4_405/Y vdd BUFX4
XBUFX4_438 BUFX4_439/A gnd BUFX4_438/Y vdd BUFX4
XBUFX4_427 d[7] gnd BUFX4_427/Y vdd BUFX4
XBUFX4_416 INVX8_16/Y gnd BUFX4_416/Y vdd BUFX4
XFILL_46_8_1 gnd vdd FILL
XBUFX4_449 d[1] gnd BUFX4_449/Y vdd BUFX4
XFILL_45_3_0 gnd vdd FILL
XOAI21X1_1306 INVX1_62/Y NOR2X1_264/Y NAND2X1_767/Y gnd DFFPOSX1_2/D vdd OAI21X1
XOAI21X1_1317 INVX1_255/Y NOR2X1_274/Y NAND2X1_779/Y gnd DFFPOSX1_37/D vdd OAI21X1
XOAI21X1_1328 INVX1_448/Y NOR2X1_284/Y NAND2X1_790/Y gnd DFFPOSX1_56/D vdd OAI21X1
XOAI21X1_1339 BUFX4_454/Y BUFX4_468/Y INVX1_321/A gnd OAI21X1_1339/Y vdd OAI21X1
XDFFPOSX1_929 MUX2X1_18/B CLKBUF1_14/Y AOI21X1_152/Y gnd vdd DFFPOSX1
XDFFPOSX1_907 NAND2X1_400/B CLKBUF1_9/Y OAI21X1_696/Y gnd vdd DFFPOSX1
XDFFPOSX1_918 INVX1_374/A CLKBUF1_87/Y OAI21X1_711/Y gnd vdd DFFPOSX1
XFILL_37_8_1 gnd vdd FILL
XFILL_36_3_0 gnd vdd FILL
XFILL_20_7_1 gnd vdd FILL
XFILL_3_8_1 gnd vdd FILL
XFILL_28_8_1 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_27_3_0 gnd vdd FILL
XFILL_11_7_1 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XBUFX4_202 BUFX4_28/Y gnd BUFX4_202/Y vdd BUFX4
XBUFX4_213 BUFX4_24/Y gnd BUFX4_213/Y vdd BUFX4
XBUFX4_235 BUFX4_29/Y gnd BUFX4_235/Y vdd BUFX4
XBUFX4_246 BUFX4_29/Y gnd BUFX4_246/Y vdd BUFX4
XFILL_19_8_1 gnd vdd FILL
XBUFX4_224 BUFX4_23/Y gnd BUFX4_224/Y vdd BUFX4
XBUFX4_268 BUFX4_29/Y gnd BUFX4_268/Y vdd BUFX4
XFILL_18_3_0 gnd vdd FILL
XBUFX4_257 BUFX4_31/Y gnd BUFX4_257/Y vdd BUFX4
XBUFX4_279 INVX8_8/Y gnd BUFX4_279/Y vdd BUFX4
XNOR2X1_306 NOR2X1_306/A NOR2X1_303/B gnd NOR2X1_306/Y vdd NOR2X1
XNOR2X1_328 NOR2X1_328/A NOR2X1_325/B gnd NOR2X1_328/Y vdd NOR2X1
XNOR2X1_339 NOR2X1_339/A NOR2X1_338/B gnd NOR2X1_339/Y vdd NOR2X1
XNOR2X1_317 NOR2X1_317/A NOR2X1_315/B gnd NOR2X1_317/Y vdd NOR2X1
XOAI21X1_1103 INVX1_315/Y BUFX4_196/Y NAND2X1_544/Y gnd MUX2X1_233/B vdd OAI21X1
XDFFPOSX1_704 NAND2X1_731/B CLKBUF1_47/Y OAI21X1_512/Y gnd vdd DFFPOSX1
XOAI21X1_1147 INVX1_359/Y MUX2X1_9/S NAND2X1_592/Y gnd MUX2X1_266/B vdd OAI21X1
XOAI21X1_1125 INVX1_337/Y BUFX4_240/Y NAND2X1_569/Y gnd MUX2X1_250/B vdd OAI21X1
XOAI21X1_1136 INVX1_348/Y BUFX4_262/Y NAND2X1_580/Y gnd MUX2X1_257/A vdd OAI21X1
XOAI21X1_1114 INVX1_326/Y BUFX4_218/Y NAND2X1_557/Y gnd MUX2X1_241/A vdd OAI21X1
XOAI21X1_1169 INVX1_381/Y BUFX4_229/Y NAND2X1_617/Y gnd MUX2X1_283/B vdd OAI21X1
XDFFPOSX1_726 INVX1_362/A CLKBUF1_94/Y OAI21X1_550/Y gnd vdd DFFPOSX1
XDFFPOSX1_715 NAND2X1_387/B CLKBUF1_26/Y OAI21X1_534/Y gnd vdd DFFPOSX1
XDFFPOSX1_748 NOR2X1_96/A CLKBUF1_26/Y AOI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_737 INVX1_59/A CLKBUF1_39/Y OAI21X1_553/Y gnd vdd DFFPOSX1
XOAI21X1_1158 INVX1_370/Y BUFX4_207/Y NAND2X1_604/Y gnd MUX2X1_274/A vdd OAI21X1
XINVX1_460 INVX1_460/A gnd INVX1_460/Y vdd INVX1
XDFFPOSX1_759 INVX1_428/A CLKBUF1_4/Y OAI21X1_567/Y gnd vdd DFFPOSX1
XINVX1_471 INVX1_471/A gnd INVX1_471/Y vdd INVX1
XINVX1_482 INVX1_482/A gnd INVX1_482/Y vdd INVX1
XNAND2X1_807 INVX8_7/A NOR2X1_309/Y gnd NAND2X1_807/Y vdd NAND2X1
XINVX1_493 INVX1_493/A gnd INVX1_493/Y vdd INVX1
XNAND2X1_818 BUFX4_334/Y NOR2X1_321/Y gnd NAND2X1_818/Y vdd NAND2X1
XNAND2X1_829 BUFX4_330/Y NOR2X1_331/Y gnd NAND2X1_829/Y vdd NAND2X1
XOAI21X1_1670 INVX1_273/Y NOR2X1_378/Y NAND2X1_867/Y gnd DFFPOSX1_325/D vdd OAI21X1
XOAI21X1_1681 BUFX4_300/Y NAND2X1_871/Y OAI21X1_1680/Y gnd DFFPOSX1_340/D vdd OAI21X1
XOAI21X1_1692 BUFX4_85/Y BUFX4_319/Y NAND2X1_294/B gnd OAI21X1_1693/C vdd OAI21X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_43/B gnd NOR2X1_46/Y vdd NOR2X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_14/B gnd NOR2X1_13/Y vdd NOR2X1
XNOR2X1_24 NOR2X1_24/A NOR2X1_27/B gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_35 NOR2X1_35/A NOR2X1_38/B gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_68 NOR2X1_68/A NOR2X1_67/B gnd NOR2X1_68/Y vdd NOR2X1
XNOR2X1_79 NOR2X1_79/A NOR2X1_77/B gnd NOR2X1_79/Y vdd NOR2X1
XNOR2X1_57 NOR2X1_57/A NOR2X1_55/B gnd NOR2X1_57/Y vdd NOR2X1
XFILL_43_6_1 gnd vdd FILL
XFILL_42_1_0 gnd vdd FILL
XMUX2X1_20 MUX2X1_19/Y MUX2X1_20/B BUFX4_48/Y gnd MUX2X1_21/A vdd MUX2X1
XMUX2X1_53 MUX2X1_53/A MUX2X1_53/B BUFX4_62/Y gnd MUX2X1_53/Y vdd MUX2X1
XNOR2X1_114 MUX2X1_2/A NOR2X1_118/B gnd NOR2X1_114/Y vdd NOR2X1
XMUX2X1_42 MUX2X1_42/A MUX2X1_40/Y MUX2X1_42/S gnd AOI22X1_8/D vdd MUX2X1
XNOR2X1_103 NOR2X1_103/A NOR2X1_103/B gnd AOI21X1_81/C vdd NOR2X1
XMUX2X1_31 MUX2X1_31/A MUX2X1_31/B BUFX4_61/Y gnd MUX2X1_33/B vdd MUX2X1
XNOR2X1_147 MUX2X1_9/A NOR2X1_153/B gnd NOR2X1_147/Y vdd NOR2X1
XNOR2X1_158 MUX2X1_11/A NOR2X1_158/B gnd NOR2X1_158/Y vdd NOR2X1
XMUX2X1_86 MUX2X1_86/A MUX2X1_86/B INVX4_1/A gnd MUX2X1_86/Y vdd MUX2X1
XNOR2X1_136 MUX2X1_5/A NOR2X1_139/B gnd NOR2X1_136/Y vdd NOR2X1
XMUX2X1_64 MUX2X1_64/A MUX2X1_64/B INVX4_1/A gnd MUX2X1_64/Y vdd MUX2X1
XMUX2X1_75 MUX2X1_74/Y MUX2X1_75/B MUX2X1_42/S gnd MUX2X1_75/Y vdd MUX2X1
XNOR2X1_125 MUX2X1_4/A NOR2X1_126/B gnd NOR2X1_125/Y vdd NOR2X1
XMUX2X1_97 MUX2X1_97/A MUX2X1_97/B BUFX4_44/Y gnd MUX2X1_99/B vdd MUX2X1
XFILL_34_6_1 gnd vdd FILL
XFILL_33_1_0 gnd vdd FILL
XNOR2X1_169 MUX2X1_12/A NOR2X1_173/B gnd NOR2X1_169/Y vdd NOR2X1
XOAI21X1_609 INVX1_175/Y NOR2X1_122/Y OAI21X1_609/C gnd OAI21X1_609/Y vdd OAI21X1
XDFFPOSX1_523 OAI21X1_245/C CLKBUF1_91/Y OAI21X1_246/Y gnd vdd DFFPOSX1
XDFFPOSX1_501 INVX1_284/A CLKBUF1_44/Y OAI21X1_221/Y gnd vdd DFFPOSX1
XDFFPOSX1_512 NOR2X1_40/A CLKBUF1_30/Y AOI21X1_32/Y gnd vdd DFFPOSX1
XMUX2X1_109 MUX2X1_109/A MUX2X1_109/B INVX4_1/A gnd MUX2X1_111/B vdd MUX2X1
XDFFPOSX1_556 NOR2X1_56/A CLKBUF1_95/Y AOI21X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_545 INVX1_47/A CLKBUF1_11/Y OAI21X1_265/Y gnd vdd DFFPOSX1
XDFFPOSX1_534 INVX1_350/A CLKBUF1_19/Y OAI21X1_262/Y gnd vdd DFFPOSX1
XDFFPOSX1_567 INVX1_416/A CLKBUF1_80/Y OAI21X1_286/Y gnd vdd DFFPOSX1
XDFFPOSX1_589 NOR2X1_67/A CLKBUF1_10/Y AOI21X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_578 INVX1_97/A CLKBUF1_83/Y OAI21X1_306/Y gnd vdd DFFPOSX1
XINVX1_290 INVX1_290/A gnd INVX1_290/Y vdd INVX1
XNAND2X1_615 AOI22X1_57/Y AOI22X1_58/Y gnd AOI22X1_59/D vdd NAND2X1
XNAND2X1_626 BUFX4_246/Y NOR2X1_329/A gnd NAND2X1_626/Y vdd NAND2X1
XNAND2X1_604 BUFX4_206/Y NOR2X1_152/A gnd NAND2X1_604/Y vdd NAND2X1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XNAND2X1_648 BUFX4_189/Y NOR2X1_29/A gnd NAND2X1_648/Y vdd NAND2X1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XNAND2X1_659 BUFX4_209/Y NOR2X1_79/A gnd NAND2X1_659/Y vdd NAND2X1
XNAND2X1_637 BUFX4_266/Y NAND2X1_637/B gnd NAND2X1_637/Y vdd NAND2X1
XNAND2X1_90 INVX8_8/A NOR2X1_71/Y gnd NAND2X1_90/Y vdd NAND2X1
XFILL_0_6_1 gnd vdd FILL
XFILL_25_6_1 gnd vdd FILL
XFILL_24_1_0 gnd vdd FILL
XAOI21X1_261 BUFX4_279/Y NOR2X1_325/B NOR2X1_329/Y gnd AOI21X1_261/Y vdd AOI21X1
XAOI21X1_250 BUFX4_297/Y NOR2X1_315/B NOR2X1_315/Y gnd AOI21X1_250/Y vdd AOI21X1
XAOI21X1_272 BUFX4_426/Y NOR2X1_342/B NOR2X1_343/Y gnd AOI21X1_272/Y vdd AOI21X1
XAOI21X1_283 BUFX4_96/Y NOR2X1_352/B NOR2X1_355/Y gnd AOI21X1_283/Y vdd AOI21X1
XAOI21X1_294 AOI21X1_1/A NOR2X1_373/B NOR2X1_370/Y gnd AOI21X1_294/Y vdd AOI21X1
XFILL_8_7_1 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XFILL_16_6_1 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XDFFPOSX1_1030 BUFX2_6/A CLKBUF1_65/Y NAND2X1_616/Y gnd vdd DFFPOSX1
XOAI21X1_439 BUFX4_83/Y INVX2_4/A OAI21X1_439/C gnd OAI21X1_440/C vdd OAI21X1
XOAI21X1_406 BUFX4_283/Y NAND2X1_82/Y OAI21X1_405/Y gnd OAI21X1_406/Y vdd OAI21X1
XOAI21X1_428 BUFX4_101/Y NAND2X1_92/Y OAI21X1_428/C gnd OAI21X1_428/Y vdd OAI21X1
XOAI21X1_417 BUFX4_403/Y BUFX4_337/Y INVX1_54/A gnd OAI21X1_418/C vdd OAI21X1
XDFFPOSX1_331 NOR2X1_382/A CLKBUF1_73/Y AOI21X1_304/Y gnd vdd DFFPOSX1
XDFFPOSX1_320 NAND2X1_706/B CLKBUF1_53/Y OAI21X1_1665/Y gnd vdd DFFPOSX1
XDFFPOSX1_353 INVX1_22/A CLKBUF1_22/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_364 OAI21X1_23/C CLKBUF1_16/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_342 INVX1_338/A CLKBUF1_45/Y DFFPOSX1_342/D gnd vdd DFFPOSX1
XNAND2X1_401 BUFX4_226/Y NOR2X1_182/A gnd NAND2X1_401/Y vdd NAND2X1
XDFFPOSX1_375 INVX1_404/A CLKBUF1_64/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_386 INVX1_85/A CLKBUF1_94/Y OAI21X1_66/Y gnd vdd DFFPOSX1
XDFFPOSX1_397 NOR2X1_7/A CLKBUF1_89/Y AOI21X1_5/Y gnd vdd DFFPOSX1
XNAND2X1_434 MUX2X1_12/S OAI21X1_55/C gnd NAND2X1_434/Y vdd NAND2X1
XNAND2X1_423 BUFX4_266/Y NOR2X1_345/A gnd OAI21X1_990/C vdd NAND2X1
XNAND2X1_412 BUFX4_244/Y NOR2X1_279/A gnd NAND2X1_412/Y vdd NAND2X1
XNAND2X1_445 BUFX4_207/Y NOR2X1_46/A gnd NAND2X1_445/Y vdd NAND2X1
XNAND2X1_467 BUFX4_249/Y NOR2X1_161/A gnd NAND2X1_467/Y vdd NAND2X1
XNAND2X1_478 AOI22X1_34/Y AOI22X1_39/Y gnd NAND2X1_478/Y vdd NAND2X1
XNAND2X1_456 BUFX4_229/Y NAND2X1_456/B gnd NAND2X1_456/Y vdd NAND2X1
XNAND2X1_489 BUFX4_190/Y NOR2X1_337/A gnd NAND2X1_489/Y vdd NAND2X1
XFILL_40_4_1 gnd vdd FILL
XOAI21X1_951 INVX1_163/Y BUFX4_189/Y NAND2X1_381/Y gnd MUX2X1_119/B vdd OAI21X1
XOAI21X1_940 INVX1_152/Y BUFX4_266/Y OAI21X1_940/C gnd MUX2X1_110/A vdd OAI21X1
XOAI21X1_973 INVX1_185/Y BUFX4_233/Y OAI21X1_973/C gnd MUX2X1_136/B vdd OAI21X1
XOAI21X1_962 INVX1_174/Y BUFX4_211/Y OAI21X1_962/C gnd MUX2X1_127/A vdd OAI21X1
XOAI21X1_984 INVX1_196/Y BUFX4_255/Y OAI21X1_984/C gnd MUX2X1_143/A vdd OAI21X1
XOAI21X1_995 INVX1_207/Y BUFX4_277/Y OAI21X1_995/C gnd MUX2X1_152/B vdd OAI21X1
XFILL_48_5_1 gnd vdd FILL
XFILL_47_0_0 gnd vdd FILL
XOAI21X1_11 BUFX4_307/Y BUFX4_314/Y INVX1_339/A gnd OAI21X1_12/C vdd OAI21X1
XOAI21X1_33 BUFX4_171/Y OAI21X1_1/B INVX1_21/A gnd OAI21X1_34/C vdd OAI21X1
XOAI21X1_22 BUFX4_109/Y NAND2X1_2/Y OAI21X1_21/Y gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_44 NAND2X1_3/Y BUFX4_101/Y OAI21X1_44/C gnd OAI21X1_44/Y vdd OAI21X1
XFILL_31_4_1 gnd vdd FILL
XOAI21X1_55 BUFX4_415/Y OAI21X1_7/B OAI21X1_55/C gnd OAI21X1_56/C vdd OAI21X1
XOAI21X1_66 INVX1_85/Y NOR2X1_1/Y NAND2X1_7/Y gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_77 NOR2X1_81/B NOR2X1_1/A INVX1_150/A gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_88 BUFX4_374/Y OAI21X1_82/B OAI21X1_88/C gnd OAI21X1_88/Y vdd OAI21X1
XOAI21X1_99 BUFX4_86/Y NOR2X1_1/A OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XFILL_39_5_1 gnd vdd FILL
XFILL_38_0_0 gnd vdd FILL
XFILL_22_4_1 gnd vdd FILL
XOAI21X1_203 INVX1_154/Y NOR2X1_11/Y NAND2X1_25/Y gnd OAI21X1_203/Y vdd OAI21X1
XOAI21X1_225 BUFX4_461/Y BUFX4_436/Y INVX1_45/A gnd OAI21X1_226/C vdd OAI21X1
XOAI21X1_236 BUFX4_97/Y NAND2X1_48/Y OAI21X1_235/Y gnd OAI21X1_236/Y vdd OAI21X1
XOAI21X1_214 INVX1_347/Y NOR2X1_21/Y NAND2X1_36/Y gnd OAI21X1_214/Y vdd OAI21X1
XOAI21X1_247 BUFX4_150/Y INVX2_2/A NAND2X1_444/B gnd OAI21X1_248/C vdd OAI21X1
XOAI21X1_269 INVX1_287/Y NOR2X1_51/Y NAND2X1_62/Y gnd OAI21X1_269/Y vdd OAI21X1
XOAI21X1_258 INVX1_94/Y NOR2X1_41/Y NAND2X1_51/Y gnd OAI21X1_258/Y vdd OAI21X1
XDFFPOSX1_150 INVX1_326/A CLKBUF1_63/Y DFFPOSX1_150/D gnd vdd DFFPOSX1
XDFFPOSX1_161 INVX1_43/A CLKBUF1_63/Y OAI21X1_1449/Y gnd vdd DFFPOSX1
XDFFPOSX1_172 NOR2X1_336/A CLKBUF1_61/Y AOI21X1_266/Y gnd vdd DFFPOSX1
XDFFPOSX1_183 INVX1_392/A CLKBUF1_78/Y OAI21X1_1470/Y gnd vdd DFFPOSX1
XNAND2X1_220 BUFX4_209/Y NAND2X1_220/B gnd NAND2X1_220/Y vdd NAND2X1
XDFFPOSX1_194 INVX1_73/A CLKBUF1_36/Y DFFPOSX1_194/D gnd vdd DFFPOSX1
XNAND2X1_231 DFFPOSX1_9/Q BUFX4_225/Y gnd OAI21X1_818/C vdd NAND2X1
XNAND2X1_242 BUFX4_41/Y NAND2X1_242/B gnd AOI21X1_203/B vdd NAND2X1
XNAND2X1_253 BUFX4_247/Y NAND2X1_253/B gnd OAI21X1_831/C vdd NAND2X1
XNAND2X1_286 BUFX4_210/Y NOR2X1_351/A gnd NAND2X1_286/Y vdd NAND2X1
XFILL_5_5_1 gnd vdd FILL
XNAND2X1_264 BUFX4_267/Y NAND2X1_264/B gnd NAND2X1_264/Y vdd NAND2X1
XNAND2X1_275 BUFX4_188/Y NOR2X1_287/A gnd NAND2X1_275/Y vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XNAND2X1_297 BUFX4_230/Y NOR2X1_4/A gnd NAND2X1_297/Y vdd NAND2X1
XFILL_29_0_0 gnd vdd FILL
XFILL_13_4_1 gnd vdd FILL
XOAI21X1_792 INVX1_124/Y NOR2X1_228/Y OAI21X1_792/C gnd OAI21X1_792/Y vdd OAI21X1
XOAI21X1_781 BUFX4_117/Y NAND2X1_201/Y OAI21X1_780/Y gnd OAI21X1_781/Y vdd OAI21X1
XOAI21X1_770 BUFX4_409/Y INVX2_5/A INVX1_378/A gnd OAI21X1_770/Y vdd OAI21X1
XMUX2X1_292 MUX2X1_292/A MUX2X1_292/B BUFX4_81/Y gnd MUX2X1_292/Y vdd MUX2X1
XMUX2X1_281 MUX2X1_281/A MUX2X1_281/B BUFX4_1/Y gnd MUX2X1_282/A vdd MUX2X1
XMUX2X1_270 MUX2X1_270/A MUX2X1_270/B BUFX4_357/Y gnd AOI22X1_56/D vdd MUX2X1
XCLKBUF1_23 BUFX4_16/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XCLKBUF1_12 BUFX4_11/Y gnd CLKBUF1_12/Y vdd CLKBUF1
XCLKBUF1_34 BUFX4_10/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XCLKBUF1_45 BUFX4_10/Y gnd CLKBUF1_45/Y vdd CLKBUF1
XCLKBUF1_56 BUFX4_13/Y gnd CLKBUF1_56/Y vdd CLKBUF1
XCLKBUF1_78 BUFX4_12/Y gnd CLKBUF1_78/Y vdd CLKBUF1
XCLKBUF1_67 BUFX4_15/Y gnd CLKBUF1_67/Y vdd CLKBUF1
XCLKBUF1_89 BUFX4_13/Y gnd CLKBUF1_89/Y vdd CLKBUF1
XINVX1_119 INVX1_119/A gnd INVX1_119/Y vdd INVX1
XINVX1_108 INVX1_108/A gnd INVX1_108/Y vdd INVX1
XBUFX4_406 INVX8_12/Y gnd BUFX4_406/Y vdd BUFX4
XBUFX4_428 d[7] gnd BUFX4_428/Y vdd BUFX4
XBUFX4_417 INVX8_16/Y gnd BUFX4_417/Y vdd BUFX4
XBUFX4_439 BUFX4_439/A gnd INVX2_5/A vdd BUFX4
XFILL_45_3_1 gnd vdd FILL
XOAI21X1_1329 BUFX4_460/Y BUFX4_465/Y INVX1_37/A gnd OAI21X1_1329/Y vdd OAI21X1
XOAI21X1_1307 INVX1_126/Y NOR2X1_264/Y NAND2X1_768/Y gnd DFFPOSX1_3/D vdd OAI21X1
XOAI21X1_1318 INVX1_319/Y NOR2X1_274/Y NAND2X1_780/Y gnd DFFPOSX1_38/D vdd OAI21X1
XDFFPOSX1_908 NAND2X1_469/B CLKBUF1_51/Y OAI21X1_698/Y gnd vdd DFFPOSX1
XDFFPOSX1_919 INVX1_438/A CLKBUF1_18/Y OAI21X1_712/Y gnd vdd DFFPOSX1
XFILL_4_1 gnd vdd FILL
XFILL_46_1 gnd vdd FILL
XFILL_36_3_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_27_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XBUFX4_203 BUFX4_30/Y gnd BUFX4_203/Y vdd BUFX4
XBUFX4_225 BUFX4_24/Y gnd BUFX4_225/Y vdd BUFX4
XBUFX4_214 BUFX4_31/Y gnd BUFX4_214/Y vdd BUFX4
XBUFX4_236 BUFX4_23/Y gnd BUFX4_236/Y vdd BUFX4
XNOR2X1_307 NOR2X1_307/A NOR2X1_303/B gnd NOR2X1_307/Y vdd NOR2X1
XBUFX4_258 BUFX4_24/Y gnd BUFX4_258/Y vdd BUFX4
XBUFX4_269 BUFX4_30/Y gnd BUFX4_269/Y vdd BUFX4
XFILL_18_3_1 gnd vdd FILL
XBUFX4_247 BUFX4_26/Y gnd BUFX4_247/Y vdd BUFX4
XNOR2X1_329 NOR2X1_329/A NOR2X1_325/B gnd NOR2X1_329/Y vdd NOR2X1
XNOR2X1_318 NOR2X1_318/A NOR2X1_315/B gnd NOR2X1_318/Y vdd NOR2X1
XOAI21X1_1104 INVX1_316/Y INVX8_1/A NAND2X1_545/Y gnd MUX2X1_233/A vdd OAI21X1
XDFFPOSX1_705 INVX1_57/A CLKBUF1_95/Y OAI21X1_514/Y gnd vdd DFFPOSX1
XOAI21X1_1126 INVX1_338/Y BUFX4_242/Y NAND2X1_570/Y gnd MUX2X1_250/A vdd OAI21X1
XOAI21X1_1115 INVX1_327/Y BUFX4_220/Y NAND2X1_558/Y gnd MUX2X1_242/B vdd OAI21X1
XOAI21X1_1137 INVX1_349/Y BUFX4_264/Y NAND2X1_582/Y gnd MUX2X1_259/B vdd OAI21X1
XOAI21X1_1148 INVX1_360/Y MUX2X1_12/S NAND2X1_593/Y gnd MUX2X1_266/A vdd OAI21X1
XDFFPOSX1_727 INVX1_426/A CLKBUF1_4/Y OAI21X1_551/Y gnd vdd DFFPOSX1
XDFFPOSX1_716 NAND2X1_456/B CLKBUF1_82/Y OAI21X1_536/Y gnd vdd DFFPOSX1
XDFFPOSX1_738 INVX1_107/A CLKBUF1_92/Y OAI21X1_554/Y gnd vdd DFFPOSX1
XOAI21X1_1159 INVX1_371/Y BUFX4_209/Y NAND2X1_605/Y gnd MUX2X1_275/B vdd OAI21X1
XDFFPOSX1_749 NOR2X1_97/A CLKBUF1_29/Y AOI21X1_77/Y gnd vdd DFFPOSX1
XINVX1_461 INVX1_461/A gnd INVX1_461/Y vdd INVX1
XINVX1_450 INVX1_450/A gnd INVX1_450/Y vdd INVX1
XINVX1_483 INVX1_483/A gnd INVX1_483/Y vdd INVX1
XNAND2X1_808 INVX8_8/A NOR2X1_309/Y gnd NAND2X1_808/Y vdd NAND2X1
XNAND2X1_819 BUFX4_144/Y NOR2X1_321/Y gnd NAND2X1_819/Y vdd NAND2X1
XINVX1_472 INVX1_472/A gnd INVX1_472/Y vdd INVX1
XINVX1_494 INVX1_494/A gnd INVX1_494/Y vdd INVX1
XOAI21X1_1660 BUFX4_412/Y BUFX4_343/Y NAND2X1_568/B gnd OAI21X1_1660/Y vdd OAI21X1
XOAI21X1_1682 BUFX4_406/Y OAI21X1_5/B INVX1_274/A gnd OAI21X1_1683/C vdd OAI21X1
XOAI21X1_1693 BUFX4_421/Y NAND2X1_872/Y OAI21X1_1693/C gnd OAI21X1_1693/Y vdd OAI21X1
XOAI21X1_1671 INVX1_337/Y NOR2X1_378/Y NAND2X1_868/Y gnd OAI21X1_1671/Y vdd OAI21X1
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_36 NOR2X1_36/A NOR2X1_38/B gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A NOR2X1_27/B gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_47 NOR2X1_47/A NOR2X1_43/B gnd NOR2X1_47/Y vdd NOR2X1
XNOR2X1_69 NOR2X1_69/A NOR2X1_67/B gnd NOR2X1_69/Y vdd NOR2X1
XNOR2X1_58 NOR2X1_58/A NOR2X1_55/B gnd NOR2X1_58/Y vdd NOR2X1
XFILL_42_1_1 gnd vdd FILL
XMUX2X1_10 MUX2X1_9/Y MUX2X1_8/Y BUFX4_19/Y gnd MUX2X1_14/B vdd MUX2X1
XMUX2X1_21 MUX2X1_21/A MUX2X1_17/Y BUFX4_357/Y gnd MUX2X1_21/Y vdd MUX2X1
XMUX2X1_54 MUX2X1_53/Y MUX2X1_54/B BUFX4_362/Y gnd MUX2X1_54/Y vdd MUX2X1
XMUX2X1_43 MUX2X1_43/A MUX2X1_43/B BUFX4_80/Y gnd MUX2X1_43/Y vdd MUX2X1
XNOR2X1_115 NOR2X1_115/A NOR2X1_118/B gnd NOR2X1_115/Y vdd NOR2X1
XMUX2X1_32 MUX2X1_32/A MUX2X1_32/B BUFX4_49/Y gnd MUX2X1_33/A vdd MUX2X1
XNOR2X1_104 NOR2X1_104/A NOR2X1_103/B gnd NOR2X1_104/Y vdd NOR2X1
XNOR2X1_137 NOR2X1_137/A NOR2X1_139/B gnd NOR2X1_137/Y vdd NOR2X1
XMUX2X1_87 MUX2X1_86/Y MUX2X1_87/B BUFX4_362/Y gnd MUX2X1_87/Y vdd MUX2X1
XMUX2X1_65 MUX2X1_65/A MUX2X1_65/B BUFX4_80/Y gnd MUX2X1_66/A vdd MUX2X1
XMUX2X1_76 MUX2X1_76/A MUX2X1_76/B BUFX4_63/Y gnd MUX2X1_76/Y vdd MUX2X1
XNOR2X1_126 NOR2X1_126/A NOR2X1_126/B gnd NOR2X1_126/Y vdd NOR2X1
XNOR2X1_148 NOR2X1_148/A NOR2X1_153/B gnd NOR2X1_148/Y vdd NOR2X1
XMUX2X1_98 MUX2X1_98/A MUX2X1_98/B BUFX4_60/Y gnd MUX2X1_99/A vdd MUX2X1
XFILL_33_1_1 gnd vdd FILL
XNOR2X1_159 NOR2X1_159/A NOR2X1_158/B gnd NOR2X1_159/Y vdd NOR2X1
XDFFPOSX1_513 INVX1_45/A CLKBUF1_91/Y OAI21X1_226/Y gnd vdd DFFPOSX1
XDFFPOSX1_502 INVX1_348/A CLKBUF1_31/Y OAI21X1_222/Y gnd vdd DFFPOSX1
XDFFPOSX1_546 INVX1_95/A CLKBUF1_46/Y OAI21X1_266/Y gnd vdd DFFPOSX1
XDFFPOSX1_535 INVX1_414/A CLKBUF1_27/Y OAI21X1_263/Y gnd vdd DFFPOSX1
XDFFPOSX1_524 NAND2X1_444/B CLKBUF1_57/Y OAI21X1_248/Y gnd vdd DFFPOSX1
XDFFPOSX1_568 INVX1_480/A CLKBUF1_80/Y OAI21X1_288/Y gnd vdd DFFPOSX1
XDFFPOSX1_579 INVX1_161/A CLKBUF1_10/Y OAI21X1_307/Y gnd vdd DFFPOSX1
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XDFFPOSX1_557 NOR2X1_57/A CLKBUF1_11/Y AOI21X1_45/Y gnd vdd DFFPOSX1
XINVX1_291 INVX1_291/A gnd INVX1_291/Y vdd INVX1
XNAND2X1_616 AOI22X1_54/Y AOI22X1_59/Y gnd NAND2X1_616/Y vdd NAND2X1
XNAND2X1_627 BUFX4_248/Y NOR2X1_339/A gnd NAND2X1_627/Y vdd NAND2X1
XNAND2X1_605 BUFX4_208/Y NOR2X1_163/A gnd NAND2X1_605/Y vdd NAND2X1
XNAND2X1_638 BUFX4_268/Y NOR2X1_386/A gnd NAND2X1_638/Y vdd NAND2X1
XNAND2X1_649 BUFX4_191/Y NOR2X1_39/A gnd NAND2X1_649/Y vdd NAND2X1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XNAND2X1_80 INVX2_3/Y INVX8_15/A gnd NAND2X1_80/Y vdd NAND2X1
XNAND2X1_91 INVX8_9/A NOR2X1_71/Y gnd NAND2X1_91/Y vdd NAND2X1
XFILL_24_1_1 gnd vdd FILL
XAOI21X1_251 BUFX4_394/Y NOR2X1_315/B NOR2X1_316/Y gnd AOI21X1_251/Y vdd AOI21X1
XAOI21X1_240 BUFX4_420/Y NOR2X1_303/B NOR2X1_301/Y gnd DFFPOSX1_90/D vdd AOI21X1
XAOI21X1_273 BUFX4_115/Y NOR2X1_342/B NOR2X1_344/Y gnd AOI21X1_273/Y vdd AOI21X1
XAOI21X1_284 BUFX4_282/Y NOR2X1_352/B NOR2X1_356/Y gnd AOI21X1_284/Y vdd AOI21X1
XAOI21X1_262 BUFX4_373/Y NOR2X1_325/B NOR2X1_330/Y gnd AOI21X1_262/Y vdd AOI21X1
XAOI21X1_295 BUFX4_420/Y NOR2X1_373/B NOR2X1_371/Y gnd AOI21X1_295/Y vdd AOI21X1
XOAI21X1_1490 BUFX4_128/Y NAND2X1_834/Y OAI21X1_1489/Y gnd OAI21X1_1490/Y vdd OAI21X1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XDFFPOSX1_1020 NOR2X1_234/A CLKBUF1_70/Y AOI21X1_190/Y gnd vdd DFFPOSX1
XDFFPOSX1_1031 BUFX2_7/A CLKBUF1_88/Y NAND2X1_685/Y gnd vdd DFFPOSX1
XOAI21X1_429 BUFX4_403/Y BUFX4_342/Y INVX1_422/A gnd OAI21X1_430/C vdd OAI21X1
XOAI21X1_418 BUFX4_124/Y NAND2X1_92/Y OAI21X1_418/C gnd OAI21X1_418/Y vdd OAI21X1
XOAI21X1_407 NOR2X1_32/B BUFX4_385/Y OAI21X1_407/C gnd OAI21X1_408/C vdd OAI21X1
XDFFPOSX1_310 INVX1_336/A CLKBUF1_32/Y DFFPOSX1_310/D gnd vdd DFFPOSX1
XDFFPOSX1_321 INVX1_24/A CLKBUF1_10/Y OAI21X1_1666/Y gnd vdd DFFPOSX1
XDFFPOSX1_343 INVX1_402/A CLKBUF1_22/Y OAI21X1_1687/Y gnd vdd DFFPOSX1
XDFFPOSX1_354 INVX1_83/A CLKBUF1_8/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_365 OAI21X1_25/C CLKBUF1_16/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_332 NOR2X1_383/A CLKBUF1_73/Y AOI21X1_305/Y gnd vdd DFFPOSX1
XNAND2X1_402 BUFX4_228/Y NOR2X1_193/A gnd NAND2X1_402/Y vdd NAND2X1
XDFFPOSX1_376 INVX1_468/A CLKBUF1_34/Y OAI21X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_387 INVX1_149/A CLKBUF1_4/Y OAI21X1_67/Y gnd vdd DFFPOSX1
XDFFPOSX1_398 NOR2X1_8/A CLKBUF1_94/Y AOI21X1_6/Y gnd vdd DFFPOSX1
XNAND2X1_424 BUFX4_268/Y NOR2X1_353/A gnd OAI21X1_991/C vdd NAND2X1
XNAND2X1_413 BUFX4_246/Y NOR2X1_289/A gnd OAI21X1_980/C vdd NAND2X1
XNAND2X1_435 BUFX4_189/Y NOR2X1_6/A gnd NAND2X1_435/Y vdd NAND2X1
XNAND2X1_468 BUFX4_251/Y NOR2X1_172/A gnd NAND2X1_468/Y vdd NAND2X1
XNAND2X1_457 BUFX4_231/Y NOR2X1_86/A gnd NAND2X1_457/Y vdd NAND2X1
XNAND2X1_446 BUFX4_209/Y NOR2X1_56/A gnd NAND2X1_446/Y vdd NAND2X1
XNAND2X1_479 BUFX4_269/Y NOR2X1_260/A gnd NAND2X1_479/Y vdd NAND2X1
XOAI21X1_952 INVX1_164/Y BUFX4_191/Y OAI21X1_952/C gnd MUX2X1_119/A vdd OAI21X1
XOAI21X1_941 INVX1_153/Y BUFX4_268/Y NAND2X1_370/Y gnd MUX2X1_112/B vdd OAI21X1
XOAI21X1_930 INVX1_142/Y BUFX4_246/Y NAND2X1_359/Y gnd MUX2X1_103/A vdd OAI21X1
XOAI21X1_974 INVX1_186/Y BUFX4_235/Y OAI21X1_974/C gnd MUX2X1_136/A vdd OAI21X1
XOAI21X1_985 INVX1_197/Y BUFX4_257/Y OAI21X1_985/C gnd MUX2X1_145/B vdd OAI21X1
XOAI21X1_963 INVX1_175/Y BUFX4_213/Y OAI21X1_963/C gnd MUX2X1_128/B vdd OAI21X1
XOAI21X1_996 INVX1_208/Y MUX2X1_1/S OAI21X1_996/C gnd MUX2X1_152/A vdd OAI21X1
XFILL_47_0_1 gnd vdd FILL
XOAI21X1_34 NAND2X1_3/Y BUFX4_128/Y OAI21X1_34/C gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_45 BUFX4_171/Y OAI21X1_1/B INVX1_404/A gnd OAI21X1_46/C vdd OAI21X1
XOAI21X1_12 BUFX4_101/Y NAND2X1_1/Y OAI21X1_12/C gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_23 BUFX4_368/Y BUFX4_319/Y OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_56 BUFX4_300/Y NAND2X1_4/Y OAI21X1_56/C gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_67 INVX1_149/Y NOR2X1_1/Y NAND2X1_8/Y gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_78 BUFX4_110/Y OAI21X1_82/B OAI21X1_77/Y gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_89 BUFX4_84/Y NOR2X1_2/A OAI21X1_89/C gnd OAI21X1_90/C vdd OAI21X1
XFILL_38_0_1 gnd vdd FILL
XOAI21X1_204 INVX1_218/Y NOR2X1_11/Y NAND2X1_26/Y gnd OAI21X1_204/Y vdd OAI21X1
XOAI21X1_226 BUFX4_126/Y NAND2X1_48/Y OAI21X1_226/C gnd OAI21X1_226/Y vdd OAI21X1
XOAI21X1_237 BUFX4_461/Y BUFX4_434/Y INVX1_413/A gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_215 INVX1_411/Y NOR2X1_21/Y NAND2X1_37/Y gnd OAI21X1_215/Y vdd OAI21X1
XOAI21X1_259 INVX1_158/Y NOR2X1_41/Y NAND2X1_52/Y gnd OAI21X1_259/Y vdd OAI21X1
XOAI21X1_248 BUFX4_297/Y NAND2X1_49/Y OAI21X1_248/C gnd OAI21X1_248/Y vdd OAI21X1
XDFFPOSX1_151 INVX1_390/A CLKBUF1_98/Y DFFPOSX1_151/D gnd vdd DFFPOSX1
XDFFPOSX1_162 INVX1_71/A CLKBUF1_61/Y DFFPOSX1_162/D gnd vdd DFFPOSX1
XDFFPOSX1_173 NOR2X1_337/A CLKBUF1_12/Y AOI21X1_267/Y gnd vdd DFFPOSX1
XDFFPOSX1_140 NAND2X1_418/B CLKBUF1_61/Y OAI21X1_1432/Y gnd vdd DFFPOSX1
XDFFPOSX1_184 INVX1_456/A CLKBUF1_78/Y DFFPOSX1_184/D gnd vdd DFFPOSX1
XDFFPOSX1_195 INVX1_137/A CLKBUF1_51/Y DFFPOSX1_195/D gnd vdd DFFPOSX1
XNAND2X1_210 MUX2X1_48/S BUFX4_5/Y gnd OR2X2_1/A vdd NAND2X1
XNAND2X1_221 BUFX4_211/Y NOR2X1_380/A gnd NAND2X1_221/Y vdd NAND2X1
XNAND2X1_232 INVX4_1/Y NAND2X1_232/B gnd AOI21X1_201/A vdd NAND2X1
XNAND2X1_243 BUFX4_237/Y NOR2X1_312/A gnd OAI21X1_825/C vdd NAND2X1
XNAND2X1_287 BUFX4_212/Y NAND2X1_287/B gnd NAND2X1_287/Y vdd NAND2X1
XNAND2X1_265 BUFX4_269/Y NAND2X1_265/B gnd NAND2X1_265/Y vdd NAND2X1
XNAND2X1_254 BUFX4_45/Y NAND2X1_254/B gnd AOI21X1_206/B vdd NAND2X1
XNAND2X1_276 BUFX4_190/Y NAND2X1_276/B gnd NAND2X1_276/Y vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XFILL_29_0_1 gnd vdd FILL
XNAND2X1_298 BUFX4_232/Y OAI21X1_91/C gnd OAI21X1_874/C vdd NAND2X1
XFILL_41_7_0 gnd vdd FILL
XOAI21X1_760 BUFX4_409/Y BUFX4_440/Y MUX2X1_23/B gnd OAI21X1_761/C vdd OAI21X1
XOAI21X1_782 BUFX4_308/Y BUFX4_443/Y INVX1_251/A gnd OAI21X1_782/Y vdd OAI21X1
XOAI21X1_793 INVX1_188/Y NOR2X1_228/Y OAI21X1_793/C gnd OAI21X1_793/Y vdd OAI21X1
XOAI21X1_771 BUFX4_103/Y OAI21X1_761/B OAI21X1_770/Y gnd OAI21X1_771/Y vdd OAI21X1
XMUX2X1_293 MUX2X1_293/A MUX2X1_293/B BUFX4_82/Y gnd MUX2X1_293/Y vdd MUX2X1
XMUX2X1_282 MUX2X1_282/A MUX2X1_282/B MUX2X1_84/S gnd AOI22X1_58/D vdd MUX2X1
XMUX2X1_271 MUX2X1_271/A MUX2X1_271/B BUFX4_82/Y gnd MUX2X1_273/B vdd MUX2X1
XMUX2X1_260 MUX2X1_260/A MUX2X1_260/B BUFX4_35/Y gnd MUX2X1_261/A vdd MUX2X1
XFILL_32_7_0 gnd vdd FILL
XCLKBUF1_24 BUFX4_11/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XCLKBUF1_13 BUFX4_9/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XCLKBUF1_46 BUFX4_18/Y gnd CLKBUF1_46/Y vdd CLKBUF1
XCLKBUF1_57 BUFX4_18/Y gnd CLKBUF1_57/Y vdd CLKBUF1
XCLKBUF1_35 BUFX4_17/Y gnd CLKBUF1_35/Y vdd CLKBUF1
XCLKBUF1_79 BUFX4_10/Y gnd CLKBUF1_79/Y vdd CLKBUF1
XCLKBUF1_68 BUFX4_12/Y gnd CLKBUF1_68/Y vdd CLKBUF1
XFILL_23_7_0 gnd vdd FILL
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XFILL_6_8_0 gnd vdd FILL
XBUFX4_407 INVX8_12/Y gnd NOR2X1_41/B vdd BUFX4
XBUFX4_418 INVX8_3/Y gnd BUFX4_418/Y vdd BUFX4
XBUFX4_429 d[7] gnd INVX8_9/A vdd BUFX4
XFILL_14_7_0 gnd vdd FILL
XOAI21X1_1308 INVX1_190/Y NOR2X1_264/Y NAND2X1_769/Y gnd DFFPOSX1_4/D vdd OAI21X1
XOAI21X1_1319 INVX1_383/Y NOR2X1_274/Y NAND2X1_781/Y gnd DFFPOSX1_39/D vdd OAI21X1
XDFFPOSX1_909 NAND2X1_538/B CLKBUF1_51/Y OAI21X1_700/Y gnd vdd DFFPOSX1
XOAI21X1_590 BUFX4_110/Y OAI21X1_590/B OAI21X1_590/C gnd OAI21X1_590/Y vdd OAI21X1
XFILL_39_1 gnd vdd FILL
XBUFX4_204 BUFX4_29/Y gnd BUFX4_204/Y vdd BUFX4
XBUFX4_237 BUFX4_31/Y gnd BUFX4_237/Y vdd BUFX4
XBUFX4_226 BUFX4_28/Y gnd BUFX4_226/Y vdd BUFX4
XBUFX4_215 BUFX4_23/Y gnd BUFX4_215/Y vdd BUFX4
XFILL_46_6_0 gnd vdd FILL
XBUFX4_248 BUFX4_28/Y gnd BUFX4_248/Y vdd BUFX4
XBUFX4_259 BUFX4_23/Y gnd BUFX4_259/Y vdd BUFX4
XNOR2X1_308 INVX4_2/Y OAI22X1_3/A gnd INVX8_14/A vdd NOR2X1
XNOR2X1_319 NOR2X1_319/A NOR2X1_315/B gnd NOR2X1_319/Y vdd NOR2X1
XOAI21X1_1116 INVX1_328/Y BUFX4_222/Y NAND2X1_559/Y gnd MUX2X1_242/A vdd OAI21X1
XOAI21X1_1127 INVX1_339/Y BUFX4_244/Y NAND2X1_571/Y gnd MUX2X1_251/B vdd OAI21X1
XOAI21X1_1105 INVX1_317/Y BUFX4_200/Y NAND2X1_548/Y gnd MUX2X1_235/B vdd OAI21X1
XOAI21X1_1138 INVX1_350/Y BUFX4_266/Y NAND2X1_583/Y gnd MUX2X1_259/A vdd OAI21X1
XDFFPOSX1_739 INVX1_171/A CLKBUF1_49/Y OAI21X1_555/Y gnd vdd DFFPOSX1
XDFFPOSX1_717 NAND2X1_525/B CLKBUF1_77/Y OAI21X1_538/Y gnd vdd DFFPOSX1
XDFFPOSX1_728 INVX1_490/A CLKBUF1_92/Y OAI21X1_552/Y gnd vdd DFFPOSX1
XOAI21X1_1149 INVX1_361/Y BUFX4_189/Y NAND2X1_594/Y gnd MUX2X1_268/B vdd OAI21X1
XDFFPOSX1_706 INVX1_105/A CLKBUF1_46/Y OAI21X1_516/Y gnd vdd DFFPOSX1
XINVX1_440 INVX1_440/A gnd INVX1_440/Y vdd INVX1
XINVX1_451 INVX1_451/A gnd INVX1_451/Y vdd INVX1
XINVX1_462 INVX1_462/A gnd INVX1_462/Y vdd INVX1
XINVX1_484 INVX1_484/A gnd INVX1_484/Y vdd INVX1
XINVX1_473 INVX1_473/A gnd INVX1_473/Y vdd INVX1
XINVX1_495 INVX1_495/A gnd INVX1_495/Y vdd INVX1
XNAND2X1_809 INVX8_9/A NOR2X1_309/Y gnd NAND2X1_809/Y vdd NAND2X1
XFILL_37_6_0 gnd vdd FILL
XFILL_20_5_0 gnd vdd FILL
XOAI21X1_1650 BUFX4_412/Y BUFX4_344/Y OAI21X1_802/B gnd OAI21X1_1650/Y vdd OAI21X1
XOAI21X1_1683 BUFX4_401/Y NAND2X1_871/Y OAI21X1_1683/C gnd DFFPOSX1_341/D vdd OAI21X1
XOAI21X1_1672 INVX1_401/Y NOR2X1_378/Y NAND2X1_869/Y gnd DFFPOSX1_327/D vdd OAI21X1
XOAI21X1_1661 BUFX4_97/Y NAND2X1_861/Y OAI21X1_1660/Y gnd DFFPOSX1_318/D vdd OAI21X1
XOAI21X1_1694 BUFX4_83/Y INVX2_11/A NAND2X1_363/B gnd OAI21X1_1694/Y vdd OAI21X1
XFILL_3_6_0 gnd vdd FILL
XNOR2X1_15 NOR2X1_15/A NOR2X1_14/B gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_26 NOR2X1_26/A NOR2X1_27/B gnd NOR2X1_26/Y vdd NOR2X1
XNOR2X1_37 NOR2X1_37/A NOR2X1_38/B gnd NOR2X1_37/Y vdd NOR2X1
XFILL_28_6_0 gnd vdd FILL
XNOR2X1_59 NOR2X1_59/A NOR2X1_55/B gnd NOR2X1_59/Y vdd NOR2X1
XNOR2X1_48 NOR2X1_48/A NOR2X1_43/B gnd NOR2X1_48/Y vdd NOR2X1
XFILL_11_5_0 gnd vdd FILL
XFILL_19_6_0 gnd vdd FILL
XMUX2X1_11 MUX2X1_11/A MUX2X1_11/B MUX2X1_11/S gnd MUX2X1_11/Y vdd MUX2X1
XMUX2X1_44 MUX2X1_44/A MUX2X1_44/B BUFX4_81/Y gnd MUX2X1_45/A vdd MUX2X1
XMUX2X1_22 MUX2X1_22/A MUX2X1_22/B BUFX4_192/Y gnd MUX2X1_24/B vdd MUX2X1
XNOR2X1_105 NOR2X1_105/A NOR2X1_103/B gnd NOR2X1_105/Y vdd NOR2X1
XMUX2X1_33 MUX2X1_33/A MUX2X1_33/B MUX2X1_7/S gnd AOI22X1_7/A vdd MUX2X1
XNOR2X1_149 NOR2X1_149/A NOR2X1_153/B gnd NOR2X1_149/Y vdd NOR2X1
XNOR2X1_138 NOR2X1_138/A NOR2X1_139/B gnd NOR2X1_138/Y vdd NOR2X1
XMUX2X1_88 MUX2X1_88/A MUX2X1_88/B BUFX4_80/Y gnd MUX2X1_88/Y vdd MUX2X1
XMUX2X1_66 MUX2X1_66/A MUX2X1_64/Y MUX2X1_7/S gnd MUX2X1_66/Y vdd MUX2X1
XMUX2X1_55 MUX2X1_55/A MUX2X1_55/B BUFX4_50/Y gnd MUX2X1_57/B vdd MUX2X1
XMUX2X1_77 MUX2X1_77/A MUX2X1_77/B BUFX4_51/Y gnd MUX2X1_78/A vdd MUX2X1
XNOR2X1_127 NOR2X1_127/A NOR2X1_126/B gnd NOR2X1_127/Y vdd NOR2X1
XNOR2X1_116 NOR2X1_116/A NOR2X1_118/B gnd NOR2X1_116/Y vdd NOR2X1
XMUX2X1_99 MUX2X1_99/A MUX2X1_99/B MUX2X1_7/S gnd MUX2X1_99/Y vdd MUX2X1
XDFFPOSX1_514 INVX1_93/A CLKBUF1_19/Y OAI21X1_228/Y gnd vdd DFFPOSX1
XDFFPOSX1_503 INVX1_412/A CLKBUF1_37/Y OAI21X1_223/Y gnd vdd DFFPOSX1
XDFFPOSX1_547 INVX1_159/A CLKBUF1_91/Y OAI21X1_267/Y gnd vdd DFFPOSX1
XDFFPOSX1_525 NAND2X1_513/B CLKBUF1_91/Y OAI21X1_250/Y gnd vdd DFFPOSX1
XDFFPOSX1_536 INVX1_478/A CLKBUF1_82/Y OAI21X1_264/Y gnd vdd DFFPOSX1
XDFFPOSX1_569 NAND2X1_258/B CLKBUF1_57/Y OAI21X1_290/Y gnd vdd DFFPOSX1
XINVX1_270 INVX1_270/A gnd INVX1_270/Y vdd INVX1
XDFFPOSX1_558 NOR2X1_58/A CLKBUF1_46/Y AOI21X1_46/Y gnd vdd DFFPOSX1
XINVX1_292 INVX1_292/A gnd INVX1_292/Y vdd INVX1
XNAND2X1_617 BUFX4_228/Y NOR2X1_262/A gnd NAND2X1_617/Y vdd NAND2X1
XINVX1_281 INVX1_281/A gnd INVX1_281/Y vdd INVX1
XNAND2X1_606 BUFX4_210/Y NOR2X1_174/A gnd NAND2X1_606/Y vdd NAND2X1
XNAND2X1_628 BUFX4_250/Y NAND2X1_628/B gnd NAND2X1_628/Y vdd NAND2X1
XNAND2X1_639 BUFX4_270/Y NAND2X1_639/B gnd NAND2X1_639/Y vdd NAND2X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XNAND2X1_70 BUFX4_450/Y NOR2X1_61/Y gnd NAND2X1_70/Y vdd NAND2X1
XNAND2X1_81 INVX2_3/Y INVX4_3/Y gnd NAND2X1_81/Y vdd NAND2X1
XNAND2X1_92 INVX2_4/Y INVX8_12/A gnd NAND2X1_92/Y vdd NAND2X1
XAOI21X1_241 BUFX4_112/Y NOR2X1_303/B NOR2X1_302/Y gnd AOI21X1_241/Y vdd AOI21X1
XAOI21X1_230 BUFX4_376/Y NOR2X1_279/B NOR2X1_283/Y gnd AOI21X1_230/Y vdd AOI21X1
XAOI21X1_252 BUFX4_97/Y NOR2X1_315/B NOR2X1_317/Y gnd AOI21X1_252/Y vdd AOI21X1
XAOI21X1_274 BUFX4_301/Y NOR2X1_342/B NOR2X1_345/Y gnd AOI21X1_274/Y vdd AOI21X1
XAOI21X1_285 BUFX4_380/Y NOR2X1_352/B NOR2X1_357/Y gnd AOI21X1_285/Y vdd AOI21X1
XAOI21X1_263 AOI21X1_1/A NOR2X1_338/B NOR2X1_333/Y gnd AOI21X1_263/Y vdd AOI21X1
XAOI21X1_296 BUFX4_114/Y NOR2X1_373/B NOR2X1_372/Y gnd AOI21X1_296/Y vdd AOI21X1
XOAI21X1_1480 BUFX4_305/Y NAND2X1_833/Y OAI21X1_1480/C gnd OAI21X1_1480/Y vdd OAI21X1
XOAI21X1_1491 NOR2X1_61/B BUFX4_94/Y INVX1_73/A gnd OAI21X1_1491/Y vdd OAI21X1
XFILL_43_4_0 gnd vdd FILL
XDFFPOSX1_1010 INVX1_124/A CLKBUF1_59/Y OAI21X1_792/Y gnd vdd DFFPOSX1
XDFFPOSX1_1021 NOR2X1_235/A CLKBUF1_22/Y AOI21X1_191/Y gnd vdd DFFPOSX1
XDFFPOSX1_1032 BUFX2_8/A CLKBUF1_65/Y NAND2X1_754/Y gnd vdd DFFPOSX1
XFILL_34_4_0 gnd vdd FILL
XOAI21X1_408 BUFX4_377/Y NAND2X1_82/Y OAI21X1_408/C gnd OAI21X1_408/Y vdd OAI21X1
XOAI21X1_419 BUFX4_403/Y BUFX4_337/Y INVX1_102/A gnd OAI21X1_420/C vdd OAI21X1
XDFFPOSX1_311 INVX1_400/A CLKBUF1_32/Y DFFPOSX1_311/D gnd vdd DFFPOSX1
XDFFPOSX1_322 INVX1_81/A CLKBUF1_97/Y OAI21X1_1667/Y gnd vdd DFFPOSX1
XDFFPOSX1_300 NOR2X1_373/A CLKBUF1_43/Y AOI21X1_297/Y gnd vdd DFFPOSX1
XDFFPOSX1_333 NOR2X1_384/A CLKBUF1_47/Y AOI21X1_306/Y gnd vdd DFFPOSX1
XDFFPOSX1_355 INVX1_147/A CLKBUF1_16/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_344 INVX1_466/A CLKBUF1_45/Y DFFPOSX1_344/D gnd vdd DFFPOSX1
XDFFPOSX1_377 OAI21X1_49/C CLKBUF1_22/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_366 OAI21X1_27/C CLKBUF1_28/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_388 INVX1_213/A CLKBUF1_33/Y OAI21X1_68/Y gnd vdd DFFPOSX1
XNAND2X1_414 BUFX4_248/Y DFFPOSX1_76/Q gnd OAI21X1_981/C vdd NAND2X1
XNAND2X1_403 BUFX4_230/Y NOR2X1_204/A gnd NAND2X1_403/Y vdd NAND2X1
XNAND2X1_425 BUFX4_270/Y NAND2X1_425/B gnd OAI21X1_992/C vdd NAND2X1
XNAND2X1_436 BUFX4_191/Y OAI21X1_95/C gnd NAND2X1_436/Y vdd NAND2X1
XDFFPOSX1_399 NOR2X1_9/A CLKBUF1_89/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XNAND2X1_469 BUFX4_253/Y NAND2X1_469/B gnd NAND2X1_469/Y vdd NAND2X1
XNAND2X1_458 BUFX4_233/Y NOR2X1_96/A gnd NAND2X1_458/Y vdd NAND2X1
XNAND2X1_447 BUFX4_211/Y NAND2X1_447/B gnd NAND2X1_447/Y vdd NAND2X1
XFILL_0_4_0 gnd vdd FILL
XFILL_25_4_0 gnd vdd FILL
XOAI21X1_942 INVX1_154/Y BUFX4_270/Y NAND2X1_371/Y gnd MUX2X1_112/A vdd OAI21X1
XOAI21X1_931 INVX1_143/Y BUFX4_248/Y NAND2X1_360/Y gnd MUX2X1_104/B vdd OAI21X1
XOAI21X1_920 INVX1_132/Y BUFX4_226/Y NAND2X1_348/Y gnd MUX2X1_95/A vdd OAI21X1
XOAI21X1_964 INVX1_176/Y BUFX4_215/Y NAND2X1_395/Y gnd MUX2X1_128/A vdd OAI21X1
XOAI21X1_975 INVX1_187/Y BUFX4_237/Y OAI21X1_975/C gnd MUX2X1_137/B vdd OAI21X1
XOAI21X1_953 INVX1_165/Y BUFX4_193/Y NAND2X1_383/Y gnd MUX2X1_121/B vdd OAI21X1
XOAI21X1_997 INVX1_209/Y MUX2X1_4/S OAI21X1_997/C gnd MUX2X1_154/B vdd OAI21X1
XOAI21X1_986 INVX1_198/Y BUFX4_259/Y OAI21X1_986/C gnd MUX2X1_145/A vdd OAI21X1
XFILL_8_5_0 gnd vdd FILL
XFILL_16_4_0 gnd vdd FILL
XOAI21X1_13 BUFX4_312/Y BUFX4_317/Y INVX1_403/A gnd OAI21X1_14/C vdd OAI21X1
XOAI21X1_24 BUFX4_300/Y NAND2X1_2/Y OAI21X1_23/Y gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_35 BUFX4_171/Y BUFX4_317/Y INVX1_84/A gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_46 NAND2X1_3/Y BUFX4_283/Y OAI21X1_46/C gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_57 BUFX4_415/Y BUFX4_314/Y OAI21X1_57/C gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_68 INVX1_213/Y NOR2X1_1/Y NAND2X1_9/Y gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_79 NOR2X1_81/B NOR2X1_1/A INVX1_214/A gnd OAI21X1_80/C vdd OAI21X1
XOAI21X1_238 BUFX4_287/Y NAND2X1_48/Y OAI21X1_237/Y gnd OAI21X1_238/Y vdd OAI21X1
XOAI21X1_227 BUFX4_461/Y BUFX4_437/Y INVX1_93/A gnd OAI21X1_227/Y vdd OAI21X1
XOAI21X1_205 INVX1_282/Y NOR2X1_11/Y NAND2X1_27/Y gnd OAI21X1_205/Y vdd OAI21X1
XOAI21X1_216 INVX1_475/Y NOR2X1_21/Y NAND2X1_38/Y gnd OAI21X1_216/Y vdd OAI21X1
XOAI21X1_249 BUFX4_150/Y BUFX4_437/Y NAND2X1_513/B gnd OAI21X1_249/Y vdd OAI21X1
XDFFPOSX1_130 INVX1_69/A CLKBUF1_98/Y OAI21X1_1412/Y gnd vdd DFFPOSX1
XDFFPOSX1_163 INVX1_135/A CLKBUF1_63/Y OAI21X1_1451/Y gnd vdd DFFPOSX1
XDFFPOSX1_152 INVX1_454/A CLKBUF1_68/Y OAI21X1_1448/Y gnd vdd DFFPOSX1
XDFFPOSX1_141 NAND2X1_487/B CLKBUF1_68/Y OAI21X1_1434/Y gnd vdd DFFPOSX1
XDFFPOSX1_196 INVX1_201/A CLKBUF1_51/Y DFFPOSX1_196/D gnd vdd DFFPOSX1
XNAND2X1_211 NAND2X1_211/A INVX1_509/A gnd OAI21X1_800/C vdd NAND2X1
XNAND2X1_200 INVX2_5/Y INVX8_12/A gnd OAI21X1_761/B vdd NAND2X1
XDFFPOSX1_174 NOR2X1_338/A CLKBUF1_68/Y AOI21X1_268/Y gnd vdd DFFPOSX1
XDFFPOSX1_185 NAND2X1_253/B CLKBUF1_84/Y OAI21X1_1474/Y gnd vdd DFFPOSX1
XNAND2X1_233 BUFX4_227/Y NOR2X1_266/A gnd NAND2X1_233/Y vdd NAND2X1
XNAND2X1_222 BUFX4_213/Y OAI21X1_121/C gnd OAI21X1_811/C vdd NAND2X1
XNAND2X1_244 INVX4_1/Y NAND2X1_244/B gnd AOI21X1_204/A vdd NAND2X1
XNAND2X1_255 BUFX4_249/Y OAI21X1_241/C gnd OAI21X1_833/C vdd NAND2X1
XNAND2X1_266 BUFX4_271/Y OAI21X1_497/C gnd NAND2X1_266/Y vdd NAND2X1
XNAND2X1_277 BUFX4_192/Y NOR2X1_301/A gnd OAI21X1_854/C vdd NAND2X1
XNAND2X1_288 AOI22X1_10/Y AOI22X1_11/Y gnd AOI22X1_14/A vdd NAND2X1
XNAND2X1_299 BUFX4_234/Y NAND2X1_299/B gnd OAI21X1_875/C vdd NAND2X1
XFILL_41_7_1 gnd vdd FILL
XFILL_40_2_0 gnd vdd FILL
XOAI21X1_750 NOR2X1_72/B BUFX4_443/Y NAND2X1_473/B gnd OAI21X1_751/C vdd OAI21X1
XOAI21X1_783 BUFX4_302/Y NAND2X1_201/Y OAI21X1_782/Y gnd OAI21X1_783/Y vdd OAI21X1
XOAI21X1_794 INVX1_252/Y NOR2X1_228/Y OAI21X1_794/C gnd OAI21X1_794/Y vdd OAI21X1
XOAI21X1_772 BUFX4_409/Y INVX2_5/A INVX1_442/A gnd OAI21X1_773/C vdd OAI21X1
XOAI21X1_761 BUFX4_130/Y OAI21X1_761/B OAI21X1_761/C gnd OAI21X1_761/Y vdd OAI21X1
XMUX2X1_250 MUX2X1_250/A MUX2X1_250/B BUFX4_43/Y gnd MUX2X1_250/Y vdd MUX2X1
XMUX2X1_283 MUX2X1_283/A MUX2X1_283/B BUFX4_32/Y gnd MUX2X1_285/B vdd MUX2X1
XMUX2X1_272 MUX2X1_272/A MUX2X1_272/B MUX2X1_3/S gnd MUX2X1_272/Y vdd MUX2X1
XMUX2X1_261 MUX2X1_261/A MUX2X1_261/B MUX2X1_96/S gnd AOI22X1_55/A vdd MUX2X1
XMUX2X1_294 MUX2X1_293/Y MUX2X1_292/Y MUX2X1_96/S gnd MUX2X1_294/Y vdd MUX2X1
XFILL_48_3_0 gnd vdd FILL
XFILL_32_7_1 gnd vdd FILL
XFILL_31_2_0 gnd vdd FILL
XCLKBUF1_14 BUFX4_16/Y gnd CLKBUF1_14/Y vdd CLKBUF1
XCLKBUF1_47 BUFX4_10/Y gnd CLKBUF1_47/Y vdd CLKBUF1
XCLKBUF1_36 BUFX4_17/Y gnd CLKBUF1_36/Y vdd CLKBUF1
XCLKBUF1_25 BUFX4_12/Y gnd CLKBUF1_25/Y vdd CLKBUF1
XCLKBUF1_69 BUFX4_15/Y gnd CLKBUF1_69/Y vdd CLKBUF1
XCLKBUF1_58 BUFX4_15/Y gnd CLKBUF1_58/Y vdd CLKBUF1
XFILL_39_3_0 gnd vdd FILL
XBUFX4_90 BUFX4_92/A gnd INVX2_9/A vdd BUFX4
XFILL_23_7_1 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XFILL_6_8_1 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XBUFX4_419 INVX8_3/Y gnd BUFX4_419/Y vdd BUFX4
XBUFX4_408 INVX8_12/Y gnd NOR2X1_81/B vdd BUFX4
XFILL_14_7_1 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XOAI21X1_1309 INVX1_254/Y NOR2X1_264/Y NAND2X1_770/Y gnd DFFPOSX1_5/D vdd OAI21X1
XOAI21X1_580 BUFX4_104/Y OAI21X1_584/B OAI21X1_580/C gnd OAI21X1_580/Y vdd OAI21X1
XOAI21X1_591 BUFX4_148/Y BUFX4_105/Y NAND2X1_461/B gnd OAI21X1_592/C vdd OAI21X1
XBUFX4_227 BUFX4_24/Y gnd BUFX4_227/Y vdd BUFX4
XBUFX4_205 BUFX4_26/Y gnd BUFX4_205/Y vdd BUFX4
XBUFX4_216 BUFX4_27/Y gnd BUFX4_216/Y vdd BUFX4
XFILL_46_6_1 gnd vdd FILL
XBUFX4_238 BUFX4_23/Y gnd BUFX4_238/Y vdd BUFX4
XBUFX4_249 BUFX4_25/Y gnd BUFX4_249/Y vdd BUFX4
XFILL_45_1_0 gnd vdd FILL
XNOR2X1_309 BUFX4_466/Y NOR2X1_51/B gnd NOR2X1_309/Y vdd NOR2X1
XOAI21X1_1128 INVX1_340/Y BUFX4_246/Y NAND2X1_572/Y gnd MUX2X1_251/A vdd OAI21X1
XOAI21X1_1106 INVX1_318/Y BUFX4_202/Y NAND2X1_549/Y gnd MUX2X1_235/A vdd OAI21X1
XOAI21X1_1117 INVX1_329/Y BUFX4_224/Y NAND2X1_560/Y gnd MUX2X1_244/B vdd OAI21X1
XDFFPOSX1_707 INVX1_169/A CLKBUF1_82/Y OAI21X1_518/Y gnd vdd DFFPOSX1
XDFFPOSX1_718 NAND2X1_594/B CLKBUF1_82/Y OAI21X1_540/Y gnd vdd DFFPOSX1
XDFFPOSX1_729 NOR2X1_83/A CLKBUF1_41/Y AOI21X1_65/Y gnd vdd DFFPOSX1
XOAI21X1_1139 INVX1_351/Y BUFX4_268/Y NAND2X1_584/Y gnd MUX2X1_260/B vdd OAI21X1
XINVX1_441 INVX1_441/A gnd INVX1_441/Y vdd INVX1
XINVX1_430 INVX1_430/A gnd INVX1_430/Y vdd INVX1
XINVX1_452 INVX1_452/A gnd INVX1_452/Y vdd INVX1
XINVX1_474 INVX1_474/A gnd INVX1_474/Y vdd INVX1
XINVX1_485 INVX1_485/A gnd INVX1_485/Y vdd INVX1
XINVX1_496 INVX1_496/A gnd INVX1_496/Y vdd INVX1
XINVX1_463 INVX1_463/A gnd INVX1_463/Y vdd INVX1
XFILL_37_6_1 gnd vdd FILL
XFILL_36_1_0 gnd vdd FILL
XFILL_20_5_1 gnd vdd FILL
XOAI21X1_1640 BUFX4_168/Y BUFX4_343/Y INVX1_208/A gnd OAI21X1_1640/Y vdd OAI21X1
XOAI21X1_1651 BUFX4_129/Y NAND2X1_861/Y OAI21X1_1650/Y gnd DFFPOSX1_313/D vdd OAI21X1
XOAI21X1_1662 BUFX4_412/Y BUFX4_344/Y NAND2X1_637/B gnd OAI21X1_1662/Y vdd OAI21X1
XOAI21X1_1684 BUFX4_406/Y OAI21X1_5/B INVX1_338/A gnd OAI21X1_1685/C vdd OAI21X1
XOAI21X1_1673 INVX1_465/Y NOR2X1_378/Y NAND2X1_870/Y gnd DFFPOSX1_328/D vdd OAI21X1
XOAI21X1_1695 BUFX4_109/Y NAND2X1_872/Y OAI21X1_1694/Y gnd DFFPOSX1_347/D vdd OAI21X1
XNOR2X1_16 NOR2X1_16/A NOR2X1_14/B gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_27 NOR2X1_27/A NOR2X1_27/B gnd NOR2X1_27/Y vdd NOR2X1
XFILL_28_6_1 gnd vdd FILL
XNOR2X1_49 NOR2X1_49/A NOR2X1_43/B gnd NOR2X1_49/Y vdd NOR2X1
XFILL_3_6_1 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B gnd NOR2X1_38/Y vdd NOR2X1
XFILL_27_1_0 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XFILL_10_0_0 gnd vdd FILL
XFILL_19_6_1 gnd vdd FILL
XMUX2X1_34 MUX2X1_34/A MUX2X1_34/B BUFX4_2/Y gnd MUX2X1_36/B vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XMUX2X1_45 MUX2X1_45/A MUX2X1_43/Y INVX2_6/A gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_23 MUX2X1_23/A MUX2X1_23/B BUFX4_193/Y gnd MUX2X1_24/A vdd MUX2X1
XNOR2X1_106 NOR2X1_106/A NOR2X1_103/B gnd AOI21X1_84/C vdd NOR2X1
XMUX2X1_12 MUX2X1_12/A MUX2X1_12/B MUX2X1_12/S gnd MUX2X1_13/A vdd MUX2X1
XMUX2X1_67 MUX2X1_67/A MUX2X1_67/B BUFX4_81/Y gnd MUX2X1_69/B vdd MUX2X1
XNOR2X1_139 NOR2X1_139/A NOR2X1_139/B gnd NOR2X1_139/Y vdd NOR2X1
XMUX2X1_78 MUX2X1_78/A MUX2X1_76/Y INVX2_6/A gnd MUX2X1_78/Y vdd MUX2X1
XNOR2X1_128 NOR2X1_128/A NOR2X1_126/B gnd NOR2X1_128/Y vdd NOR2X1
XMUX2X1_56 MUX2X1_56/A MUX2X1_56/B BUFX4_3/Y gnd MUX2X1_57/A vdd MUX2X1
XNOR2X1_117 NOR2X1_117/A NOR2X1_118/B gnd AOI21X1_93/C vdd NOR2X1
XMUX2X1_89 MUX2X1_89/A MUX2X1_89/B BUFX4_81/Y gnd MUX2X1_89/Y vdd MUX2X1
XDFFPOSX1_504 INVX1_476/A CLKBUF1_31/Y OAI21X1_224/Y gnd vdd DFFPOSX1
XDFFPOSX1_515 INVX1_157/A CLKBUF1_1/Y OAI21X1_230/Y gnd vdd DFFPOSX1
XDFFPOSX1_537 NOR2X1_43/A CLKBUF1_1/Y AOI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_526 OAI21X1_251/C CLKBUF1_19/Y OAI21X1_252/Y gnd vdd DFFPOSX1
XINVX1_260 INVX1_260/A gnd INVX1_260/Y vdd INVX1
XDFFPOSX1_548 INVX1_223/A CLKBUF1_46/Y OAI21X1_268/Y gnd vdd DFFPOSX1
XINVX1_271 INVX1_271/A gnd INVX1_271/Y vdd INVX1
XDFFPOSX1_559 NOR2X1_59/A CLKBUF1_27/Y AOI21X1_47/Y gnd vdd DFFPOSX1
XNAND2X1_607 BUFX4_212/Y NAND2X1_607/B gnd NAND2X1_607/Y vdd NAND2X1
XINVX1_282 INVX1_282/A gnd INVX1_282/Y vdd INVX1
XNAND2X1_618 BUFX4_230/Y NOR2X1_272/A gnd NAND2X1_618/Y vdd NAND2X1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XNAND2X1_629 BUFX4_252/Y NAND2X1_629/B gnd NAND2X1_629/Y vdd NAND2X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_60 NAND2X1_8/A NOR2X1_51/Y gnd NAND2X1_60/Y vdd NAND2X1
XNAND2X1_82 INVX8_16/A INVX2_3/Y gnd NAND2X1_82/Y vdd NAND2X1
XNAND2X1_93 INVX2_4/Y INVX8_13/A gnd NAND2X1_93/Y vdd NAND2X1
XNAND2X1_71 BUFX4_332/Y NOR2X1_61/Y gnd NAND2X1_71/Y vdd NAND2X1
XAOI21X1_242 BUFX4_305/Y NOR2X1_303/B NOR2X1_303/Y gnd AOI21X1_242/Y vdd AOI21X1
XAOI21X1_220 BUFX4_98/Y NOR2X1_265/Y NOR2X1_271/Y gnd AOI21X1_220/Y vdd AOI21X1
XAOI21X1_231 AOI21X1_1/A NOR2X1_289/B NOR2X1_286/Y gnd AOI21X1_231/Y vdd AOI21X1
XAOI21X1_275 BUFX4_402/Y NOR2X1_342/B NOR2X1_346/Y gnd AOI21X1_275/Y vdd AOI21X1
XAOI21X1_264 BUFX4_423/Y NOR2X1_338/B NOR2X1_334/Y gnd AOI21X1_264/Y vdd AOI21X1
XAOI21X1_253 BUFX4_280/Y NOR2X1_315/B NOR2X1_318/Y gnd AOI21X1_253/Y vdd AOI21X1
XAOI21X1_286 AOI21X1_1/A NOR2X1_367/B NOR2X1_360/Y gnd AOI21X1_286/Y vdd AOI21X1
XAOI21X1_297 BUFX4_305/Y NOR2X1_373/B NOR2X1_373/Y gnd AOI21X1_297/Y vdd AOI21X1
XOAI21X1_1470 NAND2X1_832/Y BUFX4_286/Y OAI21X1_1469/Y gnd OAI21X1_1470/Y vdd OAI21X1
XOAI21X1_1492 BUFX4_426/Y NAND2X1_834/Y OAI21X1_1491/Y gnd DFFPOSX1_194/D vdd OAI21X1
XOAI21X1_1481 BUFX4_417/Y INVX2_8/A NAND2X1_490/B gnd OAI21X1_1481/Y vdd OAI21X1
XFILL_43_4_1 gnd vdd FILL
XDFFPOSX1_1000 INVX1_507/A CLKBUF1_73/Y OAI21X1_791/Y gnd vdd DFFPOSX1
XDFFPOSX1_1011 INVX1_188/A CLKBUF1_40/Y OAI21X1_793/Y gnd vdd DFFPOSX1
XDFFPOSX1_1022 NOR2X1_236/A CLKBUF1_40/Y AOI21X1_192/Y gnd vdd DFFPOSX1
XFILL_34_4_1 gnd vdd FILL
XFILL_14_1 gnd vdd FILL
XOAI21X1_409 INVX1_53/Y NOR2X1_71/Y NAND2X1_84/Y gnd OAI21X1_409/Y vdd OAI21X1
XDFFPOSX1_312 INVX1_464/A CLKBUF1_32/Y DFFPOSX1_312/D gnd vdd DFFPOSX1
XDFFPOSX1_301 NOR2X1_374/A CLKBUF1_12/Y AOI21X1_298/Y gnd vdd DFFPOSX1
XDFFPOSX1_345 NAND2X1_220/B CLKBUF1_38/Y DFFPOSX1_345/D gnd vdd DFFPOSX1
XDFFPOSX1_356 INVX1_211/A CLKBUF1_34/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_334 NOR2X1_385/A CLKBUF1_97/Y AOI21X1_307/Y gnd vdd DFFPOSX1
XDFFPOSX1_323 INVX1_145/A CLKBUF1_85/Y OAI21X1_1668/Y gnd vdd DFFPOSX1
XDFFPOSX1_367 OAI21X1_29/C CLKBUF1_8/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_378 OAI21X1_51/C CLKBUF1_8/Y OAI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_389 INVX1_277/A CLKBUF1_12/Y OAI21X1_69/Y gnd vdd DFFPOSX1
XNAND2X1_415 BUFX4_250/Y NOR2X1_303/A gnd OAI21X1_982/C vdd NAND2X1
XNAND2X1_404 BUFX4_232/Y NAND2X1_404/B gnd OAI21X1_973/C vdd NAND2X1
XNAND2X1_426 AOI22X1_30/Y AOI22X1_31/Y gnd AOI22X1_34/A vdd NAND2X1
XNAND2X1_448 BUFX4_213/Y NOR2X1_66/A gnd NAND2X1_448/Y vdd NAND2X1
XNAND2X1_459 BUFX4_235/Y NOR2X1_106/A gnd NAND2X1_459/Y vdd NAND2X1
XNAND2X1_437 BUFX4_193/Y OAI21X1_127/C gnd NAND2X1_437/Y vdd NAND2X1
XFILL_0_4_1 gnd vdd FILL
XFILL_25_4_1 gnd vdd FILL
XOAI21X1_932 INVX1_144/Y BUFX4_250/Y NAND2X1_361/Y gnd MUX2X1_104/A vdd OAI21X1
XOAI21X1_910 INVX1_122/Y BUFX4_206/Y OAI21X1_910/C gnd MUX2X1_88/A vdd OAI21X1
XOAI21X1_943 INVX1_155/Y BUFX4_272/Y OAI21X1_943/C gnd MUX2X1_113/B vdd OAI21X1
XOAI21X1_921 INVX1_133/Y BUFX4_228/Y NAND2X1_349/Y gnd MUX2X1_97/B vdd OAI21X1
XOAI21X1_954 INVX1_166/Y BUFX4_195/Y NAND2X1_384/Y gnd MUX2X1_121/A vdd OAI21X1
XOAI21X1_976 INVX1_188/Y BUFX4_239/Y NAND2X1_407/Y gnd MUX2X1_137/A vdd OAI21X1
XOAI21X1_965 INVX1_177/Y BUFX4_217/Y OAI21X1_965/C gnd MUX2X1_130/B vdd OAI21X1
XOAI21X1_998 INVX1_210/Y MUX2X1_8/S NAND2X1_432/Y gnd MUX2X1_154/A vdd OAI21X1
XOAI21X1_987 INVX1_199/Y BUFX4_261/Y OAI21X1_987/C gnd MUX2X1_146/B vdd OAI21X1
XFILL_8_5_1 gnd vdd FILL
XDFFPOSX1_890 NOR2X1_170/A CLKBUF1_13/Y AOI21X1_136/Y gnd vdd DFFPOSX1
XFILL_7_0_0 gnd vdd FILL
XFILL_16_4_1 gnd vdd FILL
XOAI21X1_14 BUFX4_283/Y NAND2X1_1/Y OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_25 BUFX4_368/Y BUFX4_319/Y OAI21X1_25/C gnd OAI21X1_26/C vdd OAI21X1
XOAI21X1_58 BUFX4_398/Y NAND2X1_4/Y OAI21X1_57/Y gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_47 BUFX4_171/Y OAI21X1_7/B INVX1_468/A gnd OAI21X1_48/C vdd OAI21X1
XOAI21X1_36 NAND2X1_3/Y BUFX4_424/Y OAI21X1_35/Y gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_69 INVX1_277/Y NOR2X1_1/Y NAND2X1_10/Y gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_228 BUFX4_422/Y NAND2X1_48/Y OAI21X1_227/Y gnd OAI21X1_228/Y vdd OAI21X1
XOAI21X1_206 INVX1_346/Y NOR2X1_11/Y NAND2X1_28/Y gnd OAI21X1_206/Y vdd OAI21X1
XOAI21X1_217 INVX1_29/Y NOR2X1_31/Y NAND2X1_39/Y gnd OAI21X1_217/Y vdd OAI21X1
XOAI21X1_239 BUFX4_461/Y BUFX4_434/Y INVX1_477/A gnd OAI21X1_239/Y vdd OAI21X1
XDFFPOSX1_120 INVX1_452/A CLKBUF1_17/Y DFFPOSX1_120/D gnd vdd DFFPOSX1
XDFFPOSX1_142 NAND2X1_556/B CLKBUF1_63/Y OAI21X1_1436/Y gnd vdd DFFPOSX1
XDFFPOSX1_164 INVX1_199/A CLKBUF1_98/Y OAI21X1_1452/Y gnd vdd DFFPOSX1
XDFFPOSX1_153 NOR2X1_323/A CLKBUF1_98/Y AOI21X1_255/Y gnd vdd DFFPOSX1
XDFFPOSX1_131 INVX1_133/A CLKBUF1_102/Y DFFPOSX1_131/D gnd vdd DFFPOSX1
XDFFPOSX1_186 NAND2X1_283/B CLKBUF1_43/Y OAI21X1_1476/Y gnd vdd DFFPOSX1
XDFFPOSX1_197 INVX1_265/A CLKBUF1_36/Y OAI21X1_1498/Y gnd vdd DFFPOSX1
XNAND2X1_201 INVX2_5/Y INVX8_14/A gnd NAND2X1_201/Y vdd NAND2X1
XDFFPOSX1_175 NOR2X1_339/A CLKBUF1_68/Y AOI21X1_269/Y gnd vdd DFFPOSX1
XNAND2X1_212 INVX8_1/Y NOR2X1_244/Y gnd OAI22X1_3/A vdd NAND2X1
XNAND2X1_234 BUFX4_81/Y OAI21X1_819/Y gnd AOI21X1_201/B vdd NAND2X1
XNAND2X1_223 NOR2X1_244/Y NAND2X1_223/B gnd NAND3X1_3/B vdd NAND2X1
XNAND2X1_256 BUFX4_251/Y NOR2X1_43/A gnd OAI21X1_834/C vdd NAND2X1
XNAND2X1_278 BUFX4_194/Y NOR2X1_313/A gnd OAI21X1_855/C vdd NAND2X1
XNAND2X1_245 BUFX4_239/Y NAND2X1_245/B gnd OAI21X1_826/C vdd NAND2X1
XNAND2X1_267 BUFX4_273/Y NAND2X1_267/B gnd OAI21X1_845/C vdd NAND2X1
XNAND2X1_289 BUFX4_214/Y NAND2X1_289/B gnd OAI21X1_865/C vdd NAND2X1
XFILL_40_2_1 gnd vdd FILL
XOAI21X1_751 BUFX4_302/Y OAI21X1_757/B OAI21X1_751/C gnd OAI21X1_751/Y vdd OAI21X1
XOAI21X1_740 BUFX4_455/Y BUFX4_442/Y INVX1_441/A gnd OAI21X1_741/C vdd OAI21X1
XOAI21X1_784 BUFX4_308/Y BUFX4_438/Y INVX1_315/A gnd OAI21X1_785/C vdd OAI21X1
XOAI21X1_762 BUFX4_409/Y BUFX4_440/Y INVX1_122/A gnd OAI21X1_763/C vdd OAI21X1
XOAI21X1_773 BUFX4_281/Y OAI21X1_761/B OAI21X1_773/C gnd OAI21X1_773/Y vdd OAI21X1
XOAI21X1_795 INVX1_316/Y NOR2X1_228/Y OAI21X1_795/C gnd OAI21X1_795/Y vdd OAI21X1
XMUX2X1_240 MUX2X1_240/A MUX2X1_240/B MUX2X1_42/S gnd AOI22X1_50/D vdd MUX2X1
XMUX2X1_251 MUX2X1_251/A MUX2X1_251/B BUFX4_59/Y gnd MUX2X1_251/Y vdd MUX2X1
XMUX2X1_284 MUX2X1_284/A MUX2X1_284/B BUFX4_52/Y gnd MUX2X1_285/A vdd MUX2X1
XMUX2X1_262 MUX2X1_262/A MUX2X1_262/B BUFX4_55/Y gnd MUX2X1_262/Y vdd MUX2X1
XMUX2X1_273 MUX2X1_272/Y MUX2X1_273/B MUX2X1_42/S gnd AOI22X1_57/A vdd MUX2X1
XMUX2X1_295 MUX2X1_295/A MUX2X1_295/B BUFX4_41/Y gnd MUX2X1_297/B vdd MUX2X1
XFILL_48_3_1 gnd vdd FILL
XNAND2X1_790 BUFX4_427/Y NOR2X1_284/Y gnd NAND2X1_790/Y vdd NAND2X1
XFILL_31_2_1 gnd vdd FILL
XCLKBUF1_15 BUFX4_18/Y gnd CLKBUF1_15/Y vdd CLKBUF1
XCLKBUF1_37 BUFX4_11/Y gnd CLKBUF1_37/Y vdd CLKBUF1
XCLKBUF1_26 BUFX4_9/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XCLKBUF1_48 BUFX4_14/Y gnd CLKBUF1_48/Y vdd CLKBUF1
XCLKBUF1_59 BUFX4_15/Y gnd CLKBUF1_59/Y vdd CLKBUF1
XFILL_39_3_1 gnd vdd FILL
XBUFX4_80 a[1] gnd BUFX4_80/Y vdd BUFX4
XBUFX4_91 BUFX4_92/A gnd BUFX4_91/Y vdd BUFX4
XFILL_22_2_1 gnd vdd FILL
XFILL_5_3_1 gnd vdd FILL
XBUFX4_409 INVX8_12/Y gnd BUFX4_409/Y vdd BUFX4
XFILL_13_2_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XOAI21X1_581 BUFX4_455/Y BUFX4_108/Y INVX1_429/A gnd OAI21X1_582/C vdd OAI21X1
XOAI21X1_570 BUFX4_130/Y OAI21X1_584/B OAI21X1_570/C gnd OAI21X1_570/Y vdd OAI21X1
XOAI21X1_592 BUFX4_298/Y OAI21X1_590/B OAI21X1_592/C gnd OAI21X1_592/Y vdd OAI21X1
XBUFX4_217 BUFX4_31/Y gnd BUFX4_217/Y vdd BUFX4
XBUFX4_206 BUFX4_23/Y gnd BUFX4_206/Y vdd BUFX4
XBUFX4_228 BUFX4_27/Y gnd BUFX4_228/Y vdd BUFX4
XBUFX4_239 BUFX4_30/Y gnd BUFX4_239/Y vdd BUFX4
XFILL_45_1_1 gnd vdd FILL
XOAI21X1_1118 INVX1_330/Y BUFX4_226/Y NAND2X1_561/Y gnd MUX2X1_244/A vdd OAI21X1
XOAI21X1_1107 INVX1_319/Y BUFX4_204/Y NAND2X1_550/Y gnd MUX2X1_236/B vdd OAI21X1
XOAI21X1_1129 INVX1_341/Y BUFX4_248/Y NAND2X1_573/Y gnd MUX2X1_253/B vdd OAI21X1
XINVX1_420 INVX1_420/A gnd INVX1_420/Y vdd INVX1
XDFFPOSX1_719 OAI21X1_541/C CLKBUF1_29/Y OAI21X1_542/Y gnd vdd DFFPOSX1
XDFFPOSX1_708 INVX1_233/A CLKBUF1_54/Y OAI21X1_520/Y gnd vdd DFFPOSX1
XINVX1_442 INVX1_442/A gnd INVX1_442/Y vdd INVX1
XINVX1_431 INVX1_431/A gnd INVX1_431/Y vdd INVX1
XINVX1_453 INVX1_453/A gnd INVX1_453/Y vdd INVX1
XINVX1_486 INVX1_486/A gnd INVX1_486/Y vdd INVX1
XINVX1_475 INVX1_475/A gnd INVX1_475/Y vdd INVX1
XINVX1_464 INVX1_464/A gnd INVX1_464/Y vdd INVX1
XINVX1_497 INVX1_497/A gnd INVX1_497/Y vdd INVX1
XFILL_44_1 gnd vdd FILL
XFILL_36_1_1 gnd vdd FILL
XOAI21X1_1641 NAND2X1_860/Y BUFX4_305/Y OAI21X1_1640/Y gnd OAI21X1_1641/Y vdd OAI21X1
XOAI21X1_1630 INVX1_271/Y NOR2X1_368/Y NAND2X1_856/Y gnd OAI21X1_1630/Y vdd OAI21X1
XOAI21X1_1663 BUFX4_286/Y NAND2X1_861/Y OAI21X1_1662/Y gnd DFFPOSX1_319/D vdd OAI21X1
XOAI21X1_1674 BUFX4_406/Y INVX2_11/A INVX1_23/A gnd OAI21X1_1675/C vdd OAI21X1
XOAI21X1_1652 BUFX4_416/Y BUFX4_344/Y NAND2X1_292/B gnd OAI21X1_1652/Y vdd OAI21X1
XOAI21X1_1696 BUFX4_83/Y INVX2_11/A NAND2X1_432/B gnd OAI21X1_1697/C vdd OAI21X1
XOAI21X1_1685 BUFX4_101/Y NAND2X1_871/Y OAI21X1_1685/C gnd DFFPOSX1_342/D vdd OAI21X1
XNOR2X1_17 NOR2X1_17/A NOR2X1_14/B gnd NOR2X1_17/Y vdd NOR2X1
XNOR2X1_28 NOR2X1_28/A NOR2X1_27/B gnd NOR2X1_28/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XNOR2X1_39 NOR2X1_39/A NOR2X1_38/B gnd NOR2X1_39/Y vdd NOR2X1
XFILL_27_1_1 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XMUX2X1_35 MUX2X1_35/A MUX2X1_35/B BUFX4_33/Y gnd MUX2X1_35/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XMUX2X1_24 MUX2X1_24/A MUX2X1_24/B BUFX4_1/Y gnd MUX2X1_28/B vdd MUX2X1
XMUX2X1_13 MUX2X1_13/A MUX2X1_11/Y BUFX4_44/Y gnd MUX2X1_14/A vdd MUX2X1
XMUX2X1_68 MUX2X1_68/A MUX2X1_68/B BUFX4_82/Y gnd MUX2X1_69/A vdd MUX2X1
XNOR2X1_129 NOR2X1_129/A NOR2X1_126/B gnd NOR2X1_129/Y vdd NOR2X1
XMUX2X1_57 MUX2X1_57/A MUX2X1_57/B BUFX4_363/Y gnd MUX2X1_57/Y vdd MUX2X1
XNOR2X1_107 NOR2X1_107/A NOR2X1_103/B gnd AOI21X1_85/C vdd NOR2X1
XMUX2X1_79 MUX2X1_79/A MUX2X1_79/B BUFX4_4/Y gnd MUX2X1_81/B vdd MUX2X1
XMUX2X1_46 MUX2X1_46/A MUX2X1_46/B BUFX4_82/Y gnd MUX2X1_48/B vdd MUX2X1
XNOR2X1_118 NOR2X1_118/A NOR2X1_118/B gnd AOI21X1_94/C vdd NOR2X1
XFILL_30_8_0 gnd vdd FILL
XDFFPOSX1_505 NOR2X1_33/A CLKBUF1_56/Y AOI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_516 INVX1_221/A CLKBUF1_80/Y OAI21X1_232/Y gnd vdd DFFPOSX1
XDFFPOSX1_538 NOR2X1_44/A CLKBUF1_80/Y AOI21X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_527 NAND2X1_651/B CLKBUF1_41/Y OAI21X1_254/Y gnd vdd DFFPOSX1
XINVX1_250 INVX1_250/A gnd INVX1_250/Y vdd INVX1
XINVX1_261 INVX1_261/A gnd INVX1_261/Y vdd INVX1
XDFFPOSX1_549 INVX1_287/A CLKBUF1_11/Y OAI21X1_269/Y gnd vdd DFFPOSX1
XNAND2X1_608 BUFX4_214/Y NOR2X1_185/A gnd NAND2X1_608/Y vdd NAND2X1
XINVX1_294 INVX1_294/A gnd INVX1_294/Y vdd INVX1
XINVX1_283 INVX1_283/A gnd INVX1_283/Y vdd INVX1
XINVX1_272 INVX1_272/A gnd INVX1_272/Y vdd INVX1
XNAND2X1_619 BUFX4_232/Y NOR2X1_282/A gnd NAND2X1_619/Y vdd NAND2X1
XNAND2X1_50 INVX8_2/A NOR2X1_41/Y gnd NAND2X1_50/Y vdd NAND2X1
XNAND2X1_61 NAND2X1_9/A NOR2X1_51/Y gnd NAND2X1_61/Y vdd NAND2X1
XNAND2X1_94 INVX2_4/Y INVX8_14/A gnd NAND2X1_94/Y vdd NAND2X1
XNAND2X1_72 BUFX4_142/Y NOR2X1_61/Y gnd NAND2X1_72/Y vdd NAND2X1
XNAND2X1_83 BUFX4_324/Y AOI22X1_9/D gnd BUFX4_338/A vdd NAND2X1
XFILL_21_8_0 gnd vdd FILL
XAOI21X1_243 BUFX4_397/Y NOR2X1_303/B NOR2X1_304/Y gnd DFFPOSX1_93/D vdd AOI21X1
XAOI21X1_221 BUFX4_285/Y NOR2X1_265/Y NOR2X1_272/Y gnd AOI21X1_221/Y vdd AOI21X1
XAOI21X1_210 BUFX4_301/Y NOR2X1_256/B NOR2X1_259/Y gnd AOI21X1_210/Y vdd AOI21X1
XAOI21X1_232 BUFX4_423/Y NOR2X1_289/B NOR2X1_287/Y gnd DFFPOSX1_58/D vdd AOI21X1
XAOI21X1_276 BUFX4_96/Y NOR2X1_342/B NOR2X1_347/Y gnd AOI21X1_276/Y vdd AOI21X1
XAOI21X1_265 AOI21X1_3/A NOR2X1_338/B NOR2X1_335/Y gnd AOI21X1_265/Y vdd AOI21X1
XAOI21X1_254 BUFX4_376/Y NOR2X1_315/B NOR2X1_319/Y gnd AOI21X1_254/Y vdd AOI21X1
XAOI21X1_287 BUFX4_423/Y NOR2X1_367/B NOR2X1_361/Y gnd AOI21X1_287/Y vdd AOI21X1
XAOI21X1_298 BUFX4_399/Y NOR2X1_373/B NOR2X1_374/Y gnd AOI21X1_298/Y vdd AOI21X1
XAOI22X1_70 MUX2X1_333/Y BUFX4_349/Y BUFX4_156/Y AOI22X1_70/D gnd AOI22X1_70/Y vdd
+ AOI22X1
XOAI21X1_1471 BUFX4_167/Y BUFX4_393/Y INVX1_456/A gnd OAI21X1_1471/Y vdd OAI21X1
XOAI21X1_1460 NAND2X1_832/Y BUFX4_420/Y OAI21X1_1459/Y gnd OAI21X1_1460/Y vdd OAI21X1
XOAI21X1_1493 BUFX4_462/Y BUFX4_89/Y INVX1_137/A gnd OAI21X1_1494/C vdd OAI21X1
XOAI21X1_1482 BUFX4_397/Y NAND2X1_833/Y OAI21X1_1481/Y gnd OAI21X1_1482/Y vdd OAI21X1
XDFFPOSX1_1001 MUX2X1_25/A CLKBUF1_10/Y AOI21X1_178/Y gnd vdd DFFPOSX1
XFILL_12_8_0 gnd vdd FILL
XDFFPOSX1_1023 NOR2X1_237/A CLKBUF1_3/Y AOI21X1_193/Y gnd vdd DFFPOSX1
XDFFPOSX1_1012 INVX1_252/A CLKBUF1_67/Y OAI21X1_794/Y gnd vdd DFFPOSX1
XFILL_14_2 gnd vdd FILL
XDFFPOSX1_313 OAI21X1_802/B CLKBUF1_53/Y DFFPOSX1_313/D gnd vdd DFFPOSX1
XDFFPOSX1_302 NOR2X1_375/A CLKBUF1_1/Y AOI21X1_299/Y gnd vdd DFFPOSX1
XDFFPOSX1_346 NAND2X1_294/B CLKBUF1_45/Y OAI21X1_1693/Y gnd vdd DFFPOSX1
XDFFPOSX1_324 INVX1_209/A CLKBUF1_85/Y DFFPOSX1_324/D gnd vdd DFFPOSX1
XDFFPOSX1_335 NOR2X1_386/A CLKBUF1_85/Y AOI21X1_308/Y gnd vdd DFFPOSX1
XDFFPOSX1_368 OAI21X1_31/C CLKBUF1_8/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_357 INVX1_275/A CLKBUF1_16/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_379 OAI21X1_53/C CLKBUF1_16/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XNAND2X1_405 BUFX4_234/Y NOR2X1_213/A gnd OAI21X1_974/C vdd NAND2X1
XNAND2X1_427 BUFX4_272/Y NAND2X1_427/B gnd NAND2X1_427/Y vdd NAND2X1
XNAND2X1_416 BUFX4_252/Y NOR2X1_315/A gnd OAI21X1_983/C vdd NAND2X1
XNAND2X1_449 BUFX4_215/Y OAI21X1_335/C gnd NAND2X1_449/Y vdd NAND2X1
XNAND2X1_438 BUFX4_195/Y OAI21X1_159/C gnd NAND2X1_438/Y vdd NAND2X1
XOAI21X1_900 INVX1_112/Y MUX2X1_11/S NAND2X1_326/Y gnd MUX2X1_80/A vdd OAI21X1
XOAI21X1_911 INVX1_123/Y BUFX4_208/Y OAI21X1_911/C gnd MUX2X1_89/B vdd OAI21X1
XOAI21X1_933 INVX1_145/Y BUFX4_252/Y NAND2X1_362/Y gnd MUX2X1_106/B vdd OAI21X1
XOAI21X1_922 INVX1_134/Y BUFX4_230/Y OAI21X1_922/C gnd MUX2X1_97/A vdd OAI21X1
XOAI21X1_955 INVX1_167/Y BUFX4_197/Y NAND2X1_385/Y gnd MUX2X1_122/B vdd OAI21X1
XOAI21X1_944 INVX1_156/Y BUFX4_274/Y OAI21X1_944/C gnd MUX2X1_113/A vdd OAI21X1
XOAI21X1_966 INVX1_178/Y BUFX4_219/Y NAND2X1_397/Y gnd MUX2X1_130/A vdd OAI21X1
XOAI21X1_999 INVX1_211/Y MUX2X1_11/S NAND2X1_433/Y gnd MUX2X1_155/B vdd OAI21X1
XOAI21X1_977 INVX1_189/Y BUFX4_241/Y NAND2X1_410/Y gnd MUX2X1_139/B vdd OAI21X1
XOAI21X1_988 INVX1_200/Y BUFX4_263/Y OAI21X1_988/C gnd MUX2X1_146/A vdd OAI21X1
XOAI21X1_1290 INVX1_502/Y BUFX4_273/Y NAND2X1_746/Y gnd MUX2X1_373/A vdd OAI21X1
XDFFPOSX1_891 NOR2X1_171/A CLKBUF1_32/Y AOI21X1_137/Y gnd vdd DFFPOSX1
XDFFPOSX1_880 NOR2X1_165/A CLKBUF1_81/Y AOI21X1_133/Y gnd vdd DFFPOSX1
XFILL_7_0_1 gnd vdd FILL
XFILL_44_7_0 gnd vdd FILL
XOAI21X1_26 BUFX4_401/Y NAND2X1_2/Y OAI21X1_26/C gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_15 BUFX4_312/Y OAI21X1_7/B INVX1_467/A gnd OAI21X1_16/C vdd OAI21X1
XOAI21X1_59 BUFX4_415/Y BUFX4_314/Y OAI21X1_59/C gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_37 BUFX4_169/Y BUFX4_314/Y INVX1_148/A gnd OAI21X1_38/C vdd OAI21X1
XOAI21X1_48 NAND2X1_3/Y BUFX4_380/Y OAI21X1_48/C gnd OAI21X1_48/Y vdd OAI21X1
XFILL_35_7_0 gnd vdd FILL
XOAI21X1_229 BUFX4_454/Y BUFX4_436/Y INVX1_157/A gnd OAI21X1_229/Y vdd OAI21X1
XOAI21X1_218 INVX1_92/Y NOR2X1_31/Y NAND2X1_40/Y gnd OAI21X1_218/Y vdd OAI21X1
XOAI21X1_207 INVX1_410/Y NOR2X1_11/Y NAND2X1_29/Y gnd OAI21X1_207/Y vdd OAI21X1
XDFFPOSX1_110 NOR2X1_317/A CLKBUF1_39/Y AOI21X1_252/Y gnd vdd DFFPOSX1
XDFFPOSX1_121 NAND2X1_245/B CLKBUF1_20/Y OAI21X1_1394/Y gnd vdd DFFPOSX1
XDFFPOSX1_154 NOR2X1_324/A CLKBUF1_63/Y AOI21X1_256/Y gnd vdd DFFPOSX1
XDFFPOSX1_132 INVX1_197/A CLKBUF1_61/Y DFFPOSX1_132/D gnd vdd DFFPOSX1
XDFFPOSX1_143 NAND2X1_625/B CLKBUF1_102/Y OAI21X1_1438/Y gnd vdd DFFPOSX1
XDFFPOSX1_198 INVX1_329/A CLKBUF1_36/Y DFFPOSX1_198/D gnd vdd DFFPOSX1
XNAND2X1_202 BUFX4_449/Y NOR2X1_228/Y gnd OAI21X1_792/C vdd NAND2X1
XDFFPOSX1_165 INVX1_263/A CLKBUF1_61/Y OAI21X1_1453/Y gnd vdd DFFPOSX1
XDFFPOSX1_176 NOR2X1_340/A CLKBUF1_102/Y AOI21X1_270/Y gnd vdd DFFPOSX1
XDFFPOSX1_187 NAND2X1_352/B CLKBUF1_84/Y DFFPOSX1_187/D gnd vdd DFFPOSX1
XNAND2X1_213 AOI22X1_9/A AOI22X1_6/C gnd BUFX4_92/A vdd NAND2X1
XNAND2X1_235 BUFX4_229/Y NOR2X1_276/A gnd NAND2X1_235/Y vdd NAND2X1
XNAND2X1_224 BUFX4_215/Y OAI21X1_89/C gnd OAI21X1_812/C vdd NAND2X1
XNAND2X1_268 BUFX4_275/Y NOR2X1_83/A gnd OAI21X1_846/C vdd NAND2X1
XNAND2X1_246 BUFX4_57/Y NAND2X1_246/B gnd AOI21X1_204/B vdd NAND2X1
XNAND2X1_257 BUFX4_253/Y NOR2X1_53/A gnd OAI21X1_835/C vdd NAND2X1
XNAND2X1_279 BUFX4_196/Y NAND2X1_279/B gnd OAI21X1_856/C vdd NAND2X1
XFILL_26_7_0 gnd vdd FILL
XFILL_1_7_0 gnd vdd FILL
XNOR2X1_290 NOR2X1_290/A NOR2X1_289/B gnd NOR2X1_290/Y vdd NOR2X1
XOAI21X1_741 BUFX4_281/Y OAI21X1_729/B OAI21X1_741/C gnd OAI21X1_741/Y vdd OAI21X1
XOAI21X1_730 BUFX4_455/Y BUFX4_442/Y INVX1_121/A gnd OAI21X1_730/Y vdd OAI21X1
XOAI21X1_785 BUFX4_400/Y NAND2X1_201/Y OAI21X1_785/C gnd OAI21X1_785/Y vdd OAI21X1
XOAI21X1_774 BUFX4_409/Y BUFX4_443/Y INVX1_506/A gnd OAI21X1_775/C vdd OAI21X1
XOAI21X1_752 NOR2X1_72/B BUFX4_442/Y NAND2X1_542/B gnd OAI21X1_753/C vdd OAI21X1
XOAI21X1_763 BUFX4_419/Y OAI21X1_761/B OAI21X1_763/C gnd OAI21X1_763/Y vdd OAI21X1
XOAI21X1_796 INVX1_380/Y NOR2X1_228/Y NAND2X1_206/Y gnd OAI21X1_796/Y vdd OAI21X1
XMUX2X1_230 MUX2X1_230/A MUX2X1_230/B BUFX4_21/Y gnd MUX2X1_231/A vdd MUX2X1
XMUX2X1_241 MUX2X1_241/A MUX2X1_241/B BUFX4_7/Y gnd MUX2X1_243/B vdd MUX2X1
XMUX2X1_252 MUX2X1_251/Y MUX2X1_250/Y BUFX4_362/Y gnd MUX2X1_252/Y vdd MUX2X1
XMUX2X1_263 MUX2X1_263/A MUX2X1_263/B BUFX4_8/Y gnd MUX2X1_263/Y vdd MUX2X1
XMUX2X1_274 MUX2X1_274/A MUX2X1_274/B BUFX4_56/Y gnd MUX2X1_276/B vdd MUX2X1
XFILL_9_8_0 gnd vdd FILL
XMUX2X1_285 MUX2X1_285/A MUX2X1_285/B BUFX4_362/Y gnd MUX2X1_285/Y vdd MUX2X1
XMUX2X1_296 MUX2X1_296/A MUX2X1_296/B BUFX4_57/Y gnd MUX2X1_297/A vdd MUX2X1
XNAND2X1_780 BUFX4_330/Y NOR2X1_274/Y gnd NAND2X1_780/Y vdd NAND2X1
XNAND2X1_791 AOI22X1_9/A BUFX4_155/Y gnd BUFX4_467/A vdd NAND2X1
XFILL_17_7_0 gnd vdd FILL
XCLKBUF1_16 BUFX4_10/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XCLKBUF1_38 BUFX4_10/Y gnd CLKBUF1_38/Y vdd CLKBUF1
XCLKBUF1_27 BUFX4_14/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XCLKBUF1_49 BUFX4_14/Y gnd CLKBUF1_49/Y vdd CLKBUF1
XBUFX4_70 a[1] gnd BUFX4_70/Y vdd BUFX4
XBUFX4_92 BUFX4_92/A gnd BUFX4_92/Y vdd BUFX4
XBUFX4_81 a[1] gnd BUFX4_81/Y vdd BUFX4
XFILL_41_5_0 gnd vdd FILL
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XOAI21X1_582 BUFX4_281/Y OAI21X1_584/B OAI21X1_582/C gnd OAI21X1_582/Y vdd OAI21X1
XOAI21X1_571 NOR2X1_1/B BUFX4_107/Y INVX1_109/A gnd OAI21X1_572/C vdd OAI21X1
XOAI21X1_593 BUFX4_148/Y BUFX4_107/Y OAI21X1_593/C gnd OAI21X1_594/C vdd OAI21X1
XOAI21X1_560 INVX1_491/Y NOR2X1_91/Y NAND2X1_116/Y gnd OAI21X1_560/Y vdd OAI21X1
XFILL_32_5_0 gnd vdd FILL
XFILL_23_5_0 gnd vdd FILL
XFILL_6_6_0 gnd vdd FILL
XBUFX4_218 BUFX4_29/Y gnd BUFX4_218/Y vdd BUFX4
XBUFX4_207 BUFX4_25/Y gnd BUFX4_207/Y vdd BUFX4
XBUFX4_229 BUFX4_31/Y gnd BUFX4_229/Y vdd BUFX4
XFILL_14_5_0 gnd vdd FILL
XOAI21X1_1119 INVX1_331/Y BUFX4_228/Y NAND2X1_562/Y gnd MUX2X1_245/B vdd OAI21X1
XOAI21X1_1108 INVX1_320/Y BUFX4_206/Y NAND2X1_551/Y gnd MUX2X1_236/A vdd OAI21X1
XOAI21X1_390 NAND2X1_81/Y BUFX4_283/Y OAI21X1_389/Y gnd OAI21X1_390/Y vdd OAI21X1
XINVX1_410 INVX1_410/A gnd INVX1_410/Y vdd INVX1
XDFFPOSX1_709 INVX1_297/A CLKBUF1_46/Y OAI21X1_522/Y gnd vdd DFFPOSX1
XINVX1_443 INVX1_443/A gnd INVX1_443/Y vdd INVX1
XINVX1_432 INVX1_432/A gnd INVX1_432/Y vdd INVX1
XINVX1_421 INVX1_421/A gnd INVX1_421/Y vdd INVX1
XINVX1_487 INVX1_487/A gnd INVX1_487/Y vdd INVX1
XINVX1_465 INVX1_465/A gnd INVX1_465/Y vdd INVX1
XINVX1_476 INVX1_476/A gnd INVX1_476/Y vdd INVX1
XINVX1_454 INVX1_454/A gnd INVX1_454/Y vdd INVX1
XINVX1_498 INVX1_498/A gnd INVX1_498/Y vdd INVX1
XFILL_37_1 gnd vdd FILL
XOAI21X1_1620 INVX1_142/Y NOR2X1_358/Y NAND2X1_846/Y gnd DFFPOSX1_275/D vdd OAI21X1
XOAI21X1_1642 INVX4_3/A BUFX4_346/Y INVX1_272/A gnd OAI21X1_1642/Y vdd OAI21X1
XOAI21X1_1631 INVX1_335/Y NOR2X1_368/Y NAND2X1_857/Y gnd DFFPOSX1_294/D vdd OAI21X1
XOAI21X1_1675 BUFX4_124/Y NAND2X1_871/Y OAI21X1_1675/C gnd DFFPOSX1_337/D vdd OAI21X1
XOAI21X1_1653 BUFX4_420/Y NAND2X1_861/Y OAI21X1_1652/Y gnd OAI21X1_1653/Y vdd OAI21X1
XOAI21X1_1664 BUFX4_412/Y BUFX4_344/Y NAND2X1_706/B gnd OAI21X1_1665/C vdd OAI21X1
XOAI21X1_1686 BUFX4_404/Y OAI21X1_1/B INVX1_402/A gnd OAI21X1_1687/C vdd OAI21X1
XOAI21X1_1697 BUFX4_300/Y NAND2X1_872/Y OAI21X1_1697/C gnd DFFPOSX1_348/D vdd OAI21X1
XNOR2X1_18 NOR2X1_18/A NOR2X1_14/B gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_29 NOR2X1_29/A NOR2X1_27/B gnd NOR2X1_29/Y vdd NOR2X1
XFILL_46_4_0 gnd vdd FILL
XMUX2X1_25 MUX2X1_25/A MUX2X1_25/B BUFX4_194/Y gnd MUX2X1_25/Y vdd MUX2X1
XMUX2X1_36 MUX2X1_35/Y MUX2X1_36/B MUX2X1_69/S gnd MUX2X1_36/Y vdd MUX2X1
XMUX2X1_14 MUX2X1_14/A MUX2X1_14/B MUX2X1_69/S gnd OAI22X1_1/D vdd MUX2X1
XMUX2X1_58 MUX2X1_58/A MUX2X1_58/B BUFX4_34/Y gnd MUX2X1_58/Y vdd MUX2X1
XNOR2X1_108 NOR2X1_108/A NOR2X1_103/B gnd NOR2X1_108/Y vdd NOR2X1
XNOR2X1_119 NOR2X1_119/A NOR2X1_118/B gnd AOI21X1_95/C vdd NOR2X1
XMUX2X1_47 MUX2X1_47/A MUX2X1_47/B BUFX4_42/Y gnd MUX2X1_47/Y vdd MUX2X1
XMUX2X1_69 MUX2X1_69/A MUX2X1_69/B MUX2X1_69/S gnd MUX2X1_69/Y vdd MUX2X1
XFILL_30_8_1 gnd vdd FILL
XDFFPOSX1_517 INVX1_285/A CLKBUF1_1/Y OAI21X1_234/Y gnd vdd DFFPOSX1
XDFFPOSX1_528 NAND2X1_720/B CLKBUF1_57/Y OAI21X1_256/Y gnd vdd DFFPOSX1
XDFFPOSX1_506 NOR2X1_34/A CLKBUF1_24/Y AOI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_539 NOR2X1_45/A CLKBUF1_1/Y AOI21X1_35/Y gnd vdd DFFPOSX1
XINVX1_251 INVX1_251/A gnd INVX1_251/Y vdd INVX1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XINVX1_262 INVX1_262/A gnd INVX1_262/Y vdd INVX1
XNAND2X1_609 BUFX4_216/Y NOR2X1_196/A gnd NAND2X1_609/Y vdd NAND2X1
XINVX1_273 INVX1_273/A gnd INVX1_273/Y vdd INVX1
XINVX1_295 INVX1_295/A gnd INVX1_295/Y vdd INVX1
XINVX1_284 INVX1_284/A gnd INVX1_284/Y vdd INVX1
XNAND2X1_40 BUFX4_452/Y NOR2X1_31/Y gnd NAND2X1_40/Y vdd NAND2X1
XNAND2X1_51 BUFX4_453/Y NOR2X1_41/Y gnd NAND2X1_51/Y vdd NAND2X1
XNAND2X1_95 INVX2_4/Y INVX8_15/A gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_73 BUFX4_445/Y NOR2X1_61/Y gnd NAND2X1_73/Y vdd NAND2X1
XNAND2X1_84 BUFX4_164/Y NOR2X1_71/Y gnd NAND2X1_84/Y vdd NAND2X1
XFILL_37_4_0 gnd vdd FILL
XNAND2X1_62 BUFX4_444/Y NOR2X1_51/Y gnd NAND2X1_62/Y vdd NAND2X1
XAOI21X1_200 NAND2X1_5/B AOI21X1_200/B AOI21X1_195/Y gnd NAND3X1_6/B vdd AOI21X1
XAOI21X1_222 BUFX4_375/Y NOR2X1_265/Y NOR2X1_273/Y gnd DFFPOSX1_48/D vdd AOI21X1
XAOI21X1_211 BUFX4_395/Y NOR2X1_256/B NOR2X1_260/Y gnd DFFPOSX1_13/D vdd AOI21X1
XFILL_20_3_0 gnd vdd FILL
XAOI21X1_233 AOI21X1_3/A NOR2X1_289/B NOR2X1_288/Y gnd DFFPOSX1_59/D vdd AOI21X1
XFILL_21_8_1 gnd vdd FILL
XAOI21X1_266 BUFX4_304/Y NOR2X1_338/B NOR2X1_336/Y gnd AOI21X1_266/Y vdd AOI21X1
XAOI21X1_255 BUFX4_125/Y NOR2X1_325/B NOR2X1_323/Y gnd AOI21X1_255/Y vdd AOI21X1
XAOI21X1_244 BUFX4_99/Y NOR2X1_303/B NOR2X1_305/Y gnd DFFPOSX1_94/D vdd AOI21X1
XAOI21X1_277 BUFX4_282/Y NOR2X1_342/B NOR2X1_348/Y gnd AOI21X1_277/Y vdd AOI21X1
XAOI22X1_60 MUX2X1_285/Y BUFX4_354/Y BUFX4_155/Y AOI22X1_60/D gnd AOI22X1_60/Y vdd
+ AOI22X1
XAOI21X1_288 BUFX4_114/Y NOR2X1_367/B NOR2X1_362/Y gnd AOI21X1_288/Y vdd AOI21X1
XAOI21X1_299 BUFX4_97/Y NOR2X1_373/B NOR2X1_375/Y gnd AOI21X1_299/Y vdd AOI21X1
XAOI22X1_71 AOI22X1_71/A INVX1_10/A AOI22X1_6/C MUX2X1_342/Y gnd AOI22X1_71/Y vdd
+ AOI22X1
XOAI21X1_1450 INVX1_71/Y NOR2X1_331/Y NAND2X1_825/Y gnd DFFPOSX1_162/D vdd OAI21X1
XOAI21X1_1472 NAND2X1_832/Y BUFX4_373/Y OAI21X1_1471/Y gnd DFFPOSX1_184/D vdd OAI21X1
XOAI21X1_1483 BUFX4_417/Y BUFX4_392/Y NAND2X1_559/B gnd OAI21X1_1483/Y vdd OAI21X1
XOAI21X1_1461 BUFX4_167/Y BUFX4_393/Y INVX1_136/A gnd OAI21X1_1461/Y vdd OAI21X1
XOAI21X1_1494 BUFX4_115/Y NAND2X1_834/Y OAI21X1_1494/C gnd DFFPOSX1_195/D vdd OAI21X1
XFILL_3_4_0 gnd vdd FILL
XFILL_28_4_0 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XFILL_12_8_1 gnd vdd FILL
XDFFPOSX1_1002 NOR2X1_221/A CLKBUF1_85/Y AOI21X1_179/Y gnd vdd DFFPOSX1
XDFFPOSX1_1024 NOR2X1_238/A CLKBUF1_97/Y AOI21X1_194/Y gnd vdd DFFPOSX1
XDFFPOSX1_1013 INVX1_316/A CLKBUF1_3/Y OAI21X1_795/Y gnd vdd DFFPOSX1
XFILL_19_4_0 gnd vdd FILL
XDFFPOSX1_303 NOR2X1_376/A CLKBUF1_25/Y AOI21X1_300/Y gnd vdd DFFPOSX1
XDFFPOSX1_325 INVX1_273/A CLKBUF1_70/Y DFFPOSX1_325/D gnd vdd DFFPOSX1
XDFFPOSX1_347 NAND2X1_363/B CLKBUF1_38/Y DFFPOSX1_347/D gnd vdd DFFPOSX1
XDFFPOSX1_336 NOR2X1_387/A CLKBUF1_83/Y AOI21X1_309/Y gnd vdd DFFPOSX1
XDFFPOSX1_314 NAND2X1_292/B CLKBUF1_55/Y OAI21X1_1653/Y gnd vdd DFFPOSX1
XDFFPOSX1_369 INVX1_21/A CLKBUF1_8/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_358 INVX1_339/A CLKBUF1_34/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XNAND2X1_406 BUFX4_236/Y NOR2X1_222/A gnd OAI21X1_975/C vdd NAND2X1
XNAND2X1_417 BUFX4_254/Y NAND2X1_417/B gnd OAI21X1_984/C vdd NAND2X1
XNAND2X1_439 BUFX4_197/Y OAI21X1_191/C gnd NAND2X1_439/Y vdd NAND2X1
XNAND2X1_428 BUFX4_274/Y NOR2X1_363/A gnd OAI21X1_994/C vdd NAND2X1
XBUFX4_390 BUFX4_392/A gnd BUFX4_390/Y vdd BUFX4
XOAI21X1_934 INVX1_146/Y BUFX4_254/Y NAND2X1_363/Y gnd MUX2X1_106/A vdd OAI21X1
XOAI21X1_912 INVX1_124/Y BUFX4_210/Y NAND2X1_338/Y gnd MUX2X1_89/A vdd OAI21X1
XOAI21X1_923 INVX1_135/Y BUFX4_232/Y OAI21X1_923/C gnd MUX2X1_98/B vdd OAI21X1
XOAI21X1_901 INVX1_113/Y BUFX4_188/Y OAI21X1_901/C gnd MUX2X1_82/B vdd OAI21X1
XOAI21X1_945 INVX1_157/Y BUFX4_276/Y OAI21X1_945/C gnd MUX2X1_115/B vdd OAI21X1
XOAI21X1_967 INVX1_179/Y BUFX4_221/Y OAI21X1_967/C gnd MUX2X1_131/B vdd OAI21X1
XOAI21X1_956 INVX1_168/Y BUFX4_199/Y NAND2X1_386/Y gnd MUX2X1_122/A vdd OAI21X1
XOAI21X1_989 INVX1_201/Y BUFX4_265/Y NAND2X1_422/Y gnd MUX2X1_148/B vdd OAI21X1
XOAI21X1_978 INVX1_190/Y BUFX4_243/Y NAND2X1_411/Y gnd MUX2X1_139/A vdd OAI21X1
XOAI21X1_1291 INVX1_503/Y BUFX4_275/Y NAND2X1_747/Y gnd MUX2X1_374/B vdd OAI21X1
XOAI21X1_1280 INVX1_492/Y BUFX4_253/Y NAND2X1_735/Y gnd MUX2X1_365/A vdd OAI21X1
XDFFPOSX1_892 NOR2X1_172/A CLKBUF1_95/Y AOI21X1_138/Y gnd vdd DFFPOSX1
XDFFPOSX1_881 MUX2X1_12/B CLKBUF1_11/Y AOI21X1_134/Y gnd vdd DFFPOSX1
XDFFPOSX1_870 INVX1_371/A CLKBUF1_13/Y OAI21X1_665/Y gnd vdd DFFPOSX1
XFILL_44_7_1 gnd vdd FILL
XFILL_43_2_0 gnd vdd FILL
XOAI21X1_16 BUFX4_380/Y NAND2X1_1/Y OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_49 BUFX4_410/Y OAI21X1_1/B OAI21X1_49/C gnd OAI21X1_50/C vdd OAI21X1
XOAI21X1_27 BUFX4_367/Y BUFX4_314/Y OAI21X1_27/C gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_38 NAND2X1_3/Y BUFX4_109/Y OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XFILL_35_7_1 gnd vdd FILL
XFILL_34_2_0 gnd vdd FILL
XOAI21X1_208 INVX1_474/Y NOR2X1_11/Y NAND2X1_30/Y gnd OAI21X1_208/Y vdd OAI21X1
XOAI21X1_219 INVX1_156/Y NOR2X1_31/Y NAND2X1_41/Y gnd OAI21X1_219/Y vdd OAI21X1
XDFFPOSX1_100 INVX1_195/A CLKBUF1_25/Y DFFPOSX1_100/D gnd vdd DFFPOSX1
XDFFPOSX1_111 NOR2X1_318/A CLKBUF1_39/Y AOI21X1_253/Y gnd vdd DFFPOSX1
XDFFPOSX1_133 INVX1_261/A CLKBUF1_55/Y DFFPOSX1_133/D gnd vdd DFFPOSX1
XDFFPOSX1_155 NOR2X1_325/A CLKBUF1_102/Y AOI21X1_257/Y gnd vdd DFFPOSX1
XDFFPOSX1_144 NAND2X1_694/B CLKBUF1_20/Y OAI21X1_1440/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 NAND2X1_279/B CLKBUF1_17/Y DFFPOSX1_122/D gnd vdd DFFPOSX1
XDFFPOSX1_166 INVX1_327/A CLKBUF1_98/Y OAI21X1_1454/Y gnd vdd DFFPOSX1
XDFFPOSX1_188 NAND2X1_421/B CLKBUF1_78/Y OAI21X1_1480/Y gnd vdd DFFPOSX1
XDFFPOSX1_177 INVX1_44/A CLKBUF1_43/Y DFFPOSX1_177/D gnd vdd DFFPOSX1
XDFFPOSX1_199 INVX1_393/A CLKBUF1_36/Y OAI21X1_1502/Y gnd vdd DFFPOSX1
XNAND2X1_203 NAND2X1_8/A NOR2X1_228/Y gnd OAI21X1_793/C vdd NAND2X1
XNAND2X1_225 BUFX4_217/Y NOR2X1_3/A gnd OAI21X1_813/C vdd NAND2X1
XNAND2X1_214 BUFX4_201/Y NOR2X1_370/A gnd OAI21X1_803/C vdd NAND2X1
XNAND2X1_236 INVX4_1/Y NAND2X1_236/B gnd NAND2X1_236/Y vdd NAND2X1
XNAND2X1_247 BUFX4_241/Y NAND2X1_247/B gnd OAI21X1_828/C vdd NAND2X1
XNAND2X1_269 BUFX4_277/Y NOR2X1_93/A gnd OAI21X1_847/C vdd NAND2X1
XNAND2X1_258 BUFX4_255/Y NAND2X1_258/B gnd NAND2X1_258/Y vdd NAND2X1
XFILL_0_2_0 gnd vdd FILL
XFILL_1_7_1 gnd vdd FILL
XFILL_25_2_0 gnd vdd FILL
XFILL_26_7_1 gnd vdd FILL
XNOR2X1_291 NOR2X1_291/A NOR2X1_289/B gnd NOR2X1_291/Y vdd NOR2X1
XNOR2X1_280 NOR2X1_280/A NOR2X1_279/B gnd NOR2X1_280/Y vdd NOR2X1
XOAI21X1_720 INVX1_503/Y NOR2X1_189/B OAI21X1_720/C gnd OAI21X1_720/Y vdd OAI21X1
XOAI21X1_731 BUFX4_419/Y OAI21X1_729/B OAI21X1_730/Y gnd OAI21X1_731/Y vdd OAI21X1
XOAI21X1_742 BUFX4_455/Y BUFX4_440/Y INVX1_505/A gnd OAI21X1_743/C vdd OAI21X1
XOAI21X1_775 BUFX4_378/Y OAI21X1_761/B OAI21X1_775/C gnd OAI21X1_775/Y vdd OAI21X1
XOAI21X1_764 BUFX4_409/Y BUFX4_443/Y INVX1_186/A gnd OAI21X1_765/C vdd OAI21X1
XOAI21X1_753 BUFX4_400/Y OAI21X1_757/B OAI21X1_753/C gnd OAI21X1_753/Y vdd OAI21X1
XOAI21X1_797 INVX1_444/Y NOR2X1_228/Y OAI21X1_797/C gnd OAI21X1_797/Y vdd OAI21X1
XOAI21X1_786 NOR2X1_91/B BUFX4_441/Y INVX1_379/A gnd OAI21X1_787/C vdd OAI21X1
XMUX2X1_231 MUX2X1_231/A MUX2X1_229/Y MUX2X1_7/S gnd MUX2X1_231/Y vdd MUX2X1
XMUX2X1_220 MUX2X1_220/A MUX2X1_220/B BUFX4_37/Y gnd MUX2X1_222/B vdd MUX2X1
XMUX2X1_264 MUX2X1_263/Y MUX2X1_262/Y MUX2X1_7/S gnd MUX2X1_264/Y vdd MUX2X1
XMUX2X1_253 MUX2X1_253/A MUX2X1_253/B BUFX4_22/Y gnd MUX2X1_255/B vdd MUX2X1
XMUX2X1_242 MUX2X1_242/A MUX2X1_242/B BUFX4_38/Y gnd MUX2X1_243/A vdd MUX2X1
XFILL_9_8_1 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XMUX2X1_297 MUX2X1_297/A MUX2X1_297/B MUX2X1_7/S gnd AOI22X1_62/A vdd MUX2X1
XMUX2X1_286 MUX2X1_286/A MUX2X1_286/B BUFX4_5/Y gnd MUX2X1_288/B vdd MUX2X1
XMUX2X1_275 MUX2X1_275/A MUX2X1_275/B BUFX4_19/Y gnd MUX2X1_276/A vdd MUX2X1
XNAND2X1_770 BUFX4_447/Y NOR2X1_264/Y gnd NAND2X1_770/Y vdd NAND2X1
XNAND2X1_781 BUFX4_140/Y NOR2X1_274/Y gnd NAND2X1_781/Y vdd NAND2X1
XNAND2X1_792 INVX8_10/A INVX2_7/Y gnd NAND2X1_792/Y vdd NAND2X1
XFILL_16_2_0 gnd vdd FILL
XFILL_17_7_1 gnd vdd FILL
XCLKBUF1_17 BUFX4_12/Y gnd CLKBUF1_17/Y vdd CLKBUF1
XCLKBUF1_28 BUFX4_10/Y gnd CLKBUF1_28/Y vdd CLKBUF1
XCLKBUF1_39 BUFX4_14/Y gnd CLKBUF1_39/Y vdd CLKBUF1
XBUFX4_60 BUFX4_62/A gnd BUFX4_60/Y vdd BUFX4
XBUFX4_71 a[1] gnd BUFX4_71/Y vdd BUFX4
XBUFX4_82 a[1] gnd BUFX4_82/Y vdd BUFX4
XBUFX4_93 BUFX4_92/A gnd BUFX4_93/Y vdd BUFX4
XOR2X2_1 OR2X2_1/A INVX8_1/Y gnd OR2X2_1/Y vdd OR2X2
XFILL_41_5_1 gnd vdd FILL
XFILL_40_0_0 gnd vdd FILL
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XOAI21X1_550 INVX1_362/Y NOR2X1_81/Y OAI21X1_550/C gnd OAI21X1_550/Y vdd OAI21X1
XOAI21X1_572 BUFX4_418/Y OAI21X1_584/B OAI21X1_572/C gnd OAI21X1_572/Y vdd OAI21X1
XOAI21X1_583 NOR2X1_1/B INVX1_3/A INVX1_493/A gnd OAI21X1_583/Y vdd OAI21X1
XOAI21X1_561 INVX1_60/Y NOR2X1_101/Y NAND2X1_117/Y gnd OAI21X1_561/Y vdd OAI21X1
XOAI21X1_594 BUFX4_396/Y OAI21X1_590/B OAI21X1_594/C gnd OAI21X1_594/Y vdd OAI21X1
XFILL_48_1_0 gnd vdd FILL
XFILL_32_5_1 gnd vdd FILL
XFILL_31_0_0 gnd vdd FILL
XFILL_39_1_0 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XFILL_23_5_1 gnd vdd FILL
XFILL_6_6_1 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XBUFX4_219 BUFX4_24/Y gnd BUFX4_219/Y vdd BUFX4
XBUFX4_208 BUFX4_26/Y gnd BUFX4_208/Y vdd BUFX4
XFILL_13_0_0 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XOAI21X1_1109 INVX1_321/Y BUFX4_208/Y NAND2X1_552/Y gnd MUX2X1_238/B vdd OAI21X1
XINVX1_400 INVX1_400/A gnd INVX1_400/Y vdd INVX1
XOAI21X1_380 NAND2X1_81/Y BUFX4_421/Y OAI21X1_380/C gnd OAI21X1_380/Y vdd OAI21X1
XOAI21X1_391 BUFX4_169/Y BUFX4_386/Y INVX1_484/A gnd OAI21X1_392/C vdd OAI21X1
XINVX1_411 INVX1_411/A gnd INVX1_411/Y vdd INVX1
XINVX1_433 INVX1_433/A gnd INVX1_433/Y vdd INVX1
XINVX1_422 INVX1_422/A gnd INVX1_422/Y vdd INVX1
XINVX1_444 INVX1_444/A gnd INVX1_444/Y vdd INVX1
XINVX1_477 INVX1_477/A gnd INVX1_477/Y vdd INVX1
XINVX1_466 INVX1_466/A gnd INVX1_466/Y vdd INVX1
XINVX1_455 INVX1_455/A gnd INVX1_455/Y vdd INVX1
XINVX1_488 INVX1_488/A gnd INVX1_488/Y vdd INVX1
XINVX1_499 INVX1_499/A gnd INVX1_499/Y vdd INVX1
XOAI21X1_1610 NOR2X1_2/B BUFX4_345/Y NAND2X1_496/B gnd OAI21X1_1610/Y vdd OAI21X1
XOAI21X1_1621 INVX1_206/Y NOR2X1_358/Y NAND2X1_847/Y gnd DFFPOSX1_276/D vdd OAI21X1
XOAI21X1_1632 INVX1_399/Y NOR2X1_368/Y NAND2X1_858/Y gnd DFFPOSX1_295/D vdd OAI21X1
XOAI21X1_1654 BUFX4_412/Y BUFX4_343/Y NAND2X1_361/B gnd OAI21X1_1654/Y vdd OAI21X1
XOAI21X1_1643 NAND2X1_860/Y BUFX4_399/Y OAI21X1_1642/Y gnd OAI21X1_1643/Y vdd OAI21X1
XOAI21X1_1665 BUFX4_376/Y NAND2X1_861/Y OAI21X1_1665/C gnd OAI21X1_1665/Y vdd OAI21X1
XOAI21X1_1687 BUFX4_283/Y NAND2X1_871/Y OAI21X1_1687/C gnd OAI21X1_1687/Y vdd OAI21X1
XOAI21X1_1698 BUFX4_83/Y INVX2_11/A NAND2X1_501/B gnd OAI21X1_1699/C vdd OAI21X1
XOAI21X1_1676 BUFX4_406/Y OAI21X1_5/B INVX1_82/A gnd OAI21X1_1677/C vdd OAI21X1
XNOR2X1_19 NOR2X1_19/A NOR2X1_14/B gnd NOR2X1_19/Y vdd NOR2X1
XFILL_46_4_1 gnd vdd FILL
XMUX2X1_26 MUX2X1_26/A MUX2X1_26/B BUFX4_195/Y gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_15 MUX2X1_15/A MUX2X1_15/B BUFX4_188/Y gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_59 MUX2X1_59/A MUX2X1_59/B BUFX4_54/Y gnd MUX2X1_59/Y vdd MUX2X1
XMUX2X1_37 MUX2X1_37/A MUX2X1_37/B BUFX4_53/Y gnd MUX2X1_39/B vdd MUX2X1
XNOR2X1_109 NOR2X1_109/A NOR2X1_103/B gnd NOR2X1_109/Y vdd NOR2X1
XMUX2X1_48 MUX2X1_47/Y MUX2X1_48/B MUX2X1_48/S gnd MUX2X1_48/Y vdd MUX2X1
XDFFPOSX1_518 INVX1_349/A CLKBUF1_91/Y OAI21X1_236/Y gnd vdd DFFPOSX1
XDFFPOSX1_529 INVX1_46/A CLKBUF1_1/Y OAI21X1_257/Y gnd vdd DFFPOSX1
XDFFPOSX1_507 NOR2X1_35/A CLKBUF1_24/Y AOI21X1_27/Y gnd vdd DFFPOSX1
XINVX1_241 INVX1_241/A gnd INVX1_241/Y vdd INVX1
XINVX1_230 INVX1_230/A gnd INVX1_230/Y vdd INVX1
XINVX1_252 INVX1_252/A gnd INVX1_252/Y vdd INVX1
XINVX1_285 INVX1_285/A gnd INVX1_285/Y vdd INVX1
XINVX1_274 INVX1_274/A gnd INVX1_274/Y vdd INVX1
XINVX1_263 INVX1_263/A gnd INVX1_263/Y vdd INVX1
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XNAND2X1_30 BUFX4_428/Y NOR2X1_11/Y gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_41 BUFX4_334/Y NOR2X1_31/Y gnd NAND2X1_41/Y vdd NAND2X1
XNAND2X1_52 BUFX4_335/Y NOR2X1_41/Y gnd NAND2X1_52/Y vdd NAND2X1
XNAND2X1_74 BUFX4_327/Y NOR2X1_61/Y gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_85 INVX8_3/A NOR2X1_71/Y gnd NAND2X1_85/Y vdd NAND2X1
XFILL_37_4_1 gnd vdd FILL
XNAND2X1_63 BUFX4_326/Y NOR2X1_51/Y gnd NAND2X1_63/Y vdd NAND2X1
XNAND2X1_96 INVX2_4/Y INVX4_3/Y gnd NAND2X1_96/Y vdd NAND2X1
XAOI21X1_212 BUFX4_98/Y NOR2X1_256/B NOR2X1_261/Y gnd DFFPOSX1_14/D vdd AOI21X1
XAOI21X1_201 AOI21X1_201/A AOI21X1_201/B BUFX4_363/Y gnd AOI21X1_201/Y vdd AOI21X1
XAOI21X1_223 AOI21X1_1/A NOR2X1_279/B NOR2X1_276/Y gnd DFFPOSX1_17/D vdd AOI21X1
XFILL_20_3_1 gnd vdd FILL
XAOI21X1_234 BUFX4_304/Y NOR2X1_289/B NOR2X1_289/Y gnd AOI21X1_234/Y vdd AOI21X1
XAOI21X1_256 BUFX4_423/Y NOR2X1_325/B NOR2X1_324/Y gnd AOI21X1_256/Y vdd AOI21X1
XAOI21X1_267 BUFX4_397/Y NOR2X1_338/B NOR2X1_337/Y gnd AOI21X1_267/Y vdd AOI21X1
XAOI21X1_245 BUFX4_286/Y NOR2X1_303/B NOR2X1_306/Y gnd DFFPOSX1_95/D vdd AOI21X1
XAOI21X1_278 BUFX4_375/Y NOR2X1_342/B NOR2X1_349/Y gnd AOI21X1_278/Y vdd AOI21X1
XAOI22X1_50 MUX2X1_237/Y BUFX4_349/Y BUFX4_156/Y AOI22X1_50/D gnd AOI22X1_50/Y vdd
+ AOI22X1
XAOI21X1_289 BUFX4_297/Y NOR2X1_367/B NOR2X1_363/Y gnd AOI21X1_289/Y vdd AOI21X1
XAOI22X1_72 AOI22X1_72/A BUFX4_352/Y BUFX4_157/Y MUX2X1_348/Y gnd AOI22X1_72/Y vdd
+ AOI22X1
XAOI22X1_61 AOI22X1_61/A BUFX4_321/Y BUFX4_288/Y MUX2X1_294/Y gnd AOI22X1_61/Y vdd
+ AOI22X1
XOAI21X1_1440 BUFX4_373/Y NAND2X1_815/Y OAI21X1_1439/Y gnd OAI21X1_1440/Y vdd OAI21X1
XOAI21X1_1462 NAND2X1_832/Y BUFX4_112/Y OAI21X1_1461/Y gnd OAI21X1_1462/Y vdd OAI21X1
XOAI21X1_1484 BUFX4_99/Y NAND2X1_833/Y OAI21X1_1483/Y gnd OAI21X1_1484/Y vdd OAI21X1
XOAI21X1_1451 INVX1_135/Y NOR2X1_331/Y NAND2X1_826/Y gnd OAI21X1_1451/Y vdd OAI21X1
XOAI21X1_1473 BUFX4_417/Y BUFX4_392/Y NAND2X1_253/B gnd OAI21X1_1473/Y vdd OAI21X1
XOAI21X1_1495 NOR2X1_61/B BUFX4_89/Y INVX1_201/A gnd OAI21X1_1496/C vdd OAI21X1
XFILL_28_4_1 gnd vdd FILL
XFILL_3_4_1 gnd vdd FILL
XDFFPOSX1_1025 BUFX2_1/A CLKBUF1_91/Y NAND3X1_6/Y gnd vdd DFFPOSX1
XFILL_11_3_1 gnd vdd FILL
XDFFPOSX1_1003 NOR2X1_222/A CLKBUF1_40/Y AOI21X1_180/Y gnd vdd DFFPOSX1
XDFFPOSX1_1014 INVX1_380/A CLKBUF1_83/Y OAI21X1_796/Y gnd vdd DFFPOSX1
XOAI22X1_1 MUX2X1_7/Y INVX1_6/Y INVX1_8/Y OAI22X1_1/D gnd OAI22X1_1/Y vdd OAI22X1
XFILL_19_4_1 gnd vdd FILL
XDFFPOSX1_304 NOR2X1_377/A CLKBUF1_11/Y AOI21X1_301/Y gnd vdd DFFPOSX1
XDFFPOSX1_315 NAND2X1_361/B CLKBUF1_53/Y OAI21X1_1655/Y gnd vdd DFFPOSX1
XDFFPOSX1_337 INVX1_23/A CLKBUF1_47/Y DFFPOSX1_337/D gnd vdd DFFPOSX1
XDFFPOSX1_326 INVX1_337/A CLKBUF1_79/Y OAI21X1_1671/Y gnd vdd DFFPOSX1
XDFFPOSX1_348 NAND2X1_432/B CLKBUF1_47/Y DFFPOSX1_348/D gnd vdd DFFPOSX1
XDFFPOSX1_359 INVX1_403/A CLKBUF1_64/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XNAND2X1_407 BUFX4_238/Y NOR2X1_233/A gnd NAND2X1_407/Y vdd NAND2X1
XNAND2X1_418 BUFX4_256/Y NAND2X1_418/B gnd OAI21X1_985/C vdd NAND2X1
XNAND2X1_429 BUFX4_276/Y NOR2X1_373/A gnd OAI21X1_995/C vdd NAND2X1
XBUFX4_380 INVX8_9/Y gnd BUFX4_380/Y vdd BUFX4
XBUFX4_391 BUFX4_392/A gnd INVX2_8/A vdd BUFX4
XOAI21X1_924 INVX1_136/Y BUFX4_234/Y NAND2X1_352/Y gnd MUX2X1_98/A vdd OAI21X1
XOAI21X1_913 INVX1_125/Y BUFX4_212/Y NAND2X1_341/Y gnd MUX2X1_91/B vdd OAI21X1
XOAI21X1_902 INVX1_114/Y BUFX4_190/Y OAI21X1_902/C gnd MUX2X1_82/A vdd OAI21X1
XOAI21X1_935 INVX1_147/Y BUFX4_256/Y NAND2X1_364/Y gnd MUX2X1_107/B vdd OAI21X1
XOAI21X1_957 INVX1_169/Y BUFX4_201/Y OAI21X1_957/C gnd MUX2X1_124/B vdd OAI21X1
XOAI21X1_946 INVX1_158/Y BUFX4_278/Y OAI21X1_946/C gnd MUX2X1_115/A vdd OAI21X1
XOAI21X1_968 INVX1_180/Y BUFX4_223/Y OAI21X1_968/C gnd MUX2X1_131/A vdd OAI21X1
XOAI21X1_979 INVX1_191/Y BUFX4_245/Y NAND2X1_412/Y gnd MUX2X1_140/B vdd OAI21X1
XDFFPOSX1_860 NOR2X1_150/A CLKBUF1_7/Y AOI21X1_120/Y gnd vdd DFFPOSX1
XOAI21X1_1270 INVX1_482/Y BUFX4_233/Y NAND2X1_725/Y gnd MUX2X1_358/A vdd OAI21X1
XOAI21X1_1292 INVX1_504/Y BUFX4_277/Y NAND2X1_748/Y gnd MUX2X1_374/A vdd OAI21X1
XOAI21X1_1281 INVX1_493/Y BUFX4_255/Y NAND2X1_737/Y gnd MUX2X1_367/B vdd OAI21X1
XDFFPOSX1_893 NOR2X1_173/A CLKBUF1_32/Y AOI21X1_139/Y gnd vdd DFFPOSX1
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XDFFPOSX1_882 INVX1_116/A CLKBUF1_92/Y OAI21X1_668/Y gnd vdd DFFPOSX1
XDFFPOSX1_871 INVX1_435/A CLKBUF1_27/Y OAI21X1_666/Y gnd vdd DFFPOSX1
XFILL_43_2_1 gnd vdd FILL
XOAI21X1_17 BUFX4_367/Y BUFX4_317/Y OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_28 BUFX4_102/Y NAND2X1_2/Y OAI21X1_27/Y gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_39 BUFX4_169/Y OAI21X1_7/B INVX1_212/A gnd OAI21X1_40/C vdd OAI21X1
XFILL_34_2_1 gnd vdd FILL
XOAI21X1_209 INVX1_30/Y NOR2X1_21/Y NAND2X1_31/Y gnd OAI21X1_209/Y vdd OAI21X1
XDFFPOSX1_101 INVX1_259/A CLKBUF1_55/Y OAI21X1_1373/Y gnd vdd DFFPOSX1
XDFFPOSX1_112 NOR2X1_319/A CLKBUF1_25/Y AOI21X1_254/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 INVX1_42/A CLKBUF1_63/Y OAI21X1_1441/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 INVX1_325/A CLKBUF1_55/Y OAI21X1_1420/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 NAND2X1_348/B CLKBUF1_20/Y OAI21X1_1398/Y gnd vdd DFFPOSX1
XDFFPOSX1_178 INVX1_72/A CLKBUF1_43/Y OAI21X1_1460/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 NOR2X1_326/A CLKBUF1_12/Y AOI21X1_258/Y gnd vdd DFFPOSX1
XDFFPOSX1_167 INVX1_391/A CLKBUF1_98/Y OAI21X1_1455/Y gnd vdd DFFPOSX1
XDFFPOSX1_189 NAND2X1_490/B CLKBUF1_84/Y OAI21X1_1482/Y gnd vdd DFFPOSX1
XNAND2X1_204 NAND2X1_9/A NOR2X1_228/Y gnd OAI21X1_794/C vdd NAND2X1
XNAND2X1_226 BUFX4_219/Y NOR2X1_23/A gnd OAI21X1_815/C vdd NAND2X1
XNAND2X1_215 NOR2X1_244/Y NAND2X1_215/B gnd NAND3X1_1/B vdd NAND2X1
XNAND2X1_259 BUFX4_257/Y NOR2X1_63/A gnd OAI21X1_837/C vdd NAND2X1
XNAND2X1_237 BUFX4_231/Y NOR2X1_286/A gnd OAI21X1_821/C vdd NAND2X1
XNAND2X1_248 INVX4_1/Y NAND2X1_248/B gnd AOI21X1_205/A vdd NAND2X1
XFILL_25_2_1 gnd vdd FILL
XNOR2X1_270 NOR2X1_270/A NOR2X1_265/Y gnd NOR2X1_270/Y vdd NOR2X1
XFILL_0_2_1 gnd vdd FILL
XNOR2X1_292 NOR2X1_292/A NOR2X1_289/B gnd NOR2X1_292/Y vdd NOR2X1
XNOR2X1_281 NOR2X1_281/A NOR2X1_279/B gnd NOR2X1_281/Y vdd NOR2X1
XOAI21X1_721 INVX1_120/Y NOR2X1_199/Y OAI21X1_721/C gnd OAI21X1_721/Y vdd OAI21X1
XOAI21X1_710 INVX1_310/Y NOR2X1_177/Y OAI21X1_710/C gnd OAI21X1_710/Y vdd OAI21X1
XOAI21X1_732 BUFX4_455/Y BUFX4_441/Y INVX1_185/A gnd OAI21X1_733/C vdd OAI21X1
XOAI21X1_776 BUFX4_308/Y BUFX4_438/Y MUX2X1_25/B gnd OAI21X1_777/C vdd OAI21X1
XOAI21X1_765 BUFX4_117/Y OAI21X1_761/B OAI21X1_765/C gnd OAI21X1_765/Y vdd OAI21X1
XOAI21X1_754 NOR2X1_72/B BUFX4_441/Y NAND2X1_611/B gnd OAI21X1_754/Y vdd OAI21X1
XOAI21X1_743 BUFX4_378/Y OAI21X1_729/B OAI21X1_743/C gnd OAI21X1_743/Y vdd OAI21X1
XOAI21X1_798 INVX1_508/Y NOR2X1_228/Y OAI21X1_798/C gnd OAI21X1_798/Y vdd OAI21X1
XOAI21X1_787 BUFX4_103/Y NAND2X1_201/Y OAI21X1_787/C gnd OAI21X1_787/Y vdd OAI21X1
XMUX2X1_232 MUX2X1_232/A MUX2X1_232/B BUFX4_46/Y gnd MUX2X1_232/Y vdd MUX2X1
XMUX2X1_210 MUX2X1_210/A MUX2X1_208/Y INVX2_6/A gnd AOI22X1_43/D vdd MUX2X1
XMUX2X1_221 MUX2X1_221/A MUX2X1_221/B INVX4_1/A gnd MUX2X1_222/A vdd MUX2X1
XMUX2X1_265 MUX2X1_265/A MUX2X1_265/B BUFX4_39/Y gnd MUX2X1_267/B vdd MUX2X1
XMUX2X1_243 MUX2X1_243/A MUX2X1_243/B INVX2_6/A gnd AOI22X1_51/A vdd MUX2X1
XMUX2X1_254 MUX2X1_254/A MUX2X1_254/B BUFX4_47/Y gnd MUX2X1_255/A vdd MUX2X1
XDFFPOSX1_690 INVX1_104/A CLKBUF1_58/Y OAI21X1_484/Y gnd vdd DFFPOSX1
XMUX2X1_298 MUX2X1_298/A MUX2X1_298/B BUFX4_20/Y gnd MUX2X1_298/Y vdd MUX2X1
XMUX2X1_287 MUX2X1_287/A MUX2X1_287/B BUFX4_36/Y gnd MUX2X1_288/A vdd MUX2X1
XMUX2X1_276 MUX2X1_276/A MUX2X1_276/B INVX2_6/A gnd AOI22X1_57/D vdd MUX2X1
XFILL_8_3_1 gnd vdd FILL
XNAND2X1_771 BUFX4_329/Y NOR2X1_264/Y gnd NAND2X1_771/Y vdd NAND2X1
XNAND2X1_760 BUFX4_445/Y NOR2X1_254/Y gnd NAND2X1_760/Y vdd NAND2X1
XNAND2X1_782 BUFX4_431/Y NOR2X1_274/Y gnd NAND2X1_782/Y vdd NAND2X1
XNAND2X1_793 INVX8_11/A INVX2_7/Y gnd NAND2X1_793/Y vdd NAND2X1
XFILL_16_2_1 gnd vdd FILL
XCLKBUF1_18 BUFX4_16/Y gnd CLKBUF1_18/Y vdd CLKBUF1
XCLKBUF1_29 BUFX4_9/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XBUFX4_50 BUFX4_50/A gnd BUFX4_50/Y vdd BUFX4
XBUFX4_61 BUFX4_62/A gnd BUFX4_61/Y vdd BUFX4
XBUFX4_83 BUFX4_84/A gnd BUFX4_83/Y vdd BUFX4
XBUFX4_94 BUFX4_92/A gnd BUFX4_94/Y vdd BUFX4
XBUFX4_72 a[1] gnd BUFX4_62/A vdd BUFX4
XFILL_40_0_1 gnd vdd FILL
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XOAI21X1_540 AOI21X1_6/A OAI21X1_544/B OAI21X1_539/Y gnd OAI21X1_540/Y vdd OAI21X1
XOAI21X1_551 INVX1_426/Y NOR2X1_81/Y OAI21X1_551/C gnd OAI21X1_551/Y vdd OAI21X1
XOAI21X1_573 NOR2X1_1/B BUFX4_107/Y INVX1_173/A gnd OAI21X1_574/C vdd OAI21X1
XOAI21X1_584 BUFX4_372/Y OAI21X1_584/B OAI21X1_583/Y gnd OAI21X1_584/Y vdd OAI21X1
XOAI21X1_562 INVX1_108/Y NOR2X1_101/Y OAI21X1_562/C gnd OAI21X1_562/Y vdd OAI21X1
XOAI21X1_595 BUFX4_148/Y INVX1_3/A OAI21X1_595/C gnd OAI21X1_596/C vdd OAI21X1
XFILL_48_1_1 gnd vdd FILL
XNAND2X1_590 MUX2X1_1/S NOR2X1_78/A gnd NAND2X1_590/Y vdd NAND2X1
XFILL_31_0_1 gnd vdd FILL
XFILL_39_1_1 gnd vdd FILL
XFILL_22_0_1 gnd vdd FILL
XBUFX4_209 BUFX4_25/Y gnd BUFX4_209/Y vdd BUFX4
XFILL_5_1_1 gnd vdd FILL
XFILL_42_8_0 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_381 BUFX4_171/Y NOR2X1_61/A INVX1_164/A gnd OAI21X1_382/C vdd OAI21X1
XOAI21X1_370 BUFX4_398/Y NAND2X1_80/Y OAI21X1_369/Y gnd OAI21X1_370/Y vdd OAI21X1
XOAI21X1_392 NAND2X1_81/Y BUFX4_380/Y OAI21X1_392/C gnd OAI21X1_392/Y vdd OAI21X1
XINVX1_401 INVX1_401/A gnd INVX1_401/Y vdd INVX1
XINVX1_434 INVX1_434/A gnd INVX1_434/Y vdd INVX1
XINVX1_423 INVX1_423/A gnd INVX1_423/Y vdd INVX1
XINVX1_412 INVX1_412/A gnd INVX1_412/Y vdd INVX1
XINVX1_456 INVX1_456/A gnd INVX1_456/Y vdd INVX1
XINVX1_467 INVX1_467/A gnd INVX1_467/Y vdd INVX1
XINVX1_445 INVX1_445/A gnd INVX1_445/Y vdd INVX1
XINVX1_478 INVX1_478/A gnd INVX1_478/Y vdd INVX1
XINVX1_489 INVX1_489/A gnd INVX1_489/Y vdd INVX1
XFILL_33_8_0 gnd vdd FILL
XOAI21X1_1611 BUFX4_395/Y NAND2X1_843/Y OAI21X1_1610/Y gnd DFFPOSX1_269/D vdd OAI21X1
XOAI21X1_1622 INVX1_270/Y NOR2X1_358/Y NAND2X1_848/Y gnd OAI21X1_1622/Y vdd OAI21X1
XOAI21X1_1600 BUFX4_454/Y BUFX4_346/Y INVX1_461/A gnd OAI21X1_1600/Y vdd OAI21X1
XOAI21X1_1633 INVX1_463/Y NOR2X1_368/Y NAND2X1_859/Y gnd OAI21X1_1633/Y vdd OAI21X1
XOAI21X1_1644 BUFX4_168/Y BUFX4_343/Y INVX1_336/A gnd OAI21X1_1645/C vdd OAI21X1
XOAI21X1_1655 BUFX4_114/Y NAND2X1_861/Y OAI21X1_1654/Y gnd OAI21X1_1655/Y vdd OAI21X1
XOAI21X1_1666 INVX1_24/Y NOR2X1_378/Y NAND2X1_863/Y gnd OAI21X1_1666/Y vdd OAI21X1
XOAI21X1_1699 BUFX4_401/Y NAND2X1_872/Y OAI21X1_1699/C gnd DFFPOSX1_349/D vdd OAI21X1
XOAI21X1_1688 BUFX4_406/Y OAI21X1_5/B INVX1_466/A gnd OAI21X1_1689/C vdd OAI21X1
XOAI21X1_1677 BUFX4_421/Y NAND2X1_871/Y OAI21X1_1677/C gnd DFFPOSX1_338/D vdd OAI21X1
XFILL_24_8_0 gnd vdd FILL
XMUX2X1_16 MUX2X1_16/A MUX2X1_16/B BUFX4_189/Y gnd MUX2X1_17/A vdd MUX2X1
XMUX2X1_27 MUX2X1_26/Y MUX2X1_25/Y BUFX4_32/Y gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_38 MUX2X1_38/A MUX2X1_38/B BUFX4_6/Y gnd MUX2X1_38/Y vdd MUX2X1
XMUX2X1_49 MUX2X1_49/A MUX2X1_49/B BUFX4_58/Y gnd MUX2X1_51/B vdd MUX2X1
XFILL_15_8_0 gnd vdd FILL
XDFFPOSX1_519 INVX1_413/A CLKBUF1_80/Y OAI21X1_238/Y gnd vdd DFFPOSX1
XDFFPOSX1_508 NOR2X1_36/A CLKBUF1_31/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XINVX1_231 INVX1_231/A gnd INVX1_231/Y vdd INVX1
XINVX1_253 INVX1_253/A gnd INVX1_253/Y vdd INVX1
XINVX1_220 INVX1_220/A gnd INVX1_220/Y vdd INVX1
XINVX1_242 INVX1_242/A gnd INVX1_242/Y vdd INVX1
XINVX1_286 INVX1_286/A gnd INVX1_286/Y vdd INVX1
XINVX1_275 INVX1_275/A gnd INVX1_275/Y vdd INVX1
XINVX1_264 INVX1_264/A gnd INVX1_264/Y vdd INVX1
XINVX1_297 INVX1_297/A gnd INVX1_297/Y vdd INVX1
XNAND2X1_31 BUFX4_163/Y NOR2X1_21/Y gnd NAND2X1_31/Y vdd NAND2X1
XNAND2X1_42 BUFX4_144/Y NOR2X1_31/Y gnd NAND2X1_42/Y vdd NAND2X1
XNAND2X1_20 NAND2X1_5/B BUFX4_288/Y gnd BUFX4_135/A vdd NAND2X1
XNAND2X1_75 BUFX4_137/Y NOR2X1_61/Y gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_86 INVX8_4/A NOR2X1_71/Y gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_64 BUFX4_136/Y NOR2X1_51/Y gnd NAND2X1_64/Y vdd NAND2X1
XNAND2X1_53 BUFX4_145/Y NOR2X1_41/Y gnd NAND2X1_53/Y vdd NAND2X1
XNAND2X1_97 INVX8_16/A INVX2_4/Y gnd NAND2X1_97/Y vdd NAND2X1
XFILL_42_1 gnd vdd FILL
XAOI21X1_213 BUFX4_285/Y NOR2X1_256/B NOR2X1_262/Y gnd DFFPOSX1_15/D vdd AOI21X1
XAOI21X1_224 BUFX4_423/Y NOR2X1_279/B NOR2X1_277/Y gnd DFFPOSX1_18/D vdd AOI21X1
XAOI21X1_202 NAND2X1_236/Y AOI21X1_202/B INVX2_6/Y gnd OAI21X1_822/B vdd AOI21X1
XAOI21X1_246 BUFX4_373/Y NOR2X1_303/B NOR2X1_307/Y gnd DFFPOSX1_96/D vdd AOI21X1
XAOI21X1_235 BUFX4_395/Y NOR2X1_289/B NOR2X1_290/Y gnd DFFPOSX1_61/D vdd AOI21X1
XAOI21X1_257 BUFX4_112/Y NOR2X1_325/B NOR2X1_325/Y gnd AOI21X1_257/Y vdd AOI21X1
XAOI21X1_279 BUFX4_424/Y NOR2X1_352/B NOR2X1_351/Y gnd AOI21X1_279/Y vdd AOI21X1
XAOI22X1_51 AOI22X1_51/A BUFX4_323/Y BUFX4_288/Y MUX2X1_246/Y gnd AOI22X1_51/Y vdd
+ AOI22X1
XAOI22X1_40 MUX2X1_189/Y BUFX4_354/Y BUFX4_155/Y AOI22X1_40/D gnd AOI22X1_40/Y vdd
+ AOI22X1
XAOI21X1_268 BUFX4_99/Y NOR2X1_338/B NOR2X1_338/Y gnd AOI21X1_268/Y vdd AOI21X1
XAOI22X1_73 AOI22X1_73/A BUFX4_320/Y BUFX4_292/Y AOI22X1_73/D gnd AOI22X1_73/Y vdd
+ AOI22X1
XAOI22X1_62 AOI22X1_62/A BUFX4_350/Y BUFX4_156/Y MUX2X1_300/Y gnd AOI22X1_62/Y vdd
+ AOI22X1
XOAI21X1_1441 INVX1_42/Y NOR2X1_321/Y NAND2X1_816/Y gnd OAI21X1_1441/Y vdd OAI21X1
XOAI21X1_1430 BUFX4_112/Y NAND2X1_815/Y OAI21X1_1429/Y gnd DFFPOSX1_139/D vdd OAI21X1
XOAI21X1_1463 BUFX4_167/Y BUFX4_393/Y INVX1_200/A gnd OAI21X1_1464/C vdd OAI21X1
XOAI21X1_1452 INVX1_199/Y NOR2X1_331/Y NAND2X1_827/Y gnd OAI21X1_1452/Y vdd OAI21X1
XOAI21X1_1474 BUFX4_125/Y NAND2X1_833/Y OAI21X1_1473/Y gnd OAI21X1_1474/Y vdd OAI21X1
XOAI21X1_1485 BUFX4_417/Y BUFX4_392/Y NAND2X1_628/B gnd OAI21X1_1485/Y vdd OAI21X1
XOAI21X1_1496 BUFX4_301/Y NAND2X1_834/Y OAI21X1_1496/C gnd DFFPOSX1_196/D vdd OAI21X1
XDFFPOSX1_1015 INVX1_444/A CLKBUF1_3/Y OAI21X1_797/Y gnd vdd DFFPOSX1
XDFFPOSX1_1004 NOR2X1_223/A CLKBUF1_73/Y AOI21X1_181/Y gnd vdd DFFPOSX1
XDFFPOSX1_1026 BUFX2_2/A CLKBUF1_65/Y NAND2X1_340/Y gnd vdd DFFPOSX1
XOAI22X1_2 MUX2X1_21/Y INVX1_10/Y INVX1_11/Y MUX2X1_28/Y gnd OAI22X1_2/Y vdd OAI22X1
XFILL_47_7_0 gnd vdd FILL
XFILL_30_6_0 gnd vdd FILL
XDFFPOSX1_316 NAND2X1_430/B CLKBUF1_32/Y OAI21X1_1657/Y gnd vdd DFFPOSX1
XDFFPOSX1_338 INVX1_82/A CLKBUF1_99/Y DFFPOSX1_338/D gnd vdd DFFPOSX1
XDFFPOSX1_327 INVX1_401/A CLKBUF1_6/Y DFFPOSX1_327/D gnd vdd DFFPOSX1
XDFFPOSX1_305 INVX1_17/A CLKBUF1_48/Y DFFPOSX1_305/D gnd vdd DFFPOSX1
XDFFPOSX1_349 NAND2X1_501/B CLKBUF1_38/Y DFFPOSX1_349/D gnd vdd DFFPOSX1
XNAND2X1_408 AOI22X1_27/Y AOI22X1_28/Y gnd AOI22X1_29/D vdd NAND2X1
XNAND2X1_419 BUFX4_258/Y NOR2X1_326/A gnd OAI21X1_986/C vdd NAND2X1
XFILL_38_7_0 gnd vdd FILL
XBUFX4_381 BUFX4_385/A gnd BUFX4_381/Y vdd BUFX4
XBUFX4_370 INVX8_15/Y gnd BUFX4_370/Y vdd BUFX4
XBUFX4_392 BUFX4_392/A gnd BUFX4_392/Y vdd BUFX4
XOAI21X1_914 INVX1_126/Y BUFX4_214/Y NAND2X1_342/Y gnd MUX2X1_91/A vdd OAI21X1
XOAI21X1_925 INVX1_137/Y BUFX4_236/Y NAND2X1_353/Y gnd MUX2X1_100/B vdd OAI21X1
XFILL_21_6_0 gnd vdd FILL
XOAI21X1_903 INVX1_115/Y BUFX4_192/Y OAI21X1_903/C gnd MUX2X1_83/B vdd OAI21X1
XOAI21X1_947 INVX1_159/Y MUX2X1_2/S OAI21X1_947/C gnd MUX2X1_116/B vdd OAI21X1
XOAI21X1_936 INVX1_148/Y BUFX4_258/Y NAND2X1_365/Y gnd MUX2X1_107/A vdd OAI21X1
XOAI21X1_958 INVX1_170/Y BUFX4_203/Y NAND2X1_388/Y gnd MUX2X1_124/A vdd OAI21X1
XOAI21X1_969 INVX1_181/Y BUFX4_225/Y NAND2X1_400/Y gnd MUX2X1_133/B vdd OAI21X1
XOAI21X1_1271 INVX1_483/Y BUFX4_235/Y NAND2X1_726/Y gnd MUX2X1_359/B vdd OAI21X1
XOAI21X1_1260 INVX1_472/Y BUFX4_213/Y NAND2X1_714/Y gnd MUX2X1_350/A vdd OAI21X1
XOAI21X1_1282 INVX1_494/Y BUFX4_257/Y NAND2X1_738/Y gnd MUX2X1_367/A vdd OAI21X1
XDFFPOSX1_850 INVX1_114/A CLKBUF1_54/Y OAI21X1_654/Y gnd vdd DFFPOSX1
XDFFPOSX1_861 NOR2X1_151/A CLKBUF1_95/Y AOI21X1_121/Y gnd vdd DFFPOSX1
XDFFPOSX1_883 INVX1_180/A CLKBUF1_84/Y OAI21X1_669/Y gnd vdd DFFPOSX1
XDFFPOSX1_872 INVX1_499/A CLKBUF1_81/Y OAI21X1_667/Y gnd vdd DFFPOSX1
XINVX2_11 INVX2_11/A gnd INVX2_11/Y vdd INVX2
XOAI21X1_1293 INVX1_505/Y MUX2X1_1/S NAND2X1_749/Y gnd MUX2X1_376/B vdd OAI21X1
XDFFPOSX1_894 NOR2X1_174/A CLKBUF1_13/Y AOI21X1_140/Y gnd vdd DFFPOSX1
XFILL_4_7_0 gnd vdd FILL
XFILL_29_7_0 gnd vdd FILL
XOAI21X1_18 BUFX4_128/Y NAND2X1_2/Y OAI21X1_17/Y gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 BUFX4_367/Y BUFX4_317/Y OAI21X1_29/C gnd OAI21X1_30/C vdd OAI21X1
XFILL_12_6_0 gnd vdd FILL
XDFFPOSX1_102 INVX1_323/A CLKBUF1_89/Y DFFPOSX1_102/D gnd vdd DFFPOSX1
XDFFPOSX1_113 INVX1_40/A CLKBUF1_42/Y OAI21X1_1378/Y gnd vdd DFFPOSX1
XDFFPOSX1_146 INVX1_70/A CLKBUF1_63/Y OAI21X1_1442/Y gnd vdd DFFPOSX1
XDFFPOSX1_135 INVX1_389/A CLKBUF1_102/Y OAI21X1_1422/Y gnd vdd DFFPOSX1
XDFFPOSX1_124 NAND2X1_417/B CLKBUF1_17/Y DFFPOSX1_124/D gnd vdd DFFPOSX1
XDFFPOSX1_179 INVX1_136/A CLKBUF1_78/Y OAI21X1_1462/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 NOR2X1_327/A CLKBUF1_98/Y AOI21X1_259/Y gnd vdd DFFPOSX1
XDFFPOSX1_168 INVX1_455/A CLKBUF1_55/Y OAI21X1_1456/Y gnd vdd DFFPOSX1
XNAND2X1_205 BUFX4_444/Y NOR2X1_228/Y gnd OAI21X1_795/C vdd NAND2X1
XNAND2X1_216 BUFX4_203/Y NOR2X1_360/A gnd OAI21X1_804/C vdd NAND2X1
XNAND2X1_227 NOR2X1_244/Y NAND2X1_227/B gnd NAND3X1_4/B vdd NAND2X1
XNAND2X1_238 BUFX4_82/Y NAND2X1_238/B gnd AOI21X1_202/B vdd NAND2X1
XNAND2X1_249 BUFX4_243/Y NOR2X1_323/A gnd OAI21X1_829/C vdd NAND2X1
XNOR2X1_260 NOR2X1_260/A NOR2X1_256/B gnd NOR2X1_260/Y vdd NOR2X1
XNOR2X1_271 NOR2X1_271/A NOR2X1_265/Y gnd NOR2X1_271/Y vdd NOR2X1
XNOR2X1_282 NOR2X1_282/A NOR2X1_279/B gnd NOR2X1_282/Y vdd NOR2X1
XNOR2X1_293 NOR2X1_293/A NOR2X1_289/B gnd NOR2X1_293/Y vdd NOR2X1
XOAI21X1_700 BUFX4_402/Y OAI21X1_704/B OAI21X1_699/Y gnd OAI21X1_700/Y vdd OAI21X1
XOAI21X1_711 INVX1_374/Y NOR2X1_177/Y OAI21X1_711/C gnd OAI21X1_711/Y vdd OAI21X1
XOAI21X1_722 INVX1_184/Y NOR2X1_199/Y OAI21X1_722/C gnd OAI21X1_722/Y vdd OAI21X1
XOAI21X1_733 BUFX4_110/Y OAI21X1_729/B OAI21X1_733/C gnd OAI21X1_733/Y vdd OAI21X1
XOAI21X1_755 BUFX4_103/Y OAI21X1_757/B OAI21X1_754/Y gnd OAI21X1_755/Y vdd OAI21X1
XOAI21X1_766 BUFX4_409/Y BUFX4_440/Y INVX1_250/A gnd OAI21X1_767/C vdd OAI21X1
XOAI21X1_744 NOR2X1_72/B INVX2_5/A MUX2X1_22/A gnd OAI21X1_745/C vdd OAI21X1
XOAI21X1_777 BUFX4_124/Y NAND2X1_201/Y OAI21X1_777/C gnd OAI21X1_777/Y vdd OAI21X1
XOAI21X1_788 NOR2X1_91/B BUFX4_442/Y INVX1_443/A gnd OAI21X1_789/C vdd OAI21X1
XOAI21X1_799 OAI22X1_1/Y OAI22X1_2/Y AOI22X1_69/C gnd NAND3X1_6/A vdd OAI21X1
XMUX2X1_222 MUX2X1_222/A MUX2X1_222/B BUFX4_363/Y gnd AOI22X1_46/D vdd MUX2X1
XMUX2X1_200 MUX2X1_200/A MUX2X1_200/B BUFX4_80/Y gnd MUX2X1_201/A vdd MUX2X1
XMUX2X1_211 MUX2X1_211/A MUX2X1_211/B BUFX4_61/Y gnd MUX2X1_213/B vdd MUX2X1
XMUX2X1_244 MUX2X1_244/A MUX2X1_244/B INVX4_1/A gnd MUX2X1_244/Y vdd MUX2X1
XMUX2X1_233 MUX2X1_233/A MUX2X1_233/B BUFX4_62/Y gnd MUX2X1_233/Y vdd MUX2X1
XMUX2X1_255 MUX2X1_255/A MUX2X1_255/B BUFX4_363/Y gnd AOI22X1_53/A vdd MUX2X1
XOAI21X1_1090 INVX1_302/Y BUFX4_269/Y NAND2X1_531/Y gnd MUX2X1_223/A vdd OAI21X1
XDFFPOSX1_691 INVX1_168/A CLKBUF1_58/Y OAI21X1_486/Y gnd vdd DFFPOSX1
XMUX2X1_299 MUX2X1_299/A MUX2X1_299/B BUFX4_45/Y gnd MUX2X1_299/Y vdd MUX2X1
XDFFPOSX1_680 INVX1_487/A CLKBUF1_47/Y OAI21X1_464/Y gnd vdd DFFPOSX1
XMUX2X1_266 MUX2X1_266/A MUX2X1_266/B INVX4_1/A gnd MUX2X1_266/Y vdd MUX2X1
XMUX2X1_277 MUX2X1_277/A MUX2X1_277/B BUFX4_44/Y gnd MUX2X1_279/B vdd MUX2X1
XMUX2X1_288 MUX2X1_288/A MUX2X1_288/B BUFX4_363/Y gnd AOI22X1_60/D vdd MUX2X1
XNAND2X1_772 BUFX4_139/Y NOR2X1_264/Y gnd NAND2X1_772/Y vdd NAND2X1
XNAND2X1_761 BUFX4_327/Y NOR2X1_254/Y gnd NAND2X1_761/Y vdd NAND2X1
XNAND2X1_750 MUX2X1_2/S NOR2X1_218/A gnd NAND2X1_750/Y vdd NAND2X1
XNAND2X1_794 INVX8_2/A NOR2X1_297/Y gnd NAND2X1_794/Y vdd NAND2X1
XNAND2X1_783 BUFX4_164/Y NOR2X1_284/Y gnd NAND2X1_783/Y vdd NAND2X1
XFILL_44_5_0 gnd vdd FILL
XCLKBUF1_19 BUFX4_18/Y gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX4_40 BUFX4_41/A gnd MUX2X1_3/S vdd BUFX4
XBUFX4_62 BUFX4_62/A gnd BUFX4_62/Y vdd BUFX4
XBUFX4_51 BUFX4_50/A gnd BUFX4_51/Y vdd BUFX4
XBUFX4_95 BUFX4_92/A gnd BUFX4_95/Y vdd BUFX4
XBUFX4_73 a[1] gnd BUFX4_50/A vdd BUFX4
XBUFX4_84 BUFX4_84/A gnd BUFX4_84/Y vdd BUFX4
XFILL_35_5_0 gnd vdd FILL
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XINVX8_10 INVX8_10/A gnd INVX8_10/Y vdd INVX8
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOAI21X1_541 BUFX4_148/Y BUFX4_295/Y OAI21X1_541/C gnd OAI21X1_542/C vdd OAI21X1
XOAI21X1_530 BUFX4_126/Y OAI21X1_544/B OAI21X1_529/Y gnd OAI21X1_530/Y vdd OAI21X1
XOAI21X1_563 INVX1_172/Y NOR2X1_101/Y OAI21X1_563/C gnd OAI21X1_563/Y vdd OAI21X1
XOAI21X1_574 BUFX4_110/Y OAI21X1_584/B OAI21X1_574/C gnd OAI21X1_574/Y vdd OAI21X1
XOAI21X1_552 INVX1_490/Y NOR2X1_81/Y NAND2X1_108/Y gnd OAI21X1_552/Y vdd OAI21X1
XOAI21X1_585 BUFX4_148/Y BUFX4_108/Y MUX2X1_1/A gnd OAI21X1_586/C vdd OAI21X1
XOAI21X1_596 BUFX4_104/Y OAI21X1_590/B OAI21X1_596/C gnd OAI21X1_596/Y vdd OAI21X1
.ends

